
// 	Fri Dec 23 03:30:12 2022
//	vlsi
//	localhost.localdomain

module datapath__0_9 (p_0, p_1);

output [63:0] p_1;
input [63:0] p_0;
wire n_127;
wire n_125;
wire n_126;
wire n_123;
wire n_124;
wire n_5;
wire n_3;
wire n_4;
wire n_1;
wire n_2;
wire n_120;
wire n_0;
wire n_121;
wire n_11;
wire n_119;
wire n_9;
wire n_10;
wire n_7;
wire n_8;
wire n_117;
wire n_6;
wire n_118;
wire n_17;
wire n_15;
wire n_16;
wire n_13;
wire n_14;
wire n_114;
wire n_12;
wire n_115;
wire n_112;
wire n_113;
wire n_110;
wire n_108;
wire n_109;
wire n_106;
wire n_107;
wire n_104;
wire n_105;
wire n_102;
wire n_103;
wire n_100;
wire n_101;
wire n_98;
wire n_99;
wire n_96;
wire n_97;
wire n_94;
wire n_92;
wire n_93;
wire n_90;
wire n_91;
wire n_88;
wire n_89;
wire n_86;
wire n_84;
wire n_85;
wire n_82;
wire n_83;
wire n_23;
wire n_81;
wire n_21;
wire n_22;
wire n_19;
wire n_20;
wire n_31;
wire n_18;
wire n_29;
wire n_30;
wire n_27;
wire n_28;
wire n_25;
wire n_26;
wire n_77;
wire n_24;
wire n_79;
wire n_37;
wire n_76;
wire n_35;
wire n_36;
wire n_33;
wire n_34;
wire n_75;
wire n_32;
wire n_80;
wire n_73;
wire n_74;
wire n_71;
wire n_72;
wire n_69;
wire n_70;
wire n_67;
wire n_68;
wire n_43;
wire n_66;
wire n_41;
wire n_42;
wire n_45;
wire n_49;
wire n_44;
wire n_46;
wire n_129;
wire n_48;
wire n_62;
wire n_47;
wire n_63;
wire n_51;
wire n_61;
wire n_54;
wire n_52;
wire n_65;
wire n_162;
wire n_60;
wire n_161;
wire n_172;
wire n_173;
wire n_185;
wire n_58;
wire n_39;
wire n_38;
wire n_40;
wire n_50;
wire n_53;
wire n_64;
wire n_55;
wire n_56;
wire n_57;
wire n_59;
wire n_184;
wire n_183;
wire n_141;
wire n_140;
wire n_132;
wire n_134;
wire n_209;
wire n_207;
wire n_78;
wire n_204;
wire n_201;
wire n_198;
wire n_195;
wire n_128;
wire n_192;
wire n_179;
wire n_178;
wire n_181;
wire n_190;
wire n_189;
wire n_188;
wire n_130;
wire n_131;
wire n_133;
wire n_135;
wire n_137;
wire n_136;
wire n_139;
wire n_212;
wire n_160;
wire n_147;
wire n_142;
wire n_143;
wire n_145;
wire n_144;
wire n_148;
wire n_213;
wire n_146;
wire n_152;
wire n_154;
wire n_164;
wire n_158;
wire n_211;
wire n_210;
wire n_208;
wire n_166;
wire n_206;
wire n_205;
wire n_203;
wire n_202;
wire n_149;
wire n_200;
wire n_199;
wire n_197;
wire n_196;
wire n_194;
wire n_193;
wire n_176;
wire n_170;
wire n_153;
wire n_155;
wire n_156;
wire n_157;
wire n_159;
wire n_165;
wire n_167;
wire n_171;
wire n_174;
wire n_175;
wire n_177;
wire n_180;
wire n_182;
wire n_186;
wire n_187;
wire n_191;


INV_X1 i_276 (.ZN (n_213), .A (p_0[60]));
INV_X1 i_275 (.ZN (n_212), .A (p_0[47]));
INV_X1 i_274 (.ZN (n_211), .A (p_0[46]));
INV_X1 i_273 (.ZN (n_210), .A (p_0[45]));
INV_X1 i_272 (.ZN (n_209), .A (p_0[44]));
INV_X1 i_271 (.ZN (n_208), .A (n_50));
INV_X1 i_270 (.ZN (n_207), .A (p_0[31]));
INV_X1 i_269 (.ZN (n_206), .A (p_0[30]));
INV_X1 i_268 (.ZN (n_205), .A (p_0[29]));
INV_X1 i_267 (.ZN (n_204), .A (p_0[28]));
INV_X1 i_266 (.ZN (n_203), .A (p_0[27]));
INV_X1 i_265 (.ZN (n_202), .A (p_0[26]));
INV_X1 i_264 (.ZN (n_201), .A (p_0[25]));
INV_X1 i_263 (.ZN (n_200), .A (p_0[24]));
INV_X1 i_262 (.ZN (n_199), .A (p_0[23]));
INV_X1 i_261 (.ZN (n_198), .A (p_0[22]));
INV_X1 i_260 (.ZN (n_197), .A (p_0[21]));
INV_X1 i_259 (.ZN (n_196), .A (p_0[20]));
INV_X1 i_258 (.ZN (n_195), .A (p_0[19]));
INV_X1 i_257 (.ZN (n_194), .A (p_0[18]));
INV_X1 i_256 (.ZN (n_193), .A (p_0[17]));
INV_X1 i_255 (.ZN (n_192), .A (p_0[16]));
INV_X1 i_254 (.ZN (n_191), .A (p_0[3]));
INV_X1 i_253 (.ZN (n_190), .A (p_0[2]));
INV_X1 i_252 (.ZN (n_189), .A (p_0[1]));
INV_X1 i_251 (.ZN (n_188), .A (p_0[0]));
NAND4_X1 i_250 (.ZN (n_187), .A1 (n_191), .A2 (n_190), .A3 (n_189), .A4 (n_188));
INV_X1 i_249 (.ZN (n_123), .A (n_187));
INV_X1 i_248 (.ZN (n_186), .A (p_0[7]));
INV_X1 i_247 (.ZN (n_185), .A (p_0[6]));
INV_X1 i_246 (.ZN (n_184), .A (p_0[5]));
INV_X1 i_245 (.ZN (n_183), .A (p_0[4]));
NAND4_X1 i_244 (.ZN (n_182), .A1 (n_186), .A2 (n_185), .A3 (n_184), .A4 (n_183));
INV_X1 i_243 (.ZN (n_181), .A (n_182));
INV_X1 i_242 (.ZN (n_180), .A (p_0[11]));
INV_X1 i_241 (.ZN (n_179), .A (p_0[8]));
INV_X1 i_240 (.ZN (n_178), .A (n_57));
NAND3_X1 i_239 (.ZN (n_177), .A1 (n_180), .A2 (n_179), .A3 (n_178));
INV_X1 i_238 (.ZN (n_176), .A (n_177));
NAND3_X1 i_237 (.ZN (n_175), .A1 (n_123), .A2 (n_181), .A3 (n_176));
INV_X1 i_236 (.ZN (n_117), .A (n_175));
INV_X1 i_235 (.ZN (n_174), .A (p_0[15]));
INV_X1 i_234 (.ZN (n_173), .A (p_0[12]));
INV_X1 i_233 (.ZN (n_172), .A (n_56));
NAND3_X1 i_232 (.ZN (n_171), .A1 (n_174), .A2 (n_173), .A3 (n_172));
INV_X1 i_231 (.ZN (n_170), .A (n_171));
NAND4_X1 i_230 (.ZN (n_109), .A1 (n_117), .A2 (n_193), .A3 (n_192), .A4 (n_170));
NAND4_X1 i_228 (.ZN (n_103), .A1 (n_110), .A2 (n_196), .A3 (n_195), .A4 (n_194));
INV_X1 i_227 (.ZN (n_104), .A (n_103));
NAND4_X1 i_226 (.ZN (n_97), .A1 (n_104), .A2 (n_199), .A3 (n_198), .A4 (n_197));
INV_X1 i_225 (.ZN (n_98), .A (n_97));
NAND4_X1 i_224 (.ZN (n_91), .A1 (n_98), .A2 (n_202), .A3 (n_201), .A4 (n_200));
NAND4_X1 i_222 (.ZN (n_85), .A1 (n_92), .A2 (n_205), .A3 (n_204), .A4 (n_203));
INV_X1 i_221 (.ZN (n_86), .A (n_85));
OR3_X1 i_220 (.ZN (n_167), .A1 (p_0[39]), .A2 (p_0[38]), .A3 (n_53));
INV_X1 i_219 (.ZN (n_166), .A (n_167));
NAND4_X1 i_218 (.ZN (n_76), .A1 (n_86), .A2 (n_207), .A3 (n_206), .A4 (n_166));
INV_X1 i_217 (.ZN (n_77), .A (n_76));
NAND4_X1 i_216 (.ZN (n_70), .A1 (n_77), .A2 (n_210), .A3 (n_209), .A4 (n_208));
INV_X1 i_215 (.ZN (n_71), .A (n_70));
OR2_X1 i_214 (.ZN (n_165), .A1 (p_0[55]), .A2 (n_55));
INV_X1 i_213 (.ZN (n_164), .A (n_165));
NAND4_X1 i_212 (.ZN (n_61), .A1 (n_71), .A2 (n_212), .A3 (n_211), .A4 (n_164));
INV_X1 i_210 (.ZN (n_162), .A (p_0[57]));
INV_X1 i_209 (.ZN (n_161), .A (p_0[56]));
NAND2_X1 i_208 (.ZN (n_160), .A1 (n_162), .A2 (n_161));
OR3_X1 i_207 (.ZN (n_159), .A1 (n_160), .A2 (p_0[59]), .A3 (p_0[58]));
INV_X1 i_206 (.ZN (n_158), .A (n_159));
OR2_X1 i_205 (.ZN (n_157), .A1 (p_0[62]), .A2 (p_0[61]));
INV_X1 i_204 (.ZN (n_156), .A (n_157));
NAND4_X1 i_203 (.ZN (p_1[63]), .A1 (n_62), .A2 (n_213), .A3 (n_158), .A4 (n_156));
INV_X1 i_202 (.ZN (n_155), .A (p_1[63]));
INV_X1 i_201 (.ZN (n_154), .A (p_0[61]));
NAND4_X1 i_200 (.ZN (n_153), .A1 (n_62), .A2 (n_154), .A3 (n_213), .A4 (n_158));
AOI21_X1 i_199 (.ZN (p_1[62]), .A (n_155), .B1 (n_153), .B2 (p_0[62]));
INV_X1 i_198 (.ZN (n_152), .A (n_153));
NAND4_X1 i_197 (.ZN (n_113), .A1 (n_123), .A2 (n_181), .A3 (n_176), .A4 (n_170));
NAND4_X1 i_195 (.ZN (n_107), .A1 (n_114), .A2 (n_194), .A3 (n_193), .A4 (n_192));
NAND4_X1 i_193 (.ZN (n_101), .A1 (n_108), .A2 (n_197), .A3 (n_196), .A4 (n_195));
INV_X1 i_191 (.ZN (n_102), .A (n_101));
NAND4_X1 i_190 (.ZN (n_149), .A1 (n_102), .A2 (n_200), .A3 (n_199), .A4 (n_198));
INV_X1 i_189 (.ZN (n_96), .A (n_149));
NAND4_X1 i_188 (.ZN (n_89), .A1 (n_96), .A2 (n_203), .A3 (n_202), .A4 (n_201));
INV_X1 i_187 (.ZN (n_90), .A (n_89));
NAND4_X1 i_186 (.ZN (n_83), .A1 (n_90), .A2 (n_206), .A3 (n_205), .A4 (n_204));
INV_X1 i_185 (.ZN (n_84), .A (n_83));
NAND4_X1 i_184 (.ZN (n_74), .A1 (n_84), .A2 (n_207), .A3 (n_208), .A4 (n_166));
INV_X1 i_183 (.ZN (n_75), .A (n_74));
NAND4_X1 i_182 (.ZN (n_68), .A1 (n_75), .A2 (n_211), .A3 (n_210), .A4 (n_209));
INV_X1 i_181 (.ZN (n_69), .A (n_68));
NAND4_X1 i_180 (.ZN (n_148), .A1 (n_69), .A2 (n_212), .A3 (n_164), .A4 (n_158));
INV_X1 i_179 (.ZN (n_147), .A (n_148));
AOI21_X1 i_178 (.ZN (n_146), .A (n_154), .B1 (n_147), .B2 (n_213));
NOR2_X1 i_177 (.ZN (p_1[61]), .A1 (n_146), .A2 (n_152));
NAND2_X1 i_176 (.ZN (n_145), .A1 (n_147), .A2 (n_213));
NAND2_X1 i_175 (.ZN (n_144), .A1 (n_148), .A2 (p_0[60]));
NAND2_X1 i_174 (.ZN (n_143), .A1 (n_145), .A2 (n_144));
INV_X1 i_173 (.ZN (p_1[60]), .A (n_143));
INV_X1 i_172 (.ZN (n_142), .A (n_54));
AOI21_X1 i_171 (.ZN (p_1[59]), .A (n_147), .B1 (p_0[59]), .B2 (n_142));
INV_X1 i_170 (.ZN (n_141), .A (n_160));
NAND2_X1 i_169 (.ZN (n_140), .A1 (n_62), .A2 (n_161));
AOI22_X1 i_168 (.ZN (p_1[57]), .A1 (n_140), .A2 (p_0[57]), .B1 (n_62), .B2 (n_141));
INV_X1 i_167 (.ZN (n_139), .A (n_64));
NAND2_X1 i_166 (.ZN (n_66), .A1 (n_69), .A2 (n_212));
NAND2_X1 i_164 (.ZN (n_49), .A1 (n_67), .A2 (n_139));
INV_X1 i_163 (.ZN (n_137), .A (n_49));
INV_X1 i_162 (.ZN (n_136), .A (p_0[50]));
INV_X1 i_161 (.ZN (n_135), .A (p_0[49]));
INV_X1 i_160 (.ZN (n_134), .A (p_0[48]));
NAND4_X1 i_159 (.ZN (n_133), .A1 (n_67), .A2 (n_136), .A3 (n_135), .A4 (n_134));
AOI21_X1 i_158 (.ZN (p_1[51]), .A (n_137), .B1 (n_133), .B2 (p_0[51]));
NAND3_X1 i_157 (.ZN (n_132), .A1 (n_67), .A2 (n_135), .A3 (n_134));
NAND2_X1 i_156 (.ZN (n_131), .A1 (n_132), .A2 (p_0[50]));
NAND2_X1 i_155 (.ZN (n_130), .A1 (n_131), .A2 (n_133));
INV_X1 i_154 (.ZN (p_1[50]), .A (n_130));
NAND2_X1 i_153 (.ZN (n_126), .A1 (n_189), .A2 (n_188));
INV_X1 i_152 (.ZN (n_127), .A (n_126));
NAND2_X1 i_151 (.ZN (n_124), .A1 (n_127), .A2 (n_190));
INV_X1 i_150 (.ZN (n_125), .A (n_124));
NAND2_X1 i_149 (.ZN (n_119), .A1 (n_123), .A2 (n_181));
NAND2_X1 i_148 (.ZN (n_118), .A1 (n_179), .A2 (n_178));
NAND2_X1 i_147 (.ZN (n_128), .A1 (n_114), .A2 (n_192));
INV_X1 i_146 (.ZN (n_112), .A (n_128));
NAND2_X1 i_145 (.ZN (n_105), .A1 (n_108), .A2 (n_195));
INV_X1 i_144 (.ZN (n_106), .A (n_105));
NAND2_X1 i_143 (.ZN (n_99), .A1 (n_102), .A2 (n_198));
INV_X1 i_142 (.ZN (n_100), .A (n_99));
NAND2_X1 i_141 (.ZN (n_93), .A1 (n_96), .A2 (n_201));
NAND2_X1 i_140 (.ZN (n_78), .A1 (n_90), .A2 (n_204));
INV_X1 i_139 (.ZN (n_88), .A (n_78));
NAND2_X1 i_138 (.ZN (n_81), .A1 (n_84), .A2 (n_207));
INV_X1 i_137 (.ZN (n_82), .A (n_81));
NAND2_X1 i_136 (.ZN (n_72), .A1 (n_75), .A2 (n_209));
INV_X1 i_135 (.ZN (n_73), .A (n_72));
NAND2_X1 i_134 (.ZN (n_42), .A1 (n_67), .A2 (n_134));
INV_X1 i_133 (.ZN (n_43), .A (n_42));
INV_X1 i_132 (.ZN (n_41), .A (n_132));
INV_X1 i_131 (.ZN (n_51), .A (n_140));
NAND2_X1 i_130 (.ZN (n_52), .A1 (n_62), .A2 (n_141));
INV_X1 i_129 (.ZN (n_60), .A (p_0[58]));
NAND2_X1 i_128 (.ZN (n_59), .A1 (n_184), .A2 (n_183));
INV_X1 i_127 (.ZN (n_58), .A (n_59));
OR2_X1 i_126 (.ZN (n_57), .A1 (p_0[10]), .A2 (p_0[9]));
OR2_X1 i_125 (.ZN (n_56), .A1 (p_0[13]), .A2 (p_0[14]));
OR3_X1 i_124 (.ZN (n_63), .A1 (p_0[53]), .A2 (p_0[54]), .A3 (p_0[52]));
NAND2_X1 i_123 (.ZN (n_64), .A1 (n_38), .A2 (n_40));
OR2_X1 i_122 (.ZN (n_55), .A1 (n_63), .A2 (n_64));
INV_X1 i_121 (.ZN (n_110), .A (n_109));
INV_X1 i_120 (.ZN (n_94), .A (n_93));
INV_X1 i_119 (.ZN (n_62), .A (n_61));
OR4_X1 i_118 (.ZN (n_79), .A1 (p_0[35]), .A2 (p_0[34]), .A3 (p_0[33]), .A4 (p_0[32]));
OR3_X1 i_117 (.ZN (n_53), .A1 (n_79), .A2 (p_0[36]), .A3 (p_0[37]));
OR3_X1 i_116 (.ZN (n_80), .A1 (p_0[42]), .A2 (p_0[41]), .A3 (p_0[40]));
OR2_X1 i_115 (.ZN (n_50), .A1 (n_80), .A2 (p_0[43]));
INV_X1 i_114 (.ZN (n_40), .A (p_0[51]));
OR3_X1 i_112 (.ZN (n_39), .A1 (p_0[50]), .A2 (p_0[49]), .A3 (p_0[48]));
INV_X1 i_111 (.ZN (n_38), .A (n_39));
INV_X1 i_108 (.ZN (n_120), .A (n_119));
NAND2_X1 i_107 (.ZN (n_121), .A1 (n_185), .A2 (n_58));
INV_X1 i_104 (.ZN (n_114), .A (n_113));
NAND2_X1 i_94 (.ZN (n_115), .A1 (n_172), .A2 (n_173));
INV_X1 i_92 (.ZN (n_108), .A (n_107));
INV_X1 i_90 (.ZN (n_92), .A (n_91));
INV_X1 i_88 (.ZN (n_67), .A (n_66));
NAND3_X1 i_87 (.ZN (n_65), .A1 (n_162), .A2 (n_60), .A3 (n_161));
INV_X1 i_192 (.ZN (n_129), .A (p_0[53]));
NOR2_X1 i_113 (.ZN (n_54), .A1 (n_65), .A2 (n_61));
AOI21_X1 i_109 (.ZN (p_1[58]), .A (n_54), .B1 (p_0[58]), .B2 (n_52));
AOI21_X1 i_105 (.ZN (p_1[56]), .A (n_51), .B1 (p_0[56]), .B2 (n_61));
NOR2_X1 i_103 (.ZN (n_48), .A1 (n_63), .A2 (n_49));
INV_X1 i_102 (.ZN (n_47), .A (n_48));
AOI21_X1 i_101 (.ZN (p_1[55]), .A (n_62), .B1 (p_0[55]), .B2 (n_47));
OR3_X1 i_100 (.ZN (n_46), .A1 (p_0[53]), .A2 (p_0[52]), .A3 (n_49));
AOI21_X1 i_99 (.ZN (p_1[54]), .A (n_48), .B1 (p_0[54]), .B2 (n_46));
NOR2_X1 i_98 (.ZN (n_45), .A1 (p_0[52]), .A2 (n_49));
OAI21_X1 i_97 (.ZN (n_44), .A (n_46), .B1 (n_129), .B2 (n_45));
INV_X1 i_96 (.ZN (p_1[53]), .A (n_44));
AOI21_X1 i_95 (.ZN (p_1[52]), .A (n_45), .B1 (p_0[52]), .B2 (n_49));
AOI21_X1 i_86 (.ZN (p_1[49]), .A (n_41), .B1 (p_0[49]), .B2 (n_42));
AOI21_X1 i_85 (.ZN (p_1[48]), .A (n_43), .B1 (p_0[48]), .B2 (n_66));
AOI21_X1 i_84 (.ZN (p_1[47]), .A (n_67), .B1 (p_0[47]), .B2 (n_68));
AOI21_X1 i_83 (.ZN (p_1[46]), .A (n_69), .B1 (p_0[46]), .B2 (n_70));
AOI21_X1 i_82 (.ZN (p_1[45]), .A (n_71), .B1 (p_0[45]), .B2 (n_72));
AOI21_X1 i_81 (.ZN (p_1[44]), .A (n_73), .B1 (p_0[44]), .B2 (n_74));
NOR2_X1 i_80 (.ZN (n_37), .A1 (p_0[40]), .A2 (n_76));
INV_X1 i_79 (.ZN (n_36), .A (n_37));
NOR2_X1 i_78 (.ZN (n_35), .A1 (p_0[41]), .A2 (n_36));
INV_X1 i_77 (.ZN (n_34), .A (n_35));
NOR2_X1 i_76 (.ZN (n_33), .A1 (n_80), .A2 (n_76));
INV_X1 i_75 (.ZN (n_32), .A (n_33));
AOI21_X1 i_74 (.ZN (p_1[43]), .A (n_75), .B1 (p_0[43]), .B2 (n_32));
AOI21_X1 i_73 (.ZN (p_1[42]), .A (n_33), .B1 (p_0[42]), .B2 (n_34));
AOI21_X1 i_72 (.ZN (p_1[41]), .A (n_35), .B1 (p_0[41]), .B2 (n_36));
AOI21_X1 i_71 (.ZN (p_1[40]), .A (n_37), .B1 (p_0[40]), .B2 (n_76));
NOR2_X1 i_70 (.ZN (n_31), .A1 (n_81), .A2 (n_79));
INV_X1 i_69 (.ZN (n_30), .A (n_31));
NOR2_X1 i_68 (.ZN (n_29), .A1 (p_0[36]), .A2 (n_30));
INV_X1 i_67 (.ZN (n_28), .A (n_29));
NOR2_X1 i_66 (.ZN (n_27), .A1 (p_0[37]), .A2 (n_28));
INV_X1 i_65 (.ZN (n_26), .A (n_27));
NOR2_X1 i_64 (.ZN (n_25), .A1 (p_0[38]), .A2 (n_26));
INV_X1 i_63 (.ZN (n_24), .A (n_25));
AOI21_X1 i_62 (.ZN (p_1[39]), .A (n_77), .B1 (p_0[39]), .B2 (n_24));
AOI21_X1 i_61 (.ZN (p_1[38]), .A (n_25), .B1 (p_0[38]), .B2 (n_26));
AOI21_X1 i_60 (.ZN (p_1[37]), .A (n_27), .B1 (p_0[37]), .B2 (n_28));
AOI21_X1 i_59 (.ZN (p_1[36]), .A (n_29), .B1 (p_0[36]), .B2 (n_30));
NOR2_X1 i_58 (.ZN (n_23), .A1 (p_0[32]), .A2 (n_81));
INV_X1 i_57 (.ZN (n_22), .A (n_23));
NOR2_X1 i_56 (.ZN (n_21), .A1 (p_0[33]), .A2 (n_22));
INV_X1 i_55 (.ZN (n_20), .A (n_21));
NOR2_X1 i_54 (.ZN (n_19), .A1 (p_0[34]), .A2 (n_20));
INV_X1 i_53 (.ZN (n_18), .A (n_19));
AOI21_X1 i_52 (.ZN (p_1[35]), .A (n_31), .B1 (p_0[35]), .B2 (n_18));
AOI21_X1 i_51 (.ZN (p_1[34]), .A (n_19), .B1 (p_0[34]), .B2 (n_20));
AOI21_X1 i_50 (.ZN (p_1[33]), .A (n_21), .B1 (p_0[33]), .B2 (n_22));
AOI21_X1 i_49 (.ZN (p_1[32]), .A (n_23), .B1 (p_0[32]), .B2 (n_81));
AOI21_X1 i_48 (.ZN (p_1[31]), .A (n_82), .B1 (p_0[31]), .B2 (n_83));
AOI21_X1 i_47 (.ZN (p_1[30]), .A (n_84), .B1 (p_0[30]), .B2 (n_85));
AOI21_X1 i_46 (.ZN (p_1[29]), .A (n_86), .B1 (p_0[29]), .B2 (n_78));
AOI21_X1 i_45 (.ZN (p_1[28]), .A (n_88), .B1 (p_0[28]), .B2 (n_89));
AOI21_X1 i_44 (.ZN (p_1[27]), .A (n_90), .B1 (p_0[27]), .B2 (n_91));
AOI21_X1 i_43 (.ZN (p_1[26]), .A (n_92), .B1 (p_0[26]), .B2 (n_93));
AOI21_X1 i_42 (.ZN (p_1[25]), .A (n_94), .B1 (p_0[25]), .B2 (n_149));
AOI21_X1 i_41 (.ZN (p_1[24]), .A (n_96), .B1 (p_0[24]), .B2 (n_97));
AOI21_X1 i_40 (.ZN (p_1[23]), .A (n_98), .B1 (p_0[23]), .B2 (n_99));
AOI21_X1 i_39 (.ZN (p_1[22]), .A (n_100), .B1 (p_0[22]), .B2 (n_101));
AOI21_X1 i_38 (.ZN (p_1[21]), .A (n_102), .B1 (p_0[21]), .B2 (n_103));
AOI21_X1 i_37 (.ZN (p_1[20]), .A (n_104), .B1 (p_0[20]), .B2 (n_105));
AOI21_X1 i_36 (.ZN (p_1[19]), .A (n_106), .B1 (p_0[19]), .B2 (n_107));
AOI21_X1 i_35 (.ZN (p_1[18]), .A (n_108), .B1 (p_0[18]), .B2 (n_109));
AOI21_X1 i_34 (.ZN (p_1[17]), .A (n_110), .B1 (p_0[17]), .B2 (n_128));
AOI21_X1 i_33 (.ZN (p_1[16]), .A (n_112), .B1 (p_0[16]), .B2 (n_113));
NOR2_X1 i_32 (.ZN (n_17), .A1 (p_0[12]), .A2 (n_175));
INV_X1 i_31 (.ZN (n_16), .A (n_17));
NOR2_X1 i_30 (.ZN (n_15), .A1 (p_0[13]), .A2 (n_16));
INV_X1 i_29 (.ZN (n_14), .A (n_15));
NOR2_X1 i_28 (.ZN (n_13), .A1 (n_175), .A2 (n_115));
INV_X1 i_27 (.ZN (n_12), .A (n_13));
AOI21_X1 i_26 (.ZN (p_1[15]), .A (n_114), .B1 (p_0[15]), .B2 (n_12));
AOI21_X1 i_25 (.ZN (p_1[14]), .A (n_13), .B1 (p_0[14]), .B2 (n_14));
AOI21_X1 i_24 (.ZN (p_1[13]), .A (n_15), .B1 (p_0[13]), .B2 (n_16));
AOI21_X1 i_23 (.ZN (p_1[12]), .A (n_17), .B1 (p_0[12]), .B2 (n_175));
NOR2_X1 i_22 (.ZN (n_11), .A1 (p_0[8]), .A2 (n_119));
INV_X1 i_21 (.ZN (n_10), .A (n_11));
NOR2_X1 i_20 (.ZN (n_9), .A1 (p_0[9]), .A2 (n_10));
INV_X1 i_19 (.ZN (n_8), .A (n_9));
NOR2_X1 i_18 (.ZN (n_7), .A1 (n_119), .A2 (n_118));
INV_X1 i_17 (.ZN (n_6), .A (n_7));
AOI21_X1 i_16 (.ZN (p_1[11]), .A (n_117), .B1 (p_0[11]), .B2 (n_6));
AOI21_X1 i_15 (.ZN (p_1[10]), .A (n_7), .B1 (p_0[10]), .B2 (n_8));
AOI21_X1 i_14 (.ZN (p_1[9]), .A (n_9), .B1 (p_0[9]), .B2 (n_10));
AOI21_X1 i_13 (.ZN (p_1[8]), .A (n_11), .B1 (p_0[8]), .B2 (n_119));
NOR2_X1 i_12 (.ZN (n_5), .A1 (p_0[4]), .A2 (n_187));
INV_X1 i_11 (.ZN (n_4), .A (n_5));
NOR2_X1 i_10 (.ZN (n_3), .A1 (p_0[5]), .A2 (n_4));
INV_X1 i_9 (.ZN (n_2), .A (n_3));
NOR2_X1 i_8 (.ZN (n_1), .A1 (n_187), .A2 (n_121));
INV_X1 i_7 (.ZN (n_0), .A (n_1));
AOI21_X1 i_6 (.ZN (p_1[7]), .A (n_120), .B1 (p_0[7]), .B2 (n_0));
AOI21_X1 i_5 (.ZN (p_1[6]), .A (n_1), .B1 (p_0[6]), .B2 (n_2));
AOI21_X1 i_4 (.ZN (p_1[5]), .A (n_3), .B1 (p_0[5]), .B2 (n_4));
AOI21_X1 i_3 (.ZN (p_1[4]), .A (n_5), .B1 (p_0[4]), .B2 (n_187));
AOI21_X1 i_2 (.ZN (p_1[3]), .A (n_123), .B1 (p_0[3]), .B2 (n_124));
AOI21_X1 i_1 (.ZN (p_1[2]), .A (n_125), .B1 (p_0[2]), .B2 (n_126));
AOI21_X1 i_0 (.ZN (p_1[1]), .A (n_127), .B1 (p_0[1]), .B2 (p_0[0]));

endmodule //datapath__0_9

module datapath__0_6 (p_0, Accumulator, Accumulator1);

output [31:0] Accumulator1;
input [31:0] Accumulator;
input [31:0] p_0;
wire n_0;
wire n_159;
wire n_1;
wire n_158;
wire n_157;
wire n_2;
wire n_162;
wire n_156;
wire n_3;
wire n_163;
wire n_168;
wire n_165;
wire n_154;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_151;
wire n_142;
wire n_11;
wire n_5;
wire n_152;
wire n_146;
wire n_8;
wire n_149;
wire n_147;
wire n_153;
wire n_144;
wire n_140;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_137;
wire n_128;
wire n_19;
wire n_13;
wire n_138;
wire n_132;
wire n_16;
wire n_135;
wire n_133;
wire n_139;
wire n_130;
wire n_126;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_123;
wire n_114;
wire n_27;
wire n_21;
wire n_124;
wire n_118;
wire n_24;
wire n_121;
wire n_119;
wire n_125;
wire n_116;
wire n_112;
wire n_34;
wire n_33;
wire n_30;
wire n_31;
wire n_28;
wire n_109;
wire n_100;
wire n_35;
wire n_29;
wire n_110;
wire n_104;
wire n_32;
wire n_107;
wire n_105;
wire n_111;
wire n_102;
wire n_98;
wire n_42;
wire n_41;
wire n_38;
wire n_39;
wire n_36;
wire n_87;
wire n_77;
wire n_43;
wire n_37;
wire n_86;
wire n_89;
wire n_79;
wire n_40;
wire n_88;
wire n_84;
wire n_81;
wire n_91;
wire n_52;
wire n_51;
wire n_74;
wire n_66;
wire n_65;
wire n_63;
wire n_59;
wire n_64;
wire n_58;
wire n_60;
wire n_170;
wire n_167;
wire n_80;
wire n_101;
wire n_99;
wire n_108;
wire n_103;
wire n_106;
wire n_113;
wire n_117;
wire n_120;
wire n_115;
wire n_122;
wire n_127;
wire n_131;
wire n_134;
wire n_129;
wire n_136;
wire n_141;
wire n_145;
wire n_148;
wire n_143;
wire n_150;
wire n_155;
wire n_161;
wire n_160;
wire n_166;
wire n_169;
wire n_44;
wire n_45;
wire n_185;
wire n_184;
wire n_46;
wire n_53;
wire n_55;
wire n_95;
wire n_49;
wire n_47;
wire n_57;
wire n_92;
wire n_61;
wire n_48;
wire n_56;
wire n_50;
wire n_96;
wire n_54;
wire n_181;
wire n_180;
wire n_179;
wire n_182;
wire n_62;
wire n_67;
wire n_70;
wire n_68;
wire n_82;
wire n_69;
wire n_187;
wire n_78;
wire n_71;
wire n_73;
wire n_72;
wire n_75;
wire n_188;
wire n_186;
wire n_76;
wire n_83;
wire n_93;
wire n_85;
wire n_177;
wire n_90;
wire n_183;
wire n_178;
wire n_94;
wire n_174;
wire n_172;
wire n_171;
wire n_97;
wire n_164;
wire n_176;
wire n_173;
wire n_175;


INV_X1 i_220 (.ZN (n_188), .A (p_0[31]));
OR2_X1 i_219 (.ZN (n_187), .A1 (p_0[30]), .A2 (Accumulator[30]));
NAND2_X1 i_218 (.ZN (n_60), .A1 (n_170), .A2 (n_167));
NAND2_X1 i_217 (.ZN (n_186), .A1 (n_59), .A2 (n_60));
NAND2_X1 i_216 (.ZN (n_185), .A1 (p_0[28]), .A2 (Accumulator[28]));
NOR2_X1 i_215 (.ZN (n_184), .A1 (p_0[28]), .A2 (Accumulator[28]));
NOR2_X1 i_214 (.ZN (n_183), .A1 (p_0[27]), .A2 (Accumulator[27]));
INV_X1 i_213 (.ZN (n_182), .A (n_183));
INV_X1 i_212 (.ZN (n_181), .A (p_0[25]));
INV_X1 i_211 (.ZN (n_180), .A (Accumulator[25]));
NOR2_X1 i_210 (.ZN (n_179), .A1 (p_0[26]), .A2 (Accumulator[26]));
AOI21_X1 i_209 (.ZN (n_178), .A (n_179), .B1 (n_181), .B2 (n_180));
NAND2_X1 i_208 (.ZN (n_177), .A1 (n_182), .A2 (n_178));
NOR2_X1 i_207 (.ZN (n_91), .A1 (p_0[23]), .A2 (Accumulator[23]));
NOR3_X1 i_206 (.ZN (n_176), .A1 (n_91), .A2 (n_87), .A3 (n_89));
NOR4_X1 i_205 (.ZN (n_98), .A1 (n_106), .A2 (n_103), .A3 (n_102), .A4 (n_99));
NOR2_X1 i_204 (.ZN (n_175), .A1 (n_98), .A2 (n_84));
NAND2_X1 i_203 (.ZN (n_174), .A1 (n_176), .A2 (n_175));
NAND2_X1 i_196 (.ZN (n_81), .A1 (p_0[20]), .A2 (Accumulator[20]));
NAND2_X1 i_130 (.ZN (n_80), .A1 (p_0[21]), .A2 (Accumulator[21]));
NAND2_X1 i_129 (.ZN (n_173), .A1 (n_80), .A2 (n_81));
NAND2_X1 i_128 (.ZN (n_172), .A1 (n_176), .A2 (n_173));
NAND2_X1 i_127 (.ZN (n_171), .A1 (p_0[23]), .A2 (Accumulator[23]));
NAND2_X1 i_126 (.ZN (n_164), .A1 (p_0[22]), .A2 (Accumulator[22]));
INV_X1 i_125 (.ZN (n_77), .A (n_164));
OAI21_X1 i_124 (.ZN (n_97), .A (n_77), .B1 (p_0[23]), .B2 (Accumulator[23]));
NAND4_X1 i_123 (.ZN (n_52), .A1 (n_174), .A2 (n_172), .A3 (n_171), .A4 (n_97));
OAI21_X1 i_122 (.ZN (n_96), .A (n_52), .B1 (p_0[24]), .B2 (Accumulator[24]));
NAND2_X1 i_120 (.ZN (n_95), .A1 (p_0[25]), .A2 (Accumulator[25]));
NAND2_X1 i_118 (.ZN (n_94), .A1 (n_95), .A2 (n_74));
NAND3_X1 i_117 (.ZN (n_93), .A1 (n_182), .A2 (n_178), .A3 (n_94));
NAND2_X1 i_115 (.ZN (n_92), .A1 (p_0[26]), .A2 (Accumulator[26]));
OAI22_X1 i_114 (.ZN (n_90), .A1 (n_183), .A2 (n_92), .B1 (n_169), .B2 (n_166));
INV_X1 i_113 (.ZN (n_85), .A (n_90));
OAI211_X1 i_112 (.ZN (n_83), .A (n_93), .B (n_85), .C1 (n_177), .C2 (n_96));
INV_X1 i_110 (.ZN (n_66), .A (n_83));
OAI21_X1 i_109 (.ZN (n_64), .A (n_185), .B1 (n_66), .B2 (n_184));
NAND2_X1 i_108 (.ZN (n_82), .A1 (n_60), .A2 (n_64));
NAND2_X1 i_107 (.ZN (n_78), .A1 (p_0[30]), .A2 (Accumulator[30]));
AND2_X1 i_105 (.ZN (n_76), .A1 (n_82), .A2 (n_78));
NAND2_X1 i_104 (.ZN (n_75), .A1 (n_186), .A2 (n_76));
NAND3_X1 i_103 (.ZN (n_73), .A1 (n_75), .A2 (n_188), .A3 (n_187));
NAND2_X1 i_102 (.ZN (n_72), .A1 (n_75), .A2 (n_187));
NAND2_X1 i_101 (.ZN (n_71), .A1 (n_72), .A2 (p_0[31]));
NAND2_X1 i_100 (.ZN (Accumulator1[31]), .A1 (n_71), .A2 (n_73));
NAND2_X1 i_99 (.ZN (n_70), .A1 (n_187), .A2 (n_78));
NAND2_X1 i_98 (.ZN (n_69), .A1 (p_0[29]), .A2 (Accumulator[29]));
NAND2_X1 i_97 (.ZN (n_68), .A1 (n_82), .A2 (n_69));
XOR2_X1 i_96 (.Z (n_67), .A (n_70), .B (n_68));
INV_X1 i_95 (.ZN (Accumulator1[30]), .A (n_67));
NAND2_X1 i_94 (.ZN (n_62), .A1 (p_0[27]), .A2 (Accumulator[27]));
NAND2_X1 i_93 (.ZN (n_61), .A1 (n_182), .A2 (n_62));
INV_X1 i_92 (.ZN (n_57), .A (n_179));
INV_X1 i_90 (.ZN (n_56), .A (n_92));
NAND2_X1 i_89 (.ZN (n_55), .A1 (n_181), .A2 (n_180));
NOR2_X1 i_88 (.ZN (n_54), .A1 (p_0[24]), .A2 (Accumulator[24]));
OAI21_X1 i_87 (.ZN (n_53), .A (n_96), .B1 (n_74), .B2 (n_54));
NAND2_X1 i_86 (.ZN (n_50), .A1 (n_53), .A2 (n_55));
NAND2_X1 i_85 (.ZN (n_49), .A1 (n_50), .A2 (n_95));
OAI21_X1 i_84 (.ZN (n_48), .A (n_57), .B1 (n_49), .B2 (n_56));
XOR2_X1 i_81 (.Z (Accumulator1[27]), .A (n_61), .B (n_48));
NAND2_X1 i_80 (.ZN (n_47), .A1 (n_57), .A2 (n_92));
XNOR2_X1 i_78 (.ZN (Accumulator1[26]), .A (n_49), .B (n_47));
NAND2_X1 i_77 (.ZN (n_46), .A1 (n_55), .A2 (n_95));
XNOR2_X1 i_76 (.ZN (Accumulator1[25]), .A (n_46), .B (n_53));
INV_X1 i_75 (.ZN (n_86), .A (n_87));
INV_X1 i_74 (.ZN (n_88), .A (n_89));
INV_X1 i_73 (.ZN (n_45), .A (n_184));
NAND2_X1 i_72 (.ZN (n_44), .A1 (n_45), .A2 (n_185));
INV_X1 i_71 (.ZN (n_65), .A (n_44));
INV_X1 i_70 (.ZN (n_63), .A (n_64));
INV_X1 i_69 (.ZN (n_58), .A (n_59));
INV_X1 i_202 (.ZN (n_170), .A (p_0[29]));
INV_X1 i_201 (.ZN (n_169), .A (p_0[27]));
INV_X1 i_200 (.ZN (n_168), .A (p_0[3]));
INV_X1 i_199 (.ZN (n_167), .A (Accumulator[29]));
INV_X1 i_198 (.ZN (n_166), .A (Accumulator[27]));
INV_X1 i_197 (.ZN (n_165), .A (Accumulator[3]));
NAND2_X1 i_195 (.ZN (n_163), .A1 (n_168), .A2 (n_165));
NAND2_X1 i_194 (.ZN (n_162), .A1 (p_0[2]), .A2 (Accumulator[2]));
INV_X1 i_193 (.ZN (n_161), .A (n_162));
NOR2_X1 i_192 (.ZN (n_160), .A1 (p_0[1]), .A2 (Accumulator[1]));
NAND2_X1 i_191 (.ZN (n_159), .A1 (p_0[0]), .A2 (Accumulator[0]));
NAND2_X1 i_190 (.ZN (n_158), .A1 (p_0[1]), .A2 (Accumulator[1]));
AOI21_X1 i_189 (.ZN (n_157), .A (n_160), .B1 (n_159), .B2 (n_158));
OAI22_X1 i_188 (.ZN (n_156), .A1 (p_0[2]), .A2 (Accumulator[2]), .B1 (n_161), .B2 (n_157));
OAI21_X1 i_187 (.ZN (n_155), .A (n_156), .B1 (n_168), .B2 (n_165));
NAND2_X1 i_186 (.ZN (n_154), .A1 (n_163), .A2 (n_155));
NOR2_X1 i_185 (.ZN (n_153), .A1 (p_0[7]), .A2 (Accumulator[7]));
NOR2_X1 i_184 (.ZN (n_152), .A1 (p_0[5]), .A2 (Accumulator[5]));
NOR2_X1 i_183 (.ZN (n_151), .A1 (p_0[6]), .A2 (Accumulator[6]));
OR3_X1 i_182 (.ZN (n_150), .A1 (n_153), .A2 (n_151), .A3 (n_152));
NOR2_X1 i_181 (.ZN (n_149), .A1 (p_0[4]), .A2 (Accumulator[4]));
NOR3_X1 i_180 (.ZN (n_148), .A1 (n_150), .A2 (n_149), .A3 (n_154));
NAND2_X1 i_179 (.ZN (n_147), .A1 (p_0[4]), .A2 (Accumulator[4]));
NAND2_X1 i_178 (.ZN (n_146), .A1 (p_0[5]), .A2 (Accumulator[5]));
AOI21_X1 i_177 (.ZN (n_145), .A (n_150), .B1 (n_147), .B2 (n_146));
AND2_X1 i_176 (.ZN (n_144), .A1 (p_0[7]), .A2 (Accumulator[7]));
NAND2_X1 i_175 (.ZN (n_143), .A1 (p_0[6]), .A2 (Accumulator[6]));
INV_X1 i_174 (.ZN (n_142), .A (n_143));
NOR2_X1 i_173 (.ZN (n_141), .A1 (n_153), .A2 (n_143));
NOR4_X1 i_172 (.ZN (n_140), .A1 (n_144), .A2 (n_141), .A3 (n_145), .A4 (n_148));
NOR2_X1 i_171 (.ZN (n_139), .A1 (p_0[11]), .A2 (Accumulator[11]));
NOR2_X1 i_170 (.ZN (n_138), .A1 (p_0[9]), .A2 (Accumulator[9]));
NOR2_X1 i_169 (.ZN (n_137), .A1 (p_0[10]), .A2 (Accumulator[10]));
OR3_X1 i_168 (.ZN (n_136), .A1 (n_139), .A2 (n_137), .A3 (n_138));
NOR2_X1 i_167 (.ZN (n_135), .A1 (p_0[8]), .A2 (Accumulator[8]));
NOR3_X1 i_166 (.ZN (n_134), .A1 (n_136), .A2 (n_135), .A3 (n_140));
NAND2_X1 i_165 (.ZN (n_133), .A1 (p_0[8]), .A2 (Accumulator[8]));
NAND2_X1 i_164 (.ZN (n_132), .A1 (p_0[9]), .A2 (Accumulator[9]));
AOI21_X1 i_163 (.ZN (n_131), .A (n_136), .B1 (n_133), .B2 (n_132));
AND2_X1 i_162 (.ZN (n_130), .A1 (p_0[11]), .A2 (Accumulator[11]));
NAND2_X1 i_161 (.ZN (n_129), .A1 (p_0[10]), .A2 (Accumulator[10]));
INV_X1 i_160 (.ZN (n_128), .A (n_129));
NOR2_X1 i_159 (.ZN (n_127), .A1 (n_139), .A2 (n_129));
NOR4_X1 i_158 (.ZN (n_126), .A1 (n_130), .A2 (n_127), .A3 (n_131), .A4 (n_134));
NOR2_X1 i_157 (.ZN (n_125), .A1 (p_0[15]), .A2 (Accumulator[15]));
NOR2_X1 i_156 (.ZN (n_124), .A1 (p_0[13]), .A2 (Accumulator[13]));
NOR2_X1 i_155 (.ZN (n_123), .A1 (p_0[14]), .A2 (Accumulator[14]));
OR3_X1 i_154 (.ZN (n_122), .A1 (n_125), .A2 (n_123), .A3 (n_124));
NOR2_X1 i_153 (.ZN (n_121), .A1 (p_0[12]), .A2 (Accumulator[12]));
NOR3_X1 i_152 (.ZN (n_120), .A1 (n_122), .A2 (n_121), .A3 (n_126));
NAND2_X1 i_151 (.ZN (n_119), .A1 (p_0[12]), .A2 (Accumulator[12]));
NAND2_X1 i_150 (.ZN (n_118), .A1 (p_0[13]), .A2 (Accumulator[13]));
AOI21_X1 i_149 (.ZN (n_117), .A (n_122), .B1 (n_119), .B2 (n_118));
AND2_X1 i_148 (.ZN (n_116), .A1 (p_0[15]), .A2 (Accumulator[15]));
NAND2_X1 i_147 (.ZN (n_115), .A1 (p_0[14]), .A2 (Accumulator[14]));
INV_X1 i_146 (.ZN (n_114), .A (n_115));
NOR2_X1 i_145 (.ZN (n_113), .A1 (n_125), .A2 (n_115));
NOR4_X1 i_144 (.ZN (n_112), .A1 (n_116), .A2 (n_113), .A3 (n_117), .A4 (n_120));
NOR2_X1 i_143 (.ZN (n_111), .A1 (p_0[19]), .A2 (Accumulator[19]));
NOR2_X1 i_142 (.ZN (n_110), .A1 (p_0[17]), .A2 (Accumulator[17]));
NOR2_X1 i_141 (.ZN (n_109), .A1 (p_0[18]), .A2 (Accumulator[18]));
OR3_X1 i_140 (.ZN (n_108), .A1 (n_111), .A2 (n_109), .A3 (n_110));
NOR2_X1 i_139 (.ZN (n_107), .A1 (p_0[16]), .A2 (Accumulator[16]));
NOR3_X1 i_138 (.ZN (n_106), .A1 (n_108), .A2 (n_107), .A3 (n_112));
NAND2_X1 i_137 (.ZN (n_105), .A1 (p_0[16]), .A2 (Accumulator[16]));
NAND2_X1 i_136 (.ZN (n_104), .A1 (p_0[17]), .A2 (Accumulator[17]));
AOI21_X1 i_135 (.ZN (n_103), .A (n_108), .B1 (n_105), .B2 (n_104));
AND2_X1 i_134 (.ZN (n_102), .A1 (p_0[19]), .A2 (Accumulator[19]));
NAND2_X1 i_133 (.ZN (n_101), .A1 (p_0[18]), .A2 (Accumulator[18]));
INV_X1 i_132 (.ZN (n_100), .A (n_101));
NOR2_X1 i_131 (.ZN (n_99), .A1 (n_111), .A2 (n_101));
NOR2_X1 i_121 (.ZN (n_89), .A1 (p_0[21]), .A2 (Accumulator[21]));
NOR2_X1 i_119 (.ZN (n_87), .A1 (p_0[22]), .A2 (Accumulator[22]));
NOR2_X1 i_116 (.ZN (n_84), .A1 (p_0[20]), .A2 (Accumulator[20]));
INV_X1 i_111 (.ZN (n_79), .A (n_80));
NAND2_X1 i_106 (.ZN (n_74), .A1 (p_0[24]), .A2 (Accumulator[24]));
OAI21_X1 i_91 (.ZN (n_59), .A (n_60), .B1 (n_170), .B2 (n_167));
AOI22_X1 i_83 (.ZN (Accumulator1[29]), .A1 (n_63), .A2 (n_59), .B1 (n_64), .B2 (n_58));
XNOR2_X1 i_82 (.ZN (Accumulator1[28]), .A (n_66), .B (n_65));
OAI21_X1 i_79 (.ZN (n_51), .A (n_74), .B1 (p_0[24]), .B2 (Accumulator[24]));
XNOR2_X1 i_68 (.ZN (Accumulator1[24]), .A (n_52), .B (n_51));
AOI21_X1 i_67 (.ZN (n_43), .A (n_91), .B1 (p_0[23]), .B2 (Accumulator[23]));
OAI21_X1 i_66 (.ZN (n_42), .A (n_81), .B1 (p_0[20]), .B2 (Accumulator[20]));
AOI21_X1 i_65 (.ZN (n_41), .A (n_84), .B1 (n_98), .B2 (n_81));
OAI21_X1 i_64 (.ZN (n_40), .A (n_88), .B1 (n_79), .B2 (n_41));
INV_X1 i_63 (.ZN (n_39), .A (n_40));
NOR2_X1 i_62 (.ZN (n_38), .A1 (n_89), .A2 (n_79));
OAI21_X1 i_61 (.ZN (n_37), .A (n_86), .B1 (n_77), .B2 (n_39));
XNOR2_X1 i_60 (.ZN (Accumulator1[23]), .A (n_43), .B (n_37));
NOR2_X1 i_59 (.ZN (n_36), .A1 (n_87), .A2 (n_77));
XOR2_X1 i_58 (.Z (Accumulator1[22]), .A (n_39), .B (n_36));
XOR2_X1 i_57 (.Z (Accumulator1[21]), .A (n_41), .B (n_38));
XOR2_X1 i_56 (.Z (Accumulator1[20]), .A (n_98), .B (n_42));
NOR2_X1 i_55 (.ZN (n_35), .A1 (n_111), .A2 (n_102));
OAI21_X1 i_54 (.ZN (n_34), .A (n_105), .B1 (p_0[16]), .B2 (Accumulator[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_107), .B1 (n_112), .B2 (n_105));
INV_X1 i_52 (.ZN (n_32), .A (n_33));
AOI21_X1 i_51 (.ZN (n_31), .A (n_110), .B1 (n_104), .B2 (n_32));
AOI21_X1 i_50 (.ZN (n_30), .A (n_110), .B1 (p_0[17]), .B2 (Accumulator[17]));
OAI22_X1 i_49 (.ZN (n_29), .A1 (p_0[18]), .A2 (Accumulator[18]), .B1 (n_100), .B2 (n_31));
XNOR2_X1 i_48 (.ZN (Accumulator1[19]), .A (n_35), .B (n_29));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_109), .A2 (n_100));
XOR2_X1 i_46 (.Z (Accumulator1[18]), .A (n_31), .B (n_28));
XOR2_X1 i_45 (.Z (Accumulator1[17]), .A (n_33), .B (n_30));
XOR2_X1 i_44 (.Z (Accumulator1[16]), .A (n_112), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_125), .A2 (n_116));
OAI21_X1 i_42 (.ZN (n_26), .A (n_119), .B1 (p_0[12]), .B2 (Accumulator[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_121), .B1 (n_126), .B2 (n_119));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_124), .B1 (n_118), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_124), .B1 (p_0[13]), .B2 (Accumulator[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (p_0[14]), .A2 (Accumulator[14]), .B1 (n_114), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (Accumulator1[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_123), .A2 (n_114));
XOR2_X1 i_34 (.Z (Accumulator1[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (Accumulator1[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (Accumulator1[12]), .A (n_126), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_139), .A2 (n_130));
AOI21_X1 i_30 (.ZN (n_18), .A (n_135), .B1 (p_0[8]), .B2 (Accumulator[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_135), .B1 (n_140), .B2 (n_133));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_138), .B1 (n_132), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_138), .B1 (p_0[9]), .B2 (Accumulator[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (p_0[10]), .A2 (Accumulator[10]), .B1 (n_128), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (Accumulator1[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_137), .A2 (n_128));
XOR2_X1 i_22 (.Z (Accumulator1[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (Accumulator1[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (Accumulator1[8]), .A (n_140), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_153), .A2 (n_144));
OAI21_X1 i_18 (.ZN (n_10), .A (n_147), .B1 (p_0[4]), .B2 (Accumulator[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_149), .B1 (n_154), .B2 (n_147));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_152), .B1 (n_146), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_152), .B1 (p_0[5]), .B2 (Accumulator[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (p_0[6]), .A2 (Accumulator[6]), .B1 (n_142), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (Accumulator1[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_151), .A2 (n_142));
XOR2_X1 i_10 (.Z (Accumulator1[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (Accumulator1[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (Accumulator1[4]), .A (n_154), .B (n_10));
OAI21_X1 i_7 (.ZN (n_3), .A (n_163), .B1 (n_168), .B2 (n_165));
XOR2_X1 i_6 (.Z (Accumulator1[3]), .A (n_156), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_162), .B1 (p_0[2]), .B2 (Accumulator[2]));
XNOR2_X1 i_4 (.ZN (Accumulator1[2]), .A (n_157), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_158), .B1 (p_0[1]), .B2 (Accumulator[1]));
XOR2_X1 i_2 (.Z (Accumulator1[1]), .A (n_159), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_159), .B1 (p_0[0]), .B2 (Accumulator[0]));
INV_X1 i_0 (.ZN (Accumulator1[0]), .A (n_0));

endmodule //datapath__0_6

module datapath__0_2 (b, p_0);

output [31:0] p_0;
input [31:0] b;
wire n_19;
wire n_45;
wire n_18;
wire n_48;
wire n_46;
wire n_25;
wire n_44;
wire n_27;
wire n_24;
wire n_43;
wire n_26;
wire n_41;
wire n_42;
wire n_29;
wire n_40;
wire n_28;
wire n_30;
wire n_63;
wire n_32;
wire n_39;
wire n_31;
wire n_47;
wire n_34;
wire n_38;
wire n_36;
wire n_33;
wire n_37;
wire n_35;
wire n_4;
wire n_52;
wire n_0;
wire n_5;
wire n_1;
wire n_17;
wire n_50;
wire n_2;
wire n_61;
wire n_72;
wire n_6;
wire n_11;
wire n_7;
wire n_8;
wire n_10;
wire n_92;
wire n_94;
wire n_93;
wire n_12;
wire n_90;
wire n_13;
wire n_14;
wire n_16;
wire n_89;
wire n_86;
wire n_49;
wire n_81;
wire n_23;
wire n_85;
wire n_82;
wire n_77;
wire n_51;
wire n_53;
wire n_78;
wire n_56;
wire n_55;
wire n_74;
wire n_80;
wire n_57;
wire n_79;
wire n_58;
wire n_59;
wire n_60;
wire n_73;
wire n_62;
wire n_64;
wire n_66;
wire n_97;
wire n_67;
wire n_68;
wire n_71;
wire n_69;
wire n_70;
wire n_98;
wire n_99;
wire n_75;
wire n_76;
wire n_83;
wire n_84;
wire n_88;
wire n_91;
wire n_96;
wire n_95;


INV_X1 i_130 (.ZN (n_99), .A (b[17]));
INV_X1 i_129 (.ZN (n_98), .A (b[16]));
INV_X1 i_128 (.ZN (n_97), .A (n_2));
INV_X1 i_127 (.ZN (n_96), .A (b[3]));
INV_X1 i_126 (.ZN (n_95), .A (b[2]));
INV_X1 i_125 (.ZN (n_94), .A (b[1]));
INV_X1 i_124 (.ZN (n_93), .A (b[0]));
NAND3_X1 i_123 (.ZN (n_92), .A1 (n_95), .A2 (n_94), .A3 (n_93));
INV_X1 i_122 (.ZN (n_91), .A (n_92));
NAND2_X1 i_121 (.ZN (n_90), .A1 (n_91), .A2 (n_96));
INV_X1 i_120 (.ZN (n_89), .A (n_90));
INV_X1 i_119 (.ZN (n_88), .A (b[6]));
INV_X1 i_117 (.ZN (n_86), .A (b[4]));
NAND3_X1 i_116 (.ZN (n_85), .A1 (n_88), .A2 (n_1), .A3 (n_86));
OR2_X1 i_115 (.ZN (n_84), .A1 (n_85), .A2 (b[7]));
INV_X1 i_114 (.ZN (n_83), .A (n_84));
NAND2_X1 i_113 (.ZN (n_82), .A1 (n_83), .A2 (n_89));
INV_X1 i_112 (.ZN (n_81), .A (n_82));
INV_X1 i_111 (.ZN (n_80), .A (b[11]));
INV_X1 i_110 (.ZN (n_79), .A (b[10]));
INV_X1 i_109 (.ZN (n_78), .A (b[9]));
INV_X1 i_108 (.ZN (n_77), .A (b[8]));
NAND4_X1 i_107 (.ZN (n_76), .A1 (n_80), .A2 (n_79), .A3 (n_78), .A4 (n_77));
INV_X1 i_106 (.ZN (n_75), .A (n_76));
NAND2_X1 i_105 (.ZN (n_74), .A1 (n_81), .A2 (n_75));
INV_X1 i_104 (.ZN (n_73), .A (n_74));
NAND4_X1 i_103 (.ZN (n_72), .A1 (n_97), .A2 (n_99), .A3 (n_98), .A4 (n_73));
NAND3_X1 i_102 (.ZN (n_71), .A1 (n_97), .A2 (n_98), .A3 (n_73));
NAND2_X1 i_101 (.ZN (n_70), .A1 (n_71), .A2 (b[17]));
NAND2_X1 i_100 (.ZN (n_69), .A1 (n_70), .A2 (n_72));
INV_X1 i_99 (.ZN (p_0[17]), .A (n_69));
NAND2_X1 i_98 (.ZN (n_48), .A1 (n_97), .A2 (n_73));
NAND2_X1 i_97 (.ZN (n_68), .A1 (n_48), .A2 (b[16]));
NAND2_X1 i_96 (.ZN (n_67), .A1 (n_68), .A2 (n_71));
INV_X1 i_95 (.ZN (p_0[16]), .A (n_67));
OR3_X1 i_93 (.ZN (n_50), .A1 (b[14]), .A2 (b[13]), .A3 (b[12]));
OR2_X1 i_92 (.ZN (n_66), .A1 (n_74), .A2 (n_50));
AOI22_X1 i_91 (.ZN (p_0[15]), .A1 (n_97), .A2 (n_73), .B1 (b[15]), .B2 (n_66));
INV_X1 i_89 (.ZN (n_64), .A (n_66));
AOI21_X1 i_88 (.ZN (p_0[14]), .A (n_64), .B1 (n_4), .B2 (b[14]));
INV_X1 i_87 (.ZN (n_62), .A (b[12]));
NAND2_X1 i_86 (.ZN (n_61), .A1 (n_73), .A2 (n_62));
XNOR2_X1 i_85 (.ZN (n_60), .A (n_61), .B (b[13]));
INV_X1 i_84 (.ZN (p_0[13]), .A (n_60));
NAND2_X1 i_83 (.ZN (n_59), .A1 (n_74), .A2 (b[12]));
NAND2_X1 i_82 (.ZN (n_58), .A1 (n_61), .A2 (n_59));
INV_X1 i_81 (.ZN (p_0[12]), .A (n_58));
NAND4_X1 i_80 (.ZN (n_57), .A1 (n_81), .A2 (n_79), .A3 (n_78), .A4 (n_77));
INV_X1 i_79 (.ZN (n_56), .A (n_57));
OAI21_X1 i_42 (.ZN (n_55), .A (n_74), .B1 (n_56), .B2 (n_80));
INV_X1 i_41 (.ZN (p_0[11]), .A (n_55));
AOI21_X1 i_34 (.ZN (p_0[10]), .A (n_56), .B1 (n_52), .B2 (b[10]));
OAI21_X1 i_33 (.ZN (n_53), .A (b[9]), .B1 (n_82), .B2 (b[8]));
NAND3_X1 i_32 (.ZN (n_52), .A1 (n_81), .A2 (n_78), .A3 (n_77));
NAND2_X1 i_31 (.ZN (n_51), .A1 (n_53), .A2 (n_52));
INV_X1 i_30 (.ZN (p_0[9]), .A (n_51));
XNOR2_X1 i_29 (.ZN (p_0[8]), .A (n_82), .B (n_77));
INV_X1 i_28 (.ZN (n_49), .A (n_85));
NAND2_X1 i_27 (.ZN (n_23), .A1 (n_89), .A2 (n_49));
AOI21_X1 i_26 (.ZN (p_0[7]), .A (n_81), .B1 (b[7]), .B2 (n_23));
AOI22_X1 i_24 (.ZN (p_0[6]), .A1 (n_0), .A2 (b[6]), .B1 (n_89), .B2 (n_49));
NAND2_X1 i_23 (.ZN (n_17), .A1 (n_89), .A2 (n_86));
NAND2_X1 i_22 (.ZN (n_16), .A1 (n_90), .A2 (b[4]));
NAND2_X1 i_21 (.ZN (n_14), .A1 (n_17), .A2 (n_16));
INV_X1 i_20 (.ZN (p_0[4]), .A (n_14));
NAND2_X1 i_19 (.ZN (n_13), .A1 (n_92), .A2 (b[3]));
NAND2_X1 i_18 (.ZN (n_12), .A1 (n_90), .A2 (n_13));
INV_X1 i_17 (.ZN (p_0[3]), .A (n_12));
NAND2_X1 i_16 (.ZN (n_11), .A1 (n_94), .A2 (n_93));
NAND2_X1 i_15 (.ZN (n_10), .A1 (n_11), .A2 (b[2]));
NAND2_X1 i_14 (.ZN (n_8), .A1 (n_10), .A2 (n_92));
INV_X1 i_13 (.ZN (p_0[2]), .A (n_8));
NAND2_X1 i_12 (.ZN (n_7), .A1 (b[1]), .A2 (b[0]));
NAND2_X1 i_11 (.ZN (n_6), .A1 (n_11), .A2 (n_7));
INV_X1 i_10 (.ZN (p_0[1]), .A (n_6));
INV_X1 i_9 (.ZN (n_5), .A (n_17));
OR2_X1 i_7 (.ZN (n_4), .A1 (n_61), .A2 (b[13]));
OR2_X1 i_6 (.ZN (n_2), .A1 (n_50), .A2 (b[15]));
INV_X1 i_5 (.ZN (n_1), .A (b[5]));
XNOR2_X1 i_4 (.ZN (p_0[5]), .A (n_17), .B (n_1));
NAND2_X1 i_3 (.ZN (n_0), .A1 (n_5), .A2 (n_1));
INV_X1 i_94 (.ZN (n_63), .A (b[25]));
OR3_X1 i_78 (.ZN (n_47), .A1 (b[26]), .A2 (b[25]), .A3 (b[24]));
OR3_X1 i_77 (.ZN (n_46), .A1 (b[18]), .A2 (b[16]), .A3 (b[17]));
NOR3_X1 i_76 (.ZN (n_45), .A1 (b[19]), .A2 (n_46), .A3 (n_48));
INV_X1 i_75 (.ZN (n_44), .A (n_45));
NOR4_X1 i_74 (.ZN (n_43), .A1 (b[22]), .A2 (b[21]), .A3 (b[20]), .A4 (n_44));
INV_X1 i_73 (.ZN (n_42), .A (n_43));
NOR2_X1 i_72 (.ZN (n_41), .A1 (b[23]), .A2 (n_42));
INV_X1 i_71 (.ZN (n_40), .A (n_41));
NOR3_X1 i_70 (.ZN (n_39), .A1 (b[27]), .A2 (n_47), .A3 (n_40));
INV_X1 i_69 (.ZN (n_38), .A (n_39));
NOR4_X1 i_68 (.ZN (n_37), .A1 (b[29]), .A2 (b[28]), .A3 (b[30]), .A4 (n_38));
XNOR2_X1 i_67 (.ZN (p_0[31]), .A (b[31]), .B (n_37));
NOR3_X1 i_66 (.ZN (n_36), .A1 (b[29]), .A2 (b[28]), .A3 (n_38));
INV_X1 i_65 (.ZN (n_35), .A (n_36));
AOI21_X1 i_64 (.ZN (p_0[30]), .A (n_37), .B1 (b[30]), .B2 (n_35));
NOR2_X1 i_63 (.ZN (n_34), .A1 (b[28]), .A2 (n_38));
INV_X1 i_62 (.ZN (n_33), .A (n_34));
AOI21_X1 i_61 (.ZN (p_0[29]), .A (n_36), .B1 (b[29]), .B2 (n_33));
AOI21_X1 i_60 (.ZN (p_0[28]), .A (n_34), .B1 (b[28]), .B2 (n_38));
NOR2_X1 i_59 (.ZN (n_32), .A1 (n_47), .A2 (n_40));
INV_X1 i_58 (.ZN (n_31), .A (n_32));
AOI21_X1 i_57 (.ZN (p_0[27]), .A (n_39), .B1 (b[27]), .B2 (n_31));
OR3_X1 i_56 (.ZN (n_30), .A1 (b[25]), .A2 (b[24]), .A3 (n_40));
AOI21_X1 i_55 (.ZN (p_0[26]), .A (n_32), .B1 (b[26]), .B2 (n_30));
NOR2_X1 i_54 (.ZN (n_29), .A1 (b[24]), .A2 (n_40));
OAI21_X1 i_53 (.ZN (n_28), .A (n_30), .B1 (n_63), .B2 (n_29));
INV_X1 i_52 (.ZN (p_0[25]), .A (n_28));
AOI21_X1 i_51 (.ZN (p_0[24]), .A (n_29), .B1 (b[24]), .B2 (n_40));
AOI21_X1 i_50 (.ZN (p_0[23]), .A (n_41), .B1 (b[23]), .B2 (n_42));
NOR3_X1 i_49 (.ZN (n_27), .A1 (b[21]), .A2 (b[20]), .A3 (n_44));
INV_X1 i_48 (.ZN (n_26), .A (n_27));
AOI21_X1 i_47 (.ZN (p_0[22]), .A (n_43), .B1 (b[22]), .B2 (n_26));
NOR2_X1 i_46 (.ZN (n_25), .A1 (b[20]), .A2 (n_44));
INV_X1 i_45 (.ZN (n_24), .A (n_25));
AOI21_X1 i_44 (.ZN (p_0[21]), .A (n_27), .B1 (b[21]), .B2 (n_24));
AOI21_X1 i_43 (.ZN (p_0[20]), .A (n_25), .B1 (b[20]), .B2 (n_44));
NOR2_X1 i_38 (.ZN (n_19), .A1 (n_48), .A2 (n_46));
INV_X1 i_37 (.ZN (n_18), .A (n_19));
AOI21_X1 i_36 (.ZN (p_0[19]), .A (n_45), .B1 (b[19]), .B2 (n_18));
AOI21_X1 i_35 (.ZN (p_0[18]), .A (n_19), .B1 (b[18]), .B2 (n_72));

endmodule //datapath__0_2

module datapath (a, p_0);

output [31:0] p_0;
input [31:0] a;
wire n_62;
wire n_60;
wire n_61;
wire n_58;
wire n_59;
wire n_5;
wire n_57;
wire n_3;
wire n_4;
wire n_1;
wire n_2;
wire n_55;
wire n_0;
wire n_56;
wire n_11;
wire n_54;
wire n_9;
wire n_10;
wire n_7;
wire n_8;
wire n_52;
wire n_6;
wire n_53;
wire n_17;
wire n_51;
wire n_15;
wire n_16;
wire n_13;
wire n_14;
wire n_49;
wire n_12;
wire n_50;
wire n_23;
wire n_48;
wire n_21;
wire n_22;
wire n_19;
wire n_20;
wire n_45;
wire n_18;
wire n_46;
wire n_25;
wire n_44;
wire n_27;
wire n_24;
wire n_43;
wire n_26;
wire n_41;
wire n_42;
wire n_29;
wire n_40;
wire n_36;
wire n_34;
wire n_37;
wire n_35;
wire n_38;
wire n_28;
wire n_81;
wire n_80;
wire n_79;
wire n_87;
wire n_86;
wire n_85;
wire n_93;
wire n_92;
wire n_91;
wire n_99;
wire n_98;
wire n_97;
wire n_103;
wire n_102;
wire n_101;
wire n_31;
wire n_30;
wire n_32;
wire n_69;
wire n_105;
wire n_72;
wire n_39;
wire n_47;
wire n_89;
wire n_83;
wire n_77;
wire n_95;
wire n_64;
wire n_63;
wire n_67;
wire n_65;
wire n_106;
wire n_66;
wire n_68;
wire n_71;
wire n_70;
wire n_73;
wire n_76;
wire n_75;
wire n_74;
wire n_78;
wire n_82;
wire n_84;
wire n_88;
wire n_90;
wire n_94;
wire n_96;
wire n_100;
wire n_104;


INV_X1 i_137 (.ZN (n_106), .A (a[28]));
INV_X1 i_136 (.ZN (n_105), .A (a[23]));
INV_X1 i_135 (.ZN (n_104), .A (a[3]));
INV_X1 i_134 (.ZN (n_103), .A (a[2]));
INV_X1 i_133 (.ZN (n_102), .A (a[1]));
INV_X1 i_132 (.ZN (n_101), .A (a[0]));
NAND4_X1 i_131 (.ZN (n_57), .A1 (n_104), .A2 (n_103), .A3 (n_102), .A4 (n_101));
INV_X1 i_130 (.ZN (n_58), .A (n_57));
INV_X1 i_129 (.ZN (n_100), .A (a[7]));
INV_X1 i_128 (.ZN (n_99), .A (a[6]));
INV_X1 i_127 (.ZN (n_98), .A (a[5]));
INV_X1 i_126 (.ZN (n_97), .A (a[4]));
NAND4_X1 i_125 (.ZN (n_96), .A1 (n_100), .A2 (n_99), .A3 (n_98), .A4 (n_97));
INV_X1 i_124 (.ZN (n_95), .A (n_96));
INV_X1 i_123 (.ZN (n_94), .A (a[11]));
INV_X1 i_122 (.ZN (n_93), .A (a[10]));
INV_X1 i_121 (.ZN (n_92), .A (a[9]));
INV_X1 i_120 (.ZN (n_91), .A (a[8]));
NAND4_X1 i_119 (.ZN (n_90), .A1 (n_94), .A2 (n_93), .A3 (n_92), .A4 (n_91));
INV_X1 i_118 (.ZN (n_89), .A (n_90));
NAND3_X1 i_117 (.ZN (n_51), .A1 (n_58), .A2 (n_95), .A3 (n_89));
INV_X1 i_116 (.ZN (n_52), .A (n_51));
INV_X1 i_115 (.ZN (n_88), .A (a[15]));
INV_X1 i_114 (.ZN (n_87), .A (a[14]));
INV_X1 i_113 (.ZN (n_86), .A (a[13]));
INV_X1 i_112 (.ZN (n_85), .A (a[12]));
NAND4_X1 i_111 (.ZN (n_84), .A1 (n_88), .A2 (n_87), .A3 (n_86), .A4 (n_85));
INV_X1 i_110 (.ZN (n_83), .A (n_84));
INV_X1 i_109 (.ZN (n_82), .A (a[19]));
INV_X1 i_108 (.ZN (n_81), .A (a[18]));
INV_X1 i_107 (.ZN (n_80), .A (a[17]));
INV_X1 i_106 (.ZN (n_79), .A (a[16]));
NAND4_X1 i_105 (.ZN (n_78), .A1 (n_82), .A2 (n_81), .A3 (n_80), .A4 (n_79));
INV_X1 i_104 (.ZN (n_77), .A (n_78));
INV_X1 i_103 (.ZN (n_76), .A (a[22]));
INV_X1 i_102 (.ZN (n_75), .A (a[21]));
INV_X1 i_101 (.ZN (n_74), .A (a[20]));
NAND3_X1 i_100 (.ZN (n_73), .A1 (n_76), .A2 (n_75), .A3 (n_74));
INV_X1 i_99 (.ZN (n_72), .A (n_73));
NAND4_X1 i_98 (.ZN (n_42), .A1 (n_52), .A2 (n_83), .A3 (n_77), .A4 (n_72));
INV_X1 i_97 (.ZN (n_43), .A (n_42));
INV_X1 i_96 (.ZN (n_71), .A (a[27]));
OR3_X1 i_95 (.ZN (n_70), .A1 (a[26]), .A2 (a[25]), .A3 (a[24]));
INV_X1 i_94 (.ZN (n_69), .A (n_70));
NAND2_X1 i_93 (.ZN (n_68), .A1 (n_69), .A2 (n_71));
INV_X1 i_92 (.ZN (n_67), .A (n_68));
NAND4_X1 i_91 (.ZN (n_66), .A1 (n_43), .A2 (n_106), .A3 (n_105), .A4 (n_67));
INV_X1 i_90 (.ZN (n_34), .A (n_66));
NAND4_X1 i_89 (.ZN (n_48), .A1 (n_58), .A2 (n_95), .A3 (n_89), .A4 (n_83));
INV_X1 i_88 (.ZN (n_49), .A (n_48));
NAND4_X1 i_87 (.ZN (n_40), .A1 (n_49), .A2 (n_105), .A3 (n_77), .A4 (n_72));
INV_X1 i_86 (.ZN (n_41), .A (n_40));
AOI21_X1 i_85 (.ZN (n_65), .A (n_106), .B1 (n_41), .B2 (n_67));
NOR2_X1 i_84 (.ZN (p_0[28]), .A1 (n_65), .A2 (n_34));
NAND3_X1 i_83 (.ZN (n_38), .A1 (n_43), .A2 (n_105), .A3 (n_67));
INV_X1 i_82 (.ZN (n_64), .A (n_38));
NAND2_X1 i_81 (.ZN (n_63), .A1 (n_41), .A2 (n_69));
AOI21_X1 i_80 (.ZN (p_0[27]), .A (n_64), .B1 (n_63), .B2 (a[27]));
NAND2_X1 i_79 (.ZN (n_54), .A1 (n_58), .A2 (n_95));
INV_X1 i_78 (.ZN (n_55), .A (n_54));
NAND4_X1 i_77 (.ZN (n_44), .A1 (n_55), .A2 (n_89), .A3 (n_83), .A4 (n_77));
INV_X1 i_76 (.ZN (n_45), .A (n_44));
OR2_X1 i_75 (.ZN (n_47), .A1 (a[25]), .A2 (a[24]));
INV_X1 i_74 (.ZN (n_39), .A (n_47));
NAND4_X1 i_73 (.ZN (n_32), .A1 (n_45), .A2 (n_105), .A3 (n_72), .A4 (n_39));
AOI22_X1 i_72 (.ZN (p_0[26]), .A1 (n_32), .A2 (a[26]), .B1 (n_41), .B2 (n_69));
INV_X1 i_71 (.ZN (n_31), .A (n_32));
INV_X1 i_70 (.ZN (n_30), .A (a[24]));
NAND2_X1 i_69 (.ZN (n_28), .A1 (n_41), .A2 (n_30));
AOI21_X1 i_63 (.ZN (p_0[25]), .A (n_31), .B1 (n_28), .B2 (a[25]));
NAND2_X1 i_60 (.ZN (n_61), .A1 (n_102), .A2 (n_101));
INV_X1 i_59 (.ZN (n_62), .A (n_61));
NAND2_X1 i_58 (.ZN (n_59), .A1 (n_62), .A2 (n_103));
INV_X1 i_57 (.ZN (n_60), .A (n_59));
NAND3_X1 i_56 (.ZN (n_56), .A1 (n_99), .A2 (n_98), .A3 (n_97));
NAND3_X1 i_55 (.ZN (n_53), .A1 (n_93), .A2 (n_92), .A3 (n_91));
NAND3_X1 i_54 (.ZN (n_50), .A1 (n_87), .A2 (n_86), .A3 (n_85));
NAND3_X1 i_53 (.ZN (n_46), .A1 (n_81), .A2 (n_80), .A3 (n_79));
INV_X1 i_52 (.ZN (n_29), .A (n_28));
NOR4_X2 i_68 (.ZN (n_37), .A1 (a[29]), .A2 (a[28]), .A3 (a[30]), .A4 (n_38));
XNOR2_X1 i_67 (.ZN (p_0[31]), .A (a[31]), .B (n_37));
NOR3_X1 i_66 (.ZN (n_36), .A1 (a[29]), .A2 (a[28]), .A3 (n_38));
INV_X1 i_65 (.ZN (n_35), .A (n_36));
AOI21_X1 i_64 (.ZN (p_0[30]), .A (n_37), .B1 (a[30]), .B2 (n_35));
AOI21_X1 i_61 (.ZN (p_0[29]), .A (n_36), .B1 (a[29]), .B2 (n_66));
AOI21_X1 i_51 (.ZN (p_0[24]), .A (n_29), .B1 (a[24]), .B2 (n_40));
AOI21_X1 i_50 (.ZN (p_0[23]), .A (n_41), .B1 (a[23]), .B2 (n_42));
NOR3_X1 i_49 (.ZN (n_27), .A1 (a[21]), .A2 (a[20]), .A3 (n_44));
INV_X1 i_48 (.ZN (n_26), .A (n_27));
AOI21_X1 i_47 (.ZN (p_0[22]), .A (n_43), .B1 (a[22]), .B2 (n_26));
NOR2_X1 i_46 (.ZN (n_25), .A1 (a[20]), .A2 (n_44));
INV_X1 i_45 (.ZN (n_24), .A (n_25));
AOI21_X1 i_44 (.ZN (p_0[21]), .A (n_27), .B1 (a[21]), .B2 (n_24));
AOI21_X1 i_43 (.ZN (p_0[20]), .A (n_25), .B1 (a[20]), .B2 (n_44));
NOR2_X1 i_42 (.ZN (n_23), .A1 (a[16]), .A2 (n_48));
INV_X1 i_41 (.ZN (n_22), .A (n_23));
NOR2_X1 i_40 (.ZN (n_21), .A1 (a[17]), .A2 (n_22));
INV_X1 i_39 (.ZN (n_20), .A (n_21));
NOR2_X1 i_38 (.ZN (n_19), .A1 (n_48), .A2 (n_46));
INV_X1 i_37 (.ZN (n_18), .A (n_19));
AOI21_X1 i_36 (.ZN (p_0[19]), .A (n_45), .B1 (a[19]), .B2 (n_18));
AOI21_X1 i_35 (.ZN (p_0[18]), .A (n_19), .B1 (a[18]), .B2 (n_20));
AOI21_X1 i_34 (.ZN (p_0[17]), .A (n_21), .B1 (a[17]), .B2 (n_22));
AOI21_X1 i_33 (.ZN (p_0[16]), .A (n_23), .B1 (a[16]), .B2 (n_48));
NOR2_X1 i_32 (.ZN (n_17), .A1 (a[12]), .A2 (n_51));
INV_X1 i_31 (.ZN (n_16), .A (n_17));
NOR2_X1 i_30 (.ZN (n_15), .A1 (a[13]), .A2 (n_16));
INV_X1 i_29 (.ZN (n_14), .A (n_15));
NOR2_X1 i_28 (.ZN (n_13), .A1 (n_51), .A2 (n_50));
INV_X1 i_27 (.ZN (n_12), .A (n_13));
AOI21_X1 i_26 (.ZN (p_0[15]), .A (n_49), .B1 (a[15]), .B2 (n_12));
AOI21_X1 i_25 (.ZN (p_0[14]), .A (n_13), .B1 (a[14]), .B2 (n_14));
AOI21_X1 i_24 (.ZN (p_0[13]), .A (n_15), .B1 (a[13]), .B2 (n_16));
AOI21_X1 i_23 (.ZN (p_0[12]), .A (n_17), .B1 (a[12]), .B2 (n_51));
NOR2_X1 i_22 (.ZN (n_11), .A1 (a[8]), .A2 (n_54));
INV_X1 i_21 (.ZN (n_10), .A (n_11));
NOR2_X1 i_20 (.ZN (n_9), .A1 (a[9]), .A2 (n_10));
INV_X1 i_19 (.ZN (n_8), .A (n_9));
NOR2_X1 i_18 (.ZN (n_7), .A1 (n_54), .A2 (n_53));
INV_X1 i_17 (.ZN (n_6), .A (n_7));
AOI21_X1 i_16 (.ZN (p_0[11]), .A (n_52), .B1 (a[11]), .B2 (n_6));
AOI21_X1 i_15 (.ZN (p_0[10]), .A (n_7), .B1 (a[10]), .B2 (n_8));
AOI21_X1 i_14 (.ZN (p_0[9]), .A (n_9), .B1 (a[9]), .B2 (n_10));
AOI21_X1 i_13 (.ZN (p_0[8]), .A (n_11), .B1 (a[8]), .B2 (n_54));
NOR2_X1 i_12 (.ZN (n_5), .A1 (a[4]), .A2 (n_57));
INV_X1 i_11 (.ZN (n_4), .A (n_5));
NOR2_X1 i_10 (.ZN (n_3), .A1 (a[5]), .A2 (n_4));
INV_X1 i_9 (.ZN (n_2), .A (n_3));
NOR2_X1 i_8 (.ZN (n_1), .A1 (n_57), .A2 (n_56));
INV_X1 i_7 (.ZN (n_0), .A (n_1));
AOI21_X1 i_6 (.ZN (p_0[7]), .A (n_55), .B1 (a[7]), .B2 (n_0));
AOI21_X1 i_5 (.ZN (p_0[6]), .A (n_1), .B1 (a[6]), .B2 (n_2));
AOI21_X1 i_4 (.ZN (p_0[5]), .A (n_3), .B1 (a[5]), .B2 (n_4));
AOI21_X1 i_3 (.ZN (p_0[4]), .A (n_5), .B1 (a[4]), .B2 (n_57));
AOI21_X1 i_2 (.ZN (p_0[3]), .A (n_58), .B1 (a[3]), .B2 (n_59));
AOI21_X1 i_1 (.ZN (p_0[2]), .A (n_60), .B1 (a[2]), .B2 (n_61));
AOI21_X1 i_0 (.ZN (p_0[1]), .A (n_62), .B1 (a[1]), .B2 (a[0]));

endmodule //datapath

module seq_multiplier (clk, rst, a, b, c);

output [63:0] c;
input [31:0] a;
input [31:0] b;
input clk;
input rst;
wire CTS_n_tid0_168;
wire CTS_n_tid1_120;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_0_5;
wire n_0_0_0;
wire n_0_0_6;
wire n_0_0_1;
wire n_0_0_7;
wire n_0_0_2;
wire n_0_0_8;
wire n_0_0_3;
wire n_0_0_9;
wire n_0_0_4;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_0_10;
wire n_0_166;
wire n_0_0_11;
wire n_0_167;
wire n_0_0_12;
wire n_0_168;
wire n_0_0_13;
wire n_0_169;
wire n_0_0_14;
wire n_0_170;
wire n_0_0_15;
wire n_0_171;
wire n_0_0_16;
wire n_0_172;
wire n_0_0_17;
wire n_0_173;
wire n_0_0_18;
wire n_0_174;
wire n_0_0_19;
wire n_0_175;
wire n_0_0_20;
wire n_0_176;
wire n_0_0_21;
wire n_0_177;
wire n_0_0_22;
wire n_0_178;
wire n_0_0_23;
wire n_0_179;
wire n_0_0_24;
wire n_0_180;
wire n_0_0_25;
wire n_0_181;
wire n_0_0_26;
wire n_0_182;
wire n_0_0_27;
wire n_0_183;
wire n_0_0_28;
wire n_0_184;
wire n_0_0_29;
wire n_0_185;
wire n_0_0_30;
wire n_0_186;
wire n_0_0_31;
wire n_0_187;
wire n_0_0_32;
wire n_0_188;
wire n_0_0_33;
wire n_0_189;
wire n_0_0_34;
wire n_0_190;
wire n_0_0_35;
wire n_0_191;
wire n_0_0_36;
wire n_0_192;
wire n_0_0_37;
wire n_0_193;
wire n_0_0_38;
wire n_0_194;
wire n_0_0_39;
wire n_0_195;
wire n_0_0_40;
wire n_0_196;
wire n_0_0_41;
wire n_0_197;
wire n_0_0_42;
wire n_0_198;
wire n_0_0_43;
wire n_0_199;
wire n_0_0_44;
wire n_0_200;
wire n_0_0_45;
wire n_0_201;
wire n_0_0_46;
wire n_0_202;
wire n_0_0_47;
wire n_0_203;
wire n_0_0_48;
wire n_0_204;
wire n_0_0_49;
wire n_0_205;
wire n_0_0_50;
wire n_0_206;
wire n_0_0_51;
wire n_0_207;
wire n_0_0_52;
wire n_0_208;
wire n_0_0_53;
wire n_0_209;
wire n_0_0_54;
wire n_0_210;
wire n_0_0_55;
wire n_0_211;
wire n_0_0_56;
wire n_0_212;
wire n_0_0_57;
wire n_0_213;
wire n_0_0_58;
wire n_0_214;
wire n_0_0_59;
wire n_0_215;
wire n_0_0_60;
wire n_0_216;
wire n_0_0_61;
wire n_0_217;
wire n_0_0_62;
wire n_0_218;
wire n_0_0_63;
wire n_0_219;
wire n_0_0_64;
wire n_0_220;
wire n_0_0_65;
wire n_0_221;
wire n_0_0_66;
wire n_0_222;
wire n_0_0_67;
wire n_0_223;
wire n_0_0_68;
wire n_0_224;
wire n_0_0_69;
wire n_0_228;
wire n_0_229;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_233;
wire n_0_234;
wire n_0_235;
wire n_0_236;
wire n_0_237;
wire n_0_238;
wire n_0_239;
wire n_0_240;
wire n_0_241;
wire n_0_242;
wire n_0_243;
wire n_0_244;
wire n_0_245;
wire n_0_246;
wire n_0_247;
wire n_0_248;
wire n_0_249;
wire n_0_250;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_257;
wire n_0_258;
wire n_0_259;
wire n_0_260;
wire n_0_261;
wire n_0_262;
wire n_0_263;
wire n_0_264;
wire n_0_265;
wire n_0_266;
wire n_0_267;
wire n_0_268;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_272;
wire n_0_273;
wire n_0_274;
wire n_0_275;
wire n_0_276;
wire n_0_277;
wire n_0_278;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_282;
wire n_0_283;
wire n_0_284;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_288;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_296;
wire n_0_297;
wire n_0_298;
wire n_0_299;
wire n_0_300;
wire n_0_301;
wire n_0_302;
wire n_0_303;
wire n_0_304;
wire n_0_305;
wire n_0_306;
wire n_0_307;
wire n_0_308;
wire n_0_309;
wire n_0_310;
wire n_0_311;
wire n_0_312;
wire n_0_313;
wire n_0_314;
wire n_0_315;
wire n_0_316;
wire n_0_317;
wire n_0_318;
wire n_0_319;
wire n_0_320;
wire n_0_321;
wire n_0_322;
wire n_0_323;
wire n_0_324;
wire n_0_325;
wire n_0_326;
wire n_0_327;
wire n_0_328;
wire n_0_329;
wire n_0_330;
wire n_0_331;
wire n_0_332;
wire n_0_333;
wire n_0_334;
wire n_0_335;
wire n_0_336;
wire n_0_337;
wire n_0_338;
wire n_0_339;
wire n_0_340;
wire n_0_341;
wire n_0_342;
wire n_0_343;
wire n_0_344;
wire n_0_345;
wire n_0_346;
wire n_0_347;
wire n_0_348;
wire n_0_349;
wire n_0_350;
wire n_0_351;
wire n_0_352;
wire n_0_353;
wire n_0_354;
wire n_0_0_75;
wire n_0_355;
wire n_0_0_76;
wire n_0_357;
wire n_0_0_78;
wire n_0_358;
wire n_0_0_79;
wire n_0_359;
wire n_0_0_80;
wire n_0_360;
wire n_0_0_81;
wire n_0_367;
wire n_0_0_88;
wire n_0_368;
wire n_0_0_89;
wire n_0_369;
wire n_0_0_90;
wire n_0_370;
wire n_0_0_91;
wire n_0_371;
wire n_0_0_92;
wire n_0_372;
wire n_0_0_93;
wire n_0_373;
wire n_0_0_94;
wire n_0_374;
wire n_0_0_95;
wire n_0_375;
wire n_0_0_96;
wire n_0_376;
wire n_0_0_97;
wire n_0_377;
wire n_0_0_98;
wire n_0_378;
wire n_0_0_99;
wire n_0_379;
wire n_0_0_100;
wire n_0_380;
wire n_0_0_101;
wire n_0_381;
wire n_0_0_102;
wire n_0_382;
wire n_0_0_103;
wire n_0_383;
wire n_0_0_104;
wire n_0_384;
wire n_0_0_105;
wire n_0_385;
wire n_0_0_107;
wire n_0_386;
wire n_0_0_109;
wire n_0_387;
wire n_0_0_110;
wire n_0_388;
wire n_0_0_111;
wire n_0_389;
wire n_0_0_112;
wire n_0_390;
wire n_0_0_113;
wire n_0_391;
wire n_0_0_114;
wire n_0_392;
wire n_0_0_115;
wire n_0_393;
wire n_0_0_116;
wire n_0_394;
wire n_0_0_117;
wire n_0_395;
wire n_0_0_118;
wire n_0_396;
wire n_0_0_119;
wire n_0_397;
wire n_0_0_120;
wire n_0_398;
wire n_0_0_121;
wire n_0_399;
wire n_0_0_122;
wire n_0_400;
wire n_0_0_123;
wire n_0_401;
wire n_0_0_124;
wire n_0_402;
wire n_0_0_125;
wire n_0_403;
wire n_0_0_126;
wire n_0_404;
wire n_0_0_127;
wire n_0_405;
wire n_0_0_128;
wire n_0_406;
wire n_0_0_129;
wire n_0_407;
wire n_0_0_130;
wire n_0_408;
wire n_0_0_131;
wire n_0_409;
wire n_0_0_132;
wire n_0_410;
wire n_0_0_133;
wire n_0_411;
wire n_0_0_134;
wire n_0_412;
wire n_0_0_135;
wire n_0_413;
wire n_0_0_136;
wire n_0_414;
wire n_0_0_137;
wire n_0_415;
wire n_0_0_138;
wire n_0_416;
wire n_0_0_139;
wire n_0_0_140;
wire n_0_417;
wire n_0_0_141;
wire n_0_0_142;
wire n_0_0_143;
wire n_0_0_145;
wire n_0_0_146;
wire n_0_0_147;
wire n_0_418;
wire n_0_0_148;
wire n_0_0_149;
wire n_0_0_150;
wire n_0_0_151;
wire n_0_0_152;
wire n_0_0_153;
wire n_0_0_154;
wire n_0_0_155;
wire n_0_0_156;
wire n_0_226;
wire n_0_0_70;
wire n_0_0_71;
wire n_0_361;
wire n_0_0_82;
wire n_0_0_72;
wire n_0_0_158;
wire n_0_362;
wire n_0_0_83;
wire n_0_0_159;
wire n_0_0_160;
wire n_0_363;
wire n_0_0_84;
wire n_0_0_161;
wire n_0_0_162;
wire n_0_364;
wire n_0_0_85;
wire n_0_0_163;
wire n_0_0_164;
wire n_0_365;
wire n_0_0_86;
wire n_0_0_165;
wire n_0_0_166;
wire n_0_366;
wire n_0_0_87;
wire n_0_0_167;
wire n_0_0_168;
wire n_0_0_157;
wire n_0_225;
wire n_0_0_169;
wire n_0_0_170;
wire n_0_227;
wire n_0_0_171;
wire n_0_0_73;
wire n_0_0_172;
wire n_0_0_74;
wire n_0_356;
wire n_0_0_77;
wire n_0_0_173;
wire n_0_0_106;
wire n_0_0_174;
wire n_0_0_108;
wire n_0_0_144;
wire \counter[6] ;
wire \counter[5] ;
wire \counter[4] ;
wire \counter[3] ;
wire \counter[2] ;
wire \counter[1] ;
wire \counter[0] ;
wire \A_r[31] ;
wire \A_r[30] ;
wire \A_r[29] ;
wire \A_r[28] ;
wire \A_r[27] ;
wire \A_r[26] ;
wire \A_r[25] ;
wire \A_r[24] ;
wire \A_r[23] ;
wire \A_r[22] ;
wire \A_r[21] ;
wire \A_r[20] ;
wire \A_r[19] ;
wire \A_r[18] ;
wire \A_r[17] ;
wire \A_r[16] ;
wire \A_r[15] ;
wire \A_r[14] ;
wire \A_r[13] ;
wire \A_r[12] ;
wire \A_r[11] ;
wire \A_r[10] ;
wire \A_r[9] ;
wire \A_r[8] ;
wire \A_r[7] ;
wire \A_r[6] ;
wire \A_r[5] ;
wire \A_r[4] ;
wire \A_r[3] ;
wire \A_r[2] ;
wire \A_r[1] ;
wire \A_r[0] ;
wire \B_r[31] ;
wire \B_r[30] ;
wire \B_r[29] ;
wire \B_r[28] ;
wire \B_r[27] ;
wire \B_r[26] ;
wire \B_r[25] ;
wire \B_r[24] ;
wire \B_r[23] ;
wire \B_r[22] ;
wire \B_r[21] ;
wire \B_r[20] ;
wire \B_r[19] ;
wire \B_r[18] ;
wire \B_r[17] ;
wire \B_r[16] ;
wire \B_r[15] ;
wire \B_r[14] ;
wire \B_r[13] ;
wire \B_r[12] ;
wire \B_r[11] ;
wire \B_r[10] ;
wire \B_r[9] ;
wire \B_r[8] ;
wire \B_r[7] ;
wire \B_r[6] ;
wire \B_r[5] ;
wire \B_r[4] ;
wire \B_r[3] ;
wire \B_r[2] ;
wire \B_r[1] ;
wire \B_r[0] ;
wire \Accumulator[30] ;
wire \Accumulator[29] ;
wire \Accumulator[28] ;
wire \Accumulator[27] ;
wire \Accumulator[26] ;
wire \Accumulator[25] ;
wire \Accumulator[24] ;
wire \Accumulator[23] ;
wire \Accumulator[22] ;
wire \Accumulator[21] ;
wire \Accumulator[20] ;
wire \Accumulator[19] ;
wire \Accumulator[18] ;
wire \Accumulator[17] ;
wire \Accumulator[16] ;
wire \Accumulator[15] ;
wire \Accumulator[14] ;
wire \Accumulator[13] ;
wire \Accumulator[12] ;
wire \Accumulator[11] ;
wire \Accumulator[10] ;
wire \Accumulator[9] ;
wire \Accumulator[8] ;
wire \Accumulator[7] ;
wire \Accumulator[6] ;
wire \Accumulator[5] ;
wire \Accumulator[4] ;
wire \Accumulator[3] ;
wire \Accumulator[2] ;
wire \Accumulator[1] ;
wire \Accumulator[0] ;
wire negative;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire hfn_ipo_n23;
wire hfn_ipo_n24;
wire hfn_ipo_n26;
wire hfn_ipo_n27;
wire hfn_ipo_n28;
wire hfn_ipo_n29;
wire hfn_ipo_n30;
wire hfn_ipo_n31;
wire CTS_n_tid0_169;
wire CTS_n_tid1_121;
wire hfn_ipo_n25;
wire CTS_n_tid0_170;
wire drc_ipo_n35;
wire drc_ipo_n36;
wire drc_ipo_n37;
wire drc_ipo_n38;
wire drc_ipo_n39;
wire drc_ipo_n40;
wire drc_ipo_n41;
wire drc_ipo_n42;
wire drc_ipo_n43;
wire drc_ipo_n44;
wire drc_ipo_n45;
wire drc_ipo_n46;
wire drc_ipo_n47;
wire drc_ipo_n48;
wire drc_ipo_n49;
wire drc_ipo_n50;
wire drc_ipo_n51;
wire drc_ipo_n52;
wire drc_ipo_n53;
wire drc_ipo_n54;
wire drc_ipo_n55;
wire drc_ipo_n56;
wire drc_ipo_n57;
wire drc_ipo_n58;
wire drc_ipo_n59;
wire drc_ipo_n60;
wire drc_ipo_n61;
wire drc_ipo_n62;
wire drc_ipo_n63;
wire drc_ipo_n64;
wire drc_ipo_n65;
wire drc_ipo_n66;
wire drc_ipo_n67;
wire drc_ipo_n68;
wire drc_ipo_n69;
wire drc_ipo_n70;
wire drc_ipo_n71;
wire drc_ipo_n72;
wire drc_ipo_n73;
wire drc_ipo_n74;
wire drc_ipo_n75;
wire drc_ipo_n76;
wire drc_ipo_n77;
wire drc_ipo_n78;
wire drc_ipo_n79;
wire drc_ipo_n80;
wire drc_ipo_n81;
wire drc_ipo_n82;
wire drc_ipo_n83;
wire drc_ipo_n84;
wire drc_ipo_n85;
wire drc_ipo_n86;
wire drc_ipo_n87;
wire drc_ipo_n88;
wire drc_ipo_n89;
wire drc_ipo_n90;
wire drc_ipo_n91;
wire drc_ipo_n92;
wire drc_ipo_n93;
wire drc_ipo_n94;
wire drc_ipo_n95;
wire drc_ipo_n96;
wire drc_ipo_n97;
wire drc_ipo_n98;
wire drc_ipo_n99;
wire CLOCK_slh__n241;
wire CLOCK_slh__n242;
wire CLOCK_slh__n245;
wire CLOCK_slh__n246;
wire CLOCK_slh__n249;
wire CLOCK_slh__n250;
wire CLOCK_slh__n253;
wire CLOCK_slh__n254;
wire CLOCK_slh__n257;
wire CLOCK_slh__n258;
wire CLOCK_slh__n261;
wire CLOCK_slh__n263;
wire CLOCK_slh__n265;
wire CLOCK_slh__n267;
wire CLOCK_slh__n269;
wire CLOCK_slh__n271;
wire CLOCK_slh__n273;
wire CLOCK_slh__n275;
wire CLOCK_slh__n277;
wire CLOCK_slh__n279;
wire CLOCK_slh__n281;
wire CLOCK_slh__n283;
wire CLOCK_slh__n285;
wire CLOCK_slh__n287;
wire CLOCK_slh__n289;
wire CLOCK_slh__n291;
wire CLOCK_slh__n293;
wire CLOCK_slh__n295;
wire CLOCK_slh__n297;
wire CLOCK_slh__n299;
wire CLOCK_slh__n300;


DFF_X1 negative_reg (.Q (negative), .CK (CTS_n_tid0_168), .D (n_0_165));
DFF_X1 \Accumulator_reg[0]  (.Q (\Accumulator[0] ), .CK (CTS_n_tid0_168), .D (n_0_229));
DFF_X1 \Accumulator_reg[1]  (.Q (\Accumulator[1] ), .CK (CTS_n_tid0_169), .D (n_0_230));
DFF_X1 \Accumulator_reg[2]  (.Q (\Accumulator[2] ), .CK (CTS_n_tid0_169), .D (n_0_231));
DFF_X1 \Accumulator_reg[3]  (.Q (\Accumulator[3] ), .CK (CTS_n_tid0_169), .D (n_0_232));
DFF_X1 \Accumulator_reg[4]  (.Q (\Accumulator[4] ), .CK (CTS_n_tid0_169), .D (n_0_233));
DFF_X1 \Accumulator_reg[5]  (.Q (\Accumulator[5] ), .CK (CTS_n_tid0_169), .D (n_0_234));
DFF_X1 \Accumulator_reg[6]  (.Q (\Accumulator[6] ), .CK (CTS_n_tid0_169), .D (n_0_235));
DFF_X1 \Accumulator_reg[7]  (.Q (\Accumulator[7] ), .CK (CTS_n_tid0_169), .D (n_0_236));
DFF_X1 \Accumulator_reg[8]  (.Q (\Accumulator[8] ), .CK (CTS_n_tid0_169), .D (n_0_237));
DFF_X1 \Accumulator_reg[9]  (.Q (\Accumulator[9] ), .CK (CTS_n_tid0_169), .D (n_0_238));
DFF_X1 \Accumulator_reg[10]  (.Q (\Accumulator[10] ), .CK (CTS_n_tid0_169), .D (n_0_239));
DFF_X1 \Accumulator_reg[11]  (.Q (\Accumulator[11] ), .CK (CTS_n_tid0_169), .D (n_0_240));
DFF_X1 \Accumulator_reg[12]  (.Q (\Accumulator[12] ), .CK (CTS_n_tid0_169), .D (n_0_241));
DFF_X1 \Accumulator_reg[13]  (.Q (\Accumulator[13] ), .CK (CTS_n_tid0_169), .D (n_0_242));
DFF_X1 \Accumulator_reg[14]  (.Q (\Accumulator[14] ), .CK (CTS_n_tid0_169), .D (n_0_243));
DFF_X1 \Accumulator_reg[15]  (.Q (\Accumulator[15] ), .CK (CTS_n_tid0_169), .D (n_0_244));
DFF_X1 \Accumulator_reg[16]  (.Q (\Accumulator[16] ), .CK (CTS_n_tid0_169), .D (n_0_245));
DFF_X1 \Accumulator_reg[17]  (.Q (\Accumulator[17] ), .CK (CTS_n_tid0_169), .D (n_0_246));
DFF_X1 \Accumulator_reg[18]  (.Q (\Accumulator[18] ), .CK (CTS_n_tid0_169), .D (n_0_247));
DFF_X1 \Accumulator_reg[19]  (.Q (\Accumulator[19] ), .CK (CTS_n_tid0_169), .D (n_0_248));
DFF_X1 \Accumulator_reg[20]  (.Q (\Accumulator[20] ), .CK (CTS_n_tid0_169), .D (n_0_249));
DFF_X1 \Accumulator_reg[21]  (.Q (\Accumulator[21] ), .CK (CTS_n_tid0_169), .D (n_0_250));
DFF_X1 \Accumulator_reg[22]  (.Q (\Accumulator[22] ), .CK (CTS_n_tid0_169), .D (n_0_251));
DFF_X1 \Accumulator_reg[23]  (.Q (\Accumulator[23] ), .CK (CTS_n_tid0_169), .D (n_0_252));
DFF_X1 \Accumulator_reg[24]  (.Q (\Accumulator[24] ), .CK (CTS_n_tid0_168), .D (n_0_253));
DFF_X1 \Accumulator_reg[25]  (.Q (\Accumulator[25] ), .CK (CTS_n_tid0_168), .D (n_0_254));
DFF_X1 \Accumulator_reg[26]  (.Q (\Accumulator[26] ), .CK (CTS_n_tid0_168), .D (n_0_255));
DFF_X1 \Accumulator_reg[27]  (.Q (\Accumulator[27] ), .CK (CTS_n_tid0_168), .D (n_0_256));
DFF_X1 \Accumulator_reg[28]  (.Q (\Accumulator[28] ), .CK (CTS_n_tid0_168), .D (n_0_257));
DFF_X1 \Accumulator_reg[29]  (.Q (\Accumulator[29] ), .CK (CTS_n_tid0_168), .D (n_0_258));
DFF_X1 \Accumulator_reg[30]  (.Q (\Accumulator[30] ), .CK (CTS_n_tid0_168), .D (n_0_259));
DFF_X1 \B_r_reg[0]  (.Q (\B_r[0] ), .CK (CTS_n_tid0_168), .D (n_0_260));
DFF_X1 \B_r_reg[1]  (.Q (\B_r[1] ), .CK (CTS_n_tid0_168), .D (n_0_261));
DFF_X1 \B_r_reg[2]  (.Q (\B_r[2] ), .CK (CTS_n_tid0_168), .D (n_0_262));
DFF_X1 \B_r_reg[3]  (.Q (\B_r[3] ), .CK (CTS_n_tid0_168), .D (n_0_263));
DFF_X1 \B_r_reg[4]  (.Q (\B_r[4] ), .CK (CTS_n_tid0_168), .D (n_0_264));
DFF_X1 \B_r_reg[5]  (.Q (\B_r[5] ), .CK (CTS_n_tid0_168), .D (n_0_265));
DFF_X1 \B_r_reg[6]  (.Q (\B_r[6] ), .CK (CTS_n_tid0_168), .D (n_0_266));
DFF_X1 \B_r_reg[7]  (.Q (\B_r[7] ), .CK (CTS_n_tid0_168), .D (n_0_267));
DFF_X1 \B_r_reg[8]  (.Q (\B_r[8] ), .CK (CTS_n_tid0_168), .D (n_0_268));
DFF_X1 \B_r_reg[9]  (.Q (\B_r[9] ), .CK (CTS_n_tid0_168), .D (n_0_269));
DFF_X1 \B_r_reg[10]  (.Q (\B_r[10] ), .CK (CTS_n_tid0_168), .D (n_0_270));
DFF_X1 \B_r_reg[11]  (.Q (\B_r[11] ), .CK (CTS_n_tid0_168), .D (n_0_271));
DFF_X1 \B_r_reg[12]  (.Q (\B_r[12] ), .CK (CTS_n_tid0_168), .D (n_0_272));
DFF_X1 \B_r_reg[13]  (.Q (\B_r[13] ), .CK (CTS_n_tid0_168), .D (n_0_273));
DFF_X1 \B_r_reg[14]  (.Q (\B_r[14] ), .CK (CTS_n_tid0_168), .D (n_0_274));
DFF_X1 \B_r_reg[15]  (.Q (\B_r[15] ), .CK (CTS_n_tid0_168), .D (n_0_275));
DFF_X1 \B_r_reg[16]  (.Q (\B_r[16] ), .CK (CTS_n_tid0_168), .D (n_0_276));
DFF_X1 \B_r_reg[17]  (.Q (\B_r[17] ), .CK (CTS_n_tid0_168), .D (n_0_277));
DFF_X1 \B_r_reg[18]  (.Q (\B_r[18] ), .CK (CTS_n_tid0_168), .D (n_0_278));
DFF_X1 \B_r_reg[19]  (.Q (\B_r[19] ), .CK (CTS_n_tid0_168), .D (n_0_279));
DFF_X1 \B_r_reg[20]  (.Q (\B_r[20] ), .CK (CTS_n_tid0_168), .D (n_0_280));
DFF_X1 \B_r_reg[21]  (.Q (\B_r[21] ), .CK (CTS_n_tid0_168), .D (n_0_281));
DFF_X1 \B_r_reg[22]  (.Q (\B_r[22] ), .CK (CTS_n_tid0_168), .D (n_0_282));
DFF_X1 \B_r_reg[23]  (.Q (\B_r[23] ), .CK (CTS_n_tid0_168), .D (n_0_283));
DFF_X1 \B_r_reg[24]  (.Q (\B_r[24] ), .CK (CTS_n_tid0_168), .D (n_0_284));
DFF_X1 \B_r_reg[25]  (.Q (\B_r[25] ), .CK (CTS_n_tid0_168), .D (n_0_285));
DFF_X1 \B_r_reg[26]  (.Q (\B_r[26] ), .CK (CTS_n_tid0_168), .D (n_0_286));
DFF_X1 \B_r_reg[27]  (.Q (\B_r[27] ), .CK (CTS_n_tid0_168), .D (n_0_287));
DFF_X1 \B_r_reg[28]  (.Q (\B_r[28] ), .CK (CTS_n_tid0_168), .D (n_0_288));
DFF_X1 \B_r_reg[29]  (.Q (\B_r[29] ), .CK (CTS_n_tid0_168), .D (n_0_289));
DFF_X1 \B_r_reg[30]  (.Q (\B_r[30] ), .CK (CTS_n_tid0_168), .D (n_0_290));
DFF_X1 \B_r_reg[31]  (.Q (\B_r[31] ), .CK (CTS_n_tid0_169), .D (n_0_291));
DFF_X1 \A_r_reg[0]  (.Q (\A_r[0] ), .CK (CTS_n_tid0_168), .D (n_0_386));
DFF_X1 \A_r_reg[1]  (.Q (\A_r[1] ), .CK (CTS_n_tid0_169), .D (n_0_387));
DFF_X1 \A_r_reg[2]  (.Q (\A_r[2] ), .CK (CTS_n_tid0_169), .D (n_0_388));
DFF_X1 \A_r_reg[3]  (.Q (\A_r[3] ), .CK (CTS_n_tid0_169), .D (n_0_389));
DFF_X1 \A_r_reg[4]  (.Q (\A_r[4] ), .CK (CTS_n_tid0_169), .D (n_0_390));
DFF_X1 \A_r_reg[5]  (.Q (\A_r[5] ), .CK (CTS_n_tid0_169), .D (n_0_391));
DFF_X1 \A_r_reg[6]  (.Q (\A_r[6] ), .CK (CTS_n_tid0_169), .D (n_0_392));
DFF_X1 \A_r_reg[7]  (.Q (\A_r[7] ), .CK (CTS_n_tid0_169), .D (n_0_393));
DFF_X1 \A_r_reg[8]  (.Q (\A_r[8] ), .CK (CTS_n_tid0_169), .D (n_0_394));
DFF_X1 \A_r_reg[9]  (.Q (\A_r[9] ), .CK (CTS_n_tid0_169), .D (n_0_395));
DFF_X1 \A_r_reg[10]  (.Q (\A_r[10] ), .CK (CTS_n_tid0_169), .D (n_0_396));
DFF_X1 \A_r_reg[11]  (.Q (\A_r[11] ), .CK (CTS_n_tid0_169), .D (n_0_397));
DFF_X1 \A_r_reg[12]  (.Q (\A_r[12] ), .CK (CTS_n_tid0_169), .D (n_0_398));
DFF_X1 \A_r_reg[13]  (.Q (\A_r[13] ), .CK (CTS_n_tid0_169), .D (n_0_399));
DFF_X1 \A_r_reg[14]  (.Q (\A_r[14] ), .CK (CTS_n_tid0_169), .D (n_0_400));
DFF_X1 \A_r_reg[15]  (.Q (\A_r[15] ), .CK (CTS_n_tid0_169), .D (n_0_401));
DFF_X1 \A_r_reg[16]  (.Q (\A_r[16] ), .CK (CTS_n_tid0_169), .D (n_0_402));
DFF_X1 \A_r_reg[17]  (.Q (\A_r[17] ), .CK (CTS_n_tid0_169), .D (n_0_403));
DFF_X1 \A_r_reg[18]  (.Q (\A_r[18] ), .CK (CTS_n_tid0_169), .D (n_0_404));
DFF_X1 \A_r_reg[19]  (.Q (\A_r[19] ), .CK (CTS_n_tid0_169), .D (n_0_405));
DFF_X1 \A_r_reg[20]  (.Q (\A_r[20] ), .CK (CTS_n_tid0_169), .D (n_0_406));
DFF_X1 \A_r_reg[21]  (.Q (\A_r[21] ), .CK (CTS_n_tid0_169), .D (n_0_407));
DFF_X1 \A_r_reg[22]  (.Q (\A_r[22] ), .CK (CTS_n_tid0_169), .D (n_0_408));
DFF_X1 \A_r_reg[23]  (.Q (\A_r[23] ), .CK (CTS_n_tid0_169), .D (n_0_409));
DFF_X1 \A_r_reg[24]  (.Q (\A_r[24] ), .CK (CTS_n_tid0_169), .D (n_0_410));
DFF_X1 \A_r_reg[25]  (.Q (\A_r[25] ), .CK (CTS_n_tid0_169), .D (n_0_411));
DFF_X1 \A_r_reg[26]  (.Q (\A_r[26] ), .CK (CTS_n_tid0_168), .D (n_0_412));
DFF_X1 \A_r_reg[27]  (.Q (\A_r[27] ), .CK (CTS_n_tid0_169), .D (n_0_413));
DFF_X1 \A_r_reg[28]  (.Q (\A_r[28] ), .CK (CTS_n_tid0_168), .D (n_0_414));
DFF_X1 \A_r_reg[29]  (.Q (\A_r[29] ), .CK (CTS_n_tid0_168), .D (n_0_415));
DFF_X1 \A_r_reg[30]  (.Q (\A_r[30] ), .CK (CTS_n_tid0_168), .D (n_0_416));
DFF_X1 \A_r_reg[31]  (.Q (\A_r[31] ), .CK (CTS_n_tid0_168), .D (n_0_417));
DFF_X1 \counter_reg[0]  (.Q (\counter[0] ), .CK (CTS_n_tid0_168), .D (n_0_158));
DFF_X1 \counter_reg[1]  (.Q (\counter[1] ), .CK (CTS_n_tid0_168), .D (n_0_159));
DFF_X1 \counter_reg[2]  (.Q (\counter[2] ), .CK (CTS_n_tid0_168), .D (n_0_160));
DFF_X1 \counter_reg[3]  (.Q (\counter[3] ), .CK (CTS_n_tid0_169), .D (n_0_161));
DFF_X1 \counter_reg[4]  (.Q (\counter[4] ), .CK (CTS_n_tid0_168), .D (n_0_162));
DFF_X1 \counter_reg[5]  (.Q (\counter[5] ), .CK (CTS_n_tid0_168), .D (n_0_163));
DFF_X1 \counter_reg[6]  (.Q (\counter[6] ), .CK (CTS_n_tid0_169), .D (n_0_164));
NAND2_X2 i_0_0_430 (.ZN (n_0_0_144), .A1 (n_0_0_145), .A2 (n_0_0_146));
NOR2_X4 i_0_0_429 (.ZN (n_0_0_108), .A1 (n_0_0_154), .A2 (hfn_ipo_n30));
NAND2_X1 i_0_0_428 (.ZN (n_0_0_174), .A1 (n_0_33), .A2 (n_0_0_108));
NOR2_X4 i_0_0_427 (.ZN (n_0_0_106), .A1 (drc_ipo_n66), .A2 (hfn_ipo_n30));
AOI22_X1 i_0_0_426 (.ZN (n_0_0_173), .A1 (n_0_0_106), .A2 (drc_ipo_n37), .B1 (\B_r[2] ), .B2 (hfn_ipo_n29));
AND2_X1 i_0_0_425 (.ZN (n_0_0_77), .A1 (n_0_0_174), .A2 (n_0_0_173));
INV_X1 i_0_0_424 (.ZN (n_0_356), .A (n_0_0_77));
NOR3_X1 i_0_0_423 (.ZN (n_0_0_74), .A1 (n_0_0_148), .A2 (hfn_ipo_n23), .A3 (n_0_0_153));
NAND2_X1 i_0_0_422 (.ZN (n_0_0_172), .A1 (n_0_156), .A2 (hfn_ipo_n28));
AOI21_X1 i_0_0_421 (.ZN (n_0_0_73), .A (hfn_ipo_n23), .B1 (n_0_0_149), .B2 (negative));
NAND2_X1 i_0_0_420 (.ZN (n_0_0_171), .A1 (n_0_94), .A2 (hfn_ipo_n26));
NAND2_X1 i_0_0_419 (.ZN (n_0_227), .A1 (n_0_0_172), .A2 (n_0_0_171));
NAND2_X1 i_0_0_418 (.ZN (n_0_0_170), .A1 (n_0_154), .A2 (hfn_ipo_n28));
NAND2_X1 i_0_0_417 (.ZN (n_0_0_169), .A1 (n_0_92), .A2 (hfn_ipo_n26));
NAND2_X1 i_0_0_416 (.ZN (n_0_225), .A1 (n_0_0_170), .A2 (n_0_0_169));
INV_X2 i_0_0_415 (.ZN (n_0_0_157), .A (hfn_ipo_n24));
NAND2_X1 i_0_0_414 (.ZN (n_0_0_168), .A1 (n_0_43), .A2 (n_0_0_108));
AOI22_X1 i_0_0_413 (.ZN (n_0_0_167), .A1 (n_0_0_106), .A2 (drc_ipo_n47), .B1 (\B_r[12] ), .B2 (hfn_ipo_n29));
AND2_X1 i_0_0_399 (.ZN (n_0_0_87), .A1 (n_0_0_168), .A2 (n_0_0_167));
INV_X1 i_0_0_331 (.ZN (n_0_366), .A (n_0_0_87));
NAND2_X1 i_0_0_328 (.ZN (n_0_0_166), .A1 (n_0_42), .A2 (n_0_0_108));
AOI22_X1 i_0_0_291 (.ZN (n_0_0_165), .A1 (n_0_0_106), .A2 (drc_ipo_n46), .B1 (\B_r[11] ), .B2 (hfn_ipo_n29));
AND2_X1 i_0_0_290 (.ZN (n_0_0_86), .A1 (n_0_0_166), .A2 (n_0_0_165));
INV_X1 i_0_0_289 (.ZN (n_0_365), .A (n_0_0_86));
NAND2_X1 i_0_0_288 (.ZN (n_0_0_164), .A1 (n_0_41), .A2 (n_0_0_108));
AOI22_X1 i_0_0_287 (.ZN (n_0_0_163), .A1 (n_0_0_106), .A2 (drc_ipo_n45), .B1 (\B_r[10] ), .B2 (hfn_ipo_n29));
AND2_X1 i_0_0_286 (.ZN (n_0_0_85), .A1 (n_0_0_164), .A2 (n_0_0_163));
INV_X1 i_0_0_285 (.ZN (n_0_364), .A (n_0_0_85));
NAND2_X1 i_0_0_284 (.ZN (n_0_0_162), .A1 (n_0_40), .A2 (n_0_0_108));
AOI22_X1 i_0_0_283 (.ZN (n_0_0_161), .A1 (n_0_0_106), .A2 (drc_ipo_n44), .B1 (\B_r[9] ), .B2 (hfn_ipo_n29));
AND2_X1 i_0_0_282 (.ZN (n_0_0_84), .A1 (n_0_0_162), .A2 (n_0_0_161));
INV_X1 i_0_0_281 (.ZN (n_0_363), .A (n_0_0_84));
NAND2_X1 i_0_0_280 (.ZN (n_0_0_160), .A1 (n_0_39), .A2 (n_0_0_108));
AOI22_X1 i_0_0_271 (.ZN (n_0_0_159), .A1 (n_0_0_106), .A2 (drc_ipo_n43), .B1 (\B_r[8] ), .B2 (hfn_ipo_n29));
AND2_X1 i_0_0_270 (.ZN (n_0_0_83), .A1 (n_0_0_160), .A2 (n_0_0_159));
INV_X1 i_0_0_140 (.ZN (n_0_362), .A (n_0_0_83));
NAND2_X1 i_0_0_138 (.ZN (n_0_0_158), .A1 (n_0_38), .A2 (n_0_0_108));
AOI22_X1 i_0_0_137 (.ZN (n_0_0_72), .A1 (n_0_0_106), .A2 (drc_ipo_n42), .B1 (\B_r[7] ), .B2 (hfn_ipo_n29));
AND2_X1 i_0_0_136 (.ZN (n_0_0_82), .A1 (n_0_0_158), .A2 (n_0_0_72));
INV_X1 i_0_0_135 (.ZN (n_0_361), .A (n_0_0_82));
NAND2_X1 i_0_0_134 (.ZN (n_0_0_71), .A1 (n_0_155), .A2 (hfn_ipo_n28));
NAND2_X1 i_0_0_133 (.ZN (n_0_0_70), .A1 (n_0_93), .A2 (hfn_ipo_n26));
NAND2_X1 i_0_0_132 (.ZN (n_0_226), .A1 (n_0_0_71), .A2 (n_0_0_70));
INV_X1 i_0_0_412 (.ZN (n_0_0_156), .A (\counter[6] ));
INV_X1 i_0_0_411 (.ZN (n_0_0_155), .A (drc_ipo_n98));
INV_X1 i_0_0_410 (.ZN (n_0_0_154), .A (drc_ipo_n66));
INV_X1 i_0_0_409 (.ZN (n_0_0_153), .A (negative));
INV_X1 i_0_0_408 (.ZN (n_0_0_152), .A (n_0_0_4));
NAND3_X1 i_0_0_407 (.ZN (n_0_0_151), .A1 (\counter[2] ), .A2 (\counter[1] ), .A3 (\counter[0] ));
NAND2_X1 i_0_0_406 (.ZN (n_0_0_150), .A1 (\counter[4] ), .A2 (\counter[3] ));
NOR4_X1 i_0_0_405 (.ZN (n_0_0_149), .A1 (\counter[6] ), .A2 (\counter[5] ), .A3 (n_0_0_150), .A4 (n_0_0_151));
INV_X1 i_0_0_404 (.ZN (n_0_0_148), .A (n_0_0_149));
NAND2_X1 i_0_0_403 (.ZN (n_0_418), .A1 (n_0_0_157), .A2 (n_0_0_148));
INV_X1 i_0_0_402 (.ZN (n_0_0_147), .A (n_0_418));
NOR3_X1 i_0_0_401 (.ZN (n_0_0_146), .A1 (\counter[2] ), .A2 (\counter[1] ), .A3 (\counter[0] ));
NOR4_X1 i_0_0_400 (.ZN (n_0_0_145), .A1 (\counter[6] ), .A2 (\counter[5] ), .A3 (\counter[4] ), .A4 (\counter[3] ));
INV_X1 i_0_0_398 (.ZN (n_0_0_143), .A (hfn_ipo_n29));
NOR2_X4 i_0_0_397 (.ZN (n_0_0_142), .A1 (n_0_0_155), .A2 (hfn_ipo_n30));
AOI22_X1 i_0_0_396 (.ZN (n_0_0_141), .A1 (\A_r[31] ), .A2 (hfn_ipo_n30), .B1 (n_0_31), .B2 (n_0_0_142));
NOR2_X1 i_0_0_395 (.ZN (n_0_417), .A1 (hfn_ipo_n23), .A2 (n_0_0_141));
NOR2_X4 i_0_0_394 (.ZN (n_0_0_140), .A1 (drc_ipo_n98), .A2 (hfn_ipo_n30));
AOI222_X1 i_0_0_393 (.ZN (n_0_0_139), .A1 (\A_r[30] ), .A2 (hfn_ipo_n30), .B1 (drc_ipo_n97)
    , .B2 (n_0_0_140), .C1 (n_0_30), .C2 (n_0_0_142));
NOR2_X1 i_0_0_392 (.ZN (n_0_416), .A1 (hfn_ipo_n23), .A2 (n_0_0_139));
AOI222_X1 i_0_0_391 (.ZN (n_0_0_138), .A1 (\A_r[29] ), .A2 (hfn_ipo_n30), .B1 (drc_ipo_n96)
    , .B2 (n_0_0_140), .C1 (n_0_29), .C2 (n_0_0_142));
NOR2_X1 i_0_0_390 (.ZN (n_0_415), .A1 (hfn_ipo_n23), .A2 (n_0_0_138));
AOI222_X1 i_0_0_389 (.ZN (n_0_0_137), .A1 (\A_r[28] ), .A2 (hfn_ipo_n30), .B1 (drc_ipo_n95)
    , .B2 (n_0_0_140), .C1 (n_0_28), .C2 (n_0_0_142));
NOR2_X1 i_0_0_388 (.ZN (n_0_414), .A1 (hfn_ipo_n23), .A2 (n_0_0_137));
AOI222_X1 i_0_0_387 (.ZN (n_0_0_136), .A1 (\A_r[27] ), .A2 (hfn_ipo_n30), .B1 (drc_ipo_n94)
    , .B2 (n_0_0_140), .C1 (n_0_27), .C2 (n_0_0_142));
NOR2_X1 i_0_0_386 (.ZN (n_0_413), .A1 (hfn_ipo_n23), .A2 (n_0_0_136));
AOI222_X1 i_0_0_385 (.ZN (n_0_0_135), .A1 (\A_r[26] ), .A2 (hfn_ipo_n30), .B1 (drc_ipo_n93)
    , .B2 (n_0_0_140), .C1 (n_0_26), .C2 (n_0_0_142));
NOR2_X1 i_0_0_384 (.ZN (n_0_412), .A1 (hfn_ipo_n23), .A2 (n_0_0_135));
AOI222_X1 i_0_0_383 (.ZN (n_0_0_134), .A1 (\A_r[25] ), .A2 (n_0_0_144), .B1 (drc_ipo_n92)
    , .B2 (n_0_0_140), .C1 (n_0_25), .C2 (n_0_0_142));
NOR2_X1 i_0_0_382 (.ZN (n_0_411), .A1 (hfn_ipo_n23), .A2 (n_0_0_134));
AOI222_X1 i_0_0_381 (.ZN (n_0_0_133), .A1 (\A_r[24] ), .A2 (n_0_0_144), .B1 (drc_ipo_n91)
    , .B2 (n_0_0_140), .C1 (n_0_24), .C2 (n_0_0_142));
NOR2_X1 i_0_0_380 (.ZN (n_0_410), .A1 (hfn_ipo_n24), .A2 (n_0_0_133));
AOI222_X1 i_0_0_379 (.ZN (n_0_0_132), .A1 (\A_r[23] ), .A2 (n_0_0_144), .B1 (drc_ipo_n90)
    , .B2 (n_0_0_140), .C1 (n_0_23), .C2 (n_0_0_142));
NOR2_X1 i_0_0_378 (.ZN (n_0_409), .A1 (hfn_ipo_n24), .A2 (n_0_0_132));
AOI222_X1 i_0_0_377 (.ZN (n_0_0_131), .A1 (\A_r[22] ), .A2 (n_0_0_144), .B1 (drc_ipo_n89)
    , .B2 (n_0_0_140), .C1 (n_0_22), .C2 (n_0_0_142));
NOR2_X1 i_0_0_376 (.ZN (n_0_408), .A1 (hfn_ipo_n24), .A2 (n_0_0_131));
AOI222_X1 i_0_0_375 (.ZN (n_0_0_130), .A1 (\A_r[21] ), .A2 (n_0_0_144), .B1 (drc_ipo_n88)
    , .B2 (n_0_0_140), .C1 (n_0_21), .C2 (n_0_0_142));
NOR2_X1 i_0_0_374 (.ZN (n_0_407), .A1 (hfn_ipo_n24), .A2 (n_0_0_130));
AOI222_X1 i_0_0_373 (.ZN (n_0_0_129), .A1 (\A_r[20] ), .A2 (n_0_0_144), .B1 (drc_ipo_n87)
    , .B2 (n_0_0_140), .C1 (n_0_20), .C2 (n_0_0_142));
NOR2_X1 i_0_0_372 (.ZN (n_0_406), .A1 (hfn_ipo_n24), .A2 (n_0_0_129));
AOI222_X1 i_0_0_371 (.ZN (n_0_0_128), .A1 (\A_r[19] ), .A2 (n_0_0_144), .B1 (drc_ipo_n86)
    , .B2 (n_0_0_140), .C1 (n_0_19), .C2 (n_0_0_142));
NOR2_X1 i_0_0_370 (.ZN (n_0_405), .A1 (hfn_ipo_n24), .A2 (n_0_0_128));
AOI222_X1 i_0_0_369 (.ZN (n_0_0_127), .A1 (\A_r[18] ), .A2 (n_0_0_144), .B1 (drc_ipo_n85)
    , .B2 (n_0_0_140), .C1 (n_0_18), .C2 (n_0_0_142));
NOR2_X1 i_0_0_368 (.ZN (n_0_404), .A1 (hfn_ipo_n24), .A2 (n_0_0_127));
AOI222_X1 i_0_0_367 (.ZN (n_0_0_126), .A1 (\A_r[17] ), .A2 (n_0_0_144), .B1 (drc_ipo_n84)
    , .B2 (n_0_0_140), .C1 (n_0_17), .C2 (n_0_0_142));
NOR2_X1 i_0_0_366 (.ZN (n_0_403), .A1 (hfn_ipo_n24), .A2 (n_0_0_126));
AOI222_X1 i_0_0_365 (.ZN (n_0_0_125), .A1 (\A_r[16] ), .A2 (n_0_0_144), .B1 (drc_ipo_n83)
    , .B2 (n_0_0_140), .C1 (n_0_16), .C2 (n_0_0_142));
NOR2_X1 i_0_0_364 (.ZN (n_0_402), .A1 (hfn_ipo_n24), .A2 (n_0_0_125));
AOI222_X1 i_0_0_363 (.ZN (n_0_0_124), .A1 (\A_r[15] ), .A2 (n_0_0_144), .B1 (drc_ipo_n82)
    , .B2 (n_0_0_140), .C1 (n_0_15), .C2 (n_0_0_142));
NOR2_X1 i_0_0_362 (.ZN (n_0_401), .A1 (hfn_ipo_n24), .A2 (n_0_0_124));
AOI222_X1 i_0_0_361 (.ZN (n_0_0_123), .A1 (\A_r[14] ), .A2 (n_0_0_144), .B1 (drc_ipo_n81)
    , .B2 (n_0_0_140), .C1 (n_0_14), .C2 (n_0_0_142));
NOR2_X1 i_0_0_360 (.ZN (n_0_400), .A1 (hfn_ipo_n24), .A2 (n_0_0_123));
AOI222_X1 i_0_0_359 (.ZN (n_0_0_122), .A1 (\A_r[13] ), .A2 (n_0_0_144), .B1 (drc_ipo_n80)
    , .B2 (n_0_0_140), .C1 (n_0_13), .C2 (n_0_0_142));
NOR2_X1 i_0_0_358 (.ZN (n_0_399), .A1 (hfn_ipo_n24), .A2 (n_0_0_122));
AOI222_X1 i_0_0_357 (.ZN (n_0_0_121), .A1 (\A_r[12] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n79)
    , .B2 (n_0_0_140), .C1 (n_0_12), .C2 (n_0_0_142));
NOR2_X1 i_0_0_356 (.ZN (n_0_398), .A1 (hfn_ipo_n24), .A2 (n_0_0_121));
AOI222_X1 i_0_0_355 (.ZN (n_0_0_120), .A1 (\A_r[11] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n78)
    , .B2 (n_0_0_140), .C1 (n_0_11), .C2 (n_0_0_142));
NOR2_X1 i_0_0_354 (.ZN (n_0_397), .A1 (hfn_ipo_n24), .A2 (n_0_0_120));
AOI222_X1 i_0_0_353 (.ZN (n_0_0_119), .A1 (\A_r[10] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n77)
    , .B2 (n_0_0_140), .C1 (n_0_10), .C2 (n_0_0_142));
NOR2_X1 i_0_0_352 (.ZN (n_0_396), .A1 (hfn_ipo_n24), .A2 (n_0_0_119));
AOI222_X1 i_0_0_351 (.ZN (n_0_0_118), .A1 (\A_r[9] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n76)
    , .B2 (n_0_0_140), .C1 (n_0_9), .C2 (n_0_0_142));
NOR2_X1 i_0_0_350 (.ZN (n_0_395), .A1 (hfn_ipo_n24), .A2 (n_0_0_118));
AOI222_X1 i_0_0_349 (.ZN (n_0_0_117), .A1 (\A_r[8] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n75)
    , .B2 (n_0_0_140), .C1 (n_0_8), .C2 (n_0_0_142));
NOR2_X1 i_0_0_348 (.ZN (n_0_394), .A1 (hfn_ipo_n24), .A2 (n_0_0_117));
AOI222_X1 i_0_0_347 (.ZN (n_0_0_116), .A1 (\A_r[7] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n74)
    , .B2 (n_0_0_140), .C1 (n_0_7), .C2 (n_0_0_142));
NOR2_X1 i_0_0_346 (.ZN (n_0_393), .A1 (hfn_ipo_n24), .A2 (n_0_0_116));
AOI222_X1 i_0_0_345 (.ZN (n_0_0_115), .A1 (\A_r[6] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n73)
    , .B2 (n_0_0_140), .C1 (n_0_6), .C2 (n_0_0_142));
NOR2_X1 i_0_0_344 (.ZN (n_0_392), .A1 (hfn_ipo_n24), .A2 (n_0_0_115));
AOI222_X1 i_0_0_343 (.ZN (n_0_0_114), .A1 (\A_r[5] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n72)
    , .B2 (n_0_0_140), .C1 (n_0_5), .C2 (n_0_0_142));
NOR2_X1 i_0_0_342 (.ZN (n_0_391), .A1 (hfn_ipo_n24), .A2 (n_0_0_114));
AOI222_X1 i_0_0_341 (.ZN (n_0_0_113), .A1 (\A_r[4] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n71)
    , .B2 (n_0_0_140), .C1 (n_0_4), .C2 (n_0_0_142));
NOR2_X1 i_0_0_340 (.ZN (n_0_390), .A1 (hfn_ipo_n24), .A2 (n_0_0_113));
AOI222_X1 i_0_0_339 (.ZN (n_0_0_112), .A1 (\A_r[3] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n70)
    , .B2 (n_0_0_140), .C1 (n_0_3), .C2 (n_0_0_142));
NOR2_X1 i_0_0_338 (.ZN (n_0_389), .A1 (hfn_ipo_n24), .A2 (n_0_0_112));
AOI222_X1 i_0_0_337 (.ZN (n_0_0_111), .A1 (\A_r[2] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n69)
    , .B2 (n_0_0_140), .C1 (n_0_2), .C2 (n_0_0_142));
NOR2_X1 i_0_0_336 (.ZN (n_0_388), .A1 (hfn_ipo_n24), .A2 (n_0_0_111));
AOI222_X1 i_0_0_335 (.ZN (n_0_0_110), .A1 (\A_r[1] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n68)
    , .B2 (n_0_0_140), .C1 (n_0_1), .C2 (n_0_0_142));
NOR2_X1 i_0_0_334 (.ZN (n_0_387), .A1 (hfn_ipo_n24), .A2 (n_0_0_110));
AOI22_X1 i_0_0_333 (.ZN (n_0_0_109), .A1 (\A_r[0] ), .A2 (hfn_ipo_n31), .B1 (drc_ipo_n67), .B2 (n_0_0_143));
NOR2_X1 i_0_0_332 (.ZN (CLOCK_slh__n273), .A1 (hfn_ipo_n23), .A2 (n_0_0_109));
AOI22_X1 i_0_0_330 (.ZN (n_0_0_107), .A1 (\B_r[31] ), .A2 (hfn_ipo_n29), .B1 (n_0_62), .B2 (n_0_0_108));
INV_X1 i_0_0_329 (.ZN (n_0_385), .A (n_0_0_107));
AOI222_X1 i_0_0_327 (.ZN (n_0_0_105), .A1 (\B_r[30] ), .A2 (hfn_ipo_n29), .B1 (n_0_61)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n65), .C2 (n_0_0_106));
INV_X1 i_0_0_326 (.ZN (n_0_384), .A (n_0_0_105));
AOI222_X1 i_0_0_325 (.ZN (n_0_0_104), .A1 (\B_r[29] ), .A2 (hfn_ipo_n29), .B1 (n_0_60)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n64), .C2 (n_0_0_106));
INV_X1 i_0_0_324 (.ZN (n_0_383), .A (n_0_0_104));
AOI222_X1 i_0_0_323 (.ZN (n_0_0_103), .A1 (\B_r[28] ), .A2 (hfn_ipo_n29), .B1 (n_0_59)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n63), .C2 (n_0_0_106));
INV_X1 i_0_0_322 (.ZN (n_0_382), .A (n_0_0_103));
AOI222_X1 i_0_0_321 (.ZN (n_0_0_102), .A1 (\B_r[27] ), .A2 (hfn_ipo_n29), .B1 (n_0_58)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n62), .C2 (n_0_0_106));
INV_X1 i_0_0_320 (.ZN (n_0_381), .A (n_0_0_102));
AOI222_X1 i_0_0_319 (.ZN (n_0_0_101), .A1 (\B_r[26] ), .A2 (hfn_ipo_n29), .B1 (n_0_57)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n61), .C2 (n_0_0_106));
INV_X1 i_0_0_318 (.ZN (n_0_380), .A (n_0_0_101));
AOI222_X1 i_0_0_317 (.ZN (n_0_0_100), .A1 (\B_r[25] ), .A2 (hfn_ipo_n29), .B1 (n_0_56)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n60), .C2 (n_0_0_106));
INV_X1 i_0_0_316 (.ZN (n_0_379), .A (n_0_0_100));
AOI222_X1 i_0_0_315 (.ZN (n_0_0_99), .A1 (\B_r[24] ), .A2 (hfn_ipo_n29), .B1 (n_0_55)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n59), .C2 (n_0_0_106));
INV_X1 i_0_0_314 (.ZN (n_0_378), .A (n_0_0_99));
AOI222_X1 i_0_0_313 (.ZN (n_0_0_98), .A1 (\B_r[23] ), .A2 (hfn_ipo_n29), .B1 (n_0_54)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n58), .C2 (n_0_0_106));
INV_X1 i_0_0_312 (.ZN (n_0_377), .A (n_0_0_98));
AOI222_X1 i_0_0_311 (.ZN (n_0_0_97), .A1 (\B_r[22] ), .A2 (hfn_ipo_n29), .B1 (n_0_53)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n57), .C2 (n_0_0_106));
INV_X1 i_0_0_310 (.ZN (n_0_376), .A (n_0_0_97));
AOI222_X1 i_0_0_309 (.ZN (n_0_0_96), .A1 (\B_r[21] ), .A2 (hfn_ipo_n29), .B1 (n_0_52)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n56), .C2 (n_0_0_106));
INV_X1 i_0_0_308 (.ZN (n_0_375), .A (n_0_0_96));
AOI222_X1 i_0_0_307 (.ZN (n_0_0_95), .A1 (\B_r[20] ), .A2 (hfn_ipo_n29), .B1 (n_0_51)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n55), .C2 (n_0_0_106));
INV_X1 i_0_0_306 (.ZN (n_0_374), .A (n_0_0_95));
AOI222_X1 i_0_0_305 (.ZN (n_0_0_94), .A1 (\B_r[19] ), .A2 (hfn_ipo_n30), .B1 (n_0_50)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n54), .C2 (n_0_0_106));
INV_X1 i_0_0_304 (.ZN (n_0_373), .A (n_0_0_94));
AOI222_X1 i_0_0_303 (.ZN (n_0_0_93), .A1 (\B_r[18] ), .A2 (hfn_ipo_n30), .B1 (n_0_49)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n53), .C2 (n_0_0_106));
INV_X1 i_0_0_302 (.ZN (n_0_372), .A (n_0_0_93));
AOI222_X1 i_0_0_301 (.ZN (n_0_0_92), .A1 (\B_r[17] ), .A2 (hfn_ipo_n30), .B1 (n_0_48)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n52), .C2 (n_0_0_106));
INV_X1 i_0_0_300 (.ZN (n_0_371), .A (n_0_0_92));
AOI222_X1 i_0_0_299 (.ZN (n_0_0_91), .A1 (\B_r[16] ), .A2 (hfn_ipo_n30), .B1 (n_0_47)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n51), .C2 (n_0_0_106));
INV_X1 i_0_0_298 (.ZN (n_0_370), .A (n_0_0_91));
AOI222_X1 i_0_0_297 (.ZN (n_0_0_90), .A1 (\B_r[15] ), .A2 (hfn_ipo_n30), .B1 (n_0_46)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n50), .C2 (n_0_0_106));
INV_X1 i_0_0_296 (.ZN (n_0_369), .A (n_0_0_90));
AOI222_X1 i_0_0_295 (.ZN (n_0_0_89), .A1 (\B_r[14] ), .A2 (hfn_ipo_n30), .B1 (n_0_45)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n49), .C2 (n_0_0_106));
INV_X1 i_0_0_294 (.ZN (n_0_368), .A (n_0_0_89));
AOI222_X1 i_0_0_293 (.ZN (n_0_0_88), .A1 (\B_r[13] ), .A2 (hfn_ipo_n30), .B1 (n_0_44)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n48), .C2 (n_0_0_106));
INV_X1 i_0_0_292 (.ZN (n_0_367), .A (n_0_0_88));
AOI222_X1 i_0_0_279 (.ZN (n_0_0_81), .A1 (\B_r[6] ), .A2 (hfn_ipo_n29), .B1 (n_0_37)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n41), .C2 (n_0_0_106));
INV_X1 i_0_0_278 (.ZN (n_0_360), .A (n_0_0_81));
AOI222_X1 i_0_0_277 (.ZN (n_0_0_80), .A1 (\B_r[5] ), .A2 (hfn_ipo_n29), .B1 (n_0_36)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n40), .C2 (n_0_0_106));
INV_X1 i_0_0_276 (.ZN (n_0_359), .A (n_0_0_80));
AOI222_X1 i_0_0_275 (.ZN (n_0_0_79), .A1 (\B_r[4] ), .A2 (hfn_ipo_n29), .B1 (n_0_35)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n39), .C2 (n_0_0_106));
INV_X1 i_0_0_274 (.ZN (n_0_358), .A (n_0_0_79));
AOI222_X1 i_0_0_273 (.ZN (n_0_0_78), .A1 (\B_r[3] ), .A2 (hfn_ipo_n29), .B1 (n_0_34)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n38), .C2 (n_0_0_106));
INV_X1 i_0_0_272 (.ZN (n_0_357), .A (n_0_0_78));
AOI222_X1 i_0_0_269 (.ZN (n_0_0_76), .A1 (\B_r[1] ), .A2 (hfn_ipo_n29), .B1 (n_0_32)
    , .B2 (n_0_0_108), .C1 (drc_ipo_n36), .C2 (n_0_0_106));
INV_X1 i_0_0_268 (.ZN (n_0_355), .A (n_0_0_76));
AOI22_X4 i_0_0_267 (.ZN (n_0_0_75), .A1 (\B_r[0] ), .A2 (hfn_ipo_n29), .B1 (drc_ipo_n35), .B2 (n_0_0_143));
NOR2_X1 i_0_0_266 (.ZN (n_0_354), .A1 (n_0_0_141), .A2 (n_0_0_75));
NOR2_X1 i_0_0_265 (.ZN (n_0_353), .A1 (n_0_0_139), .A2 (n_0_0_75));
NOR2_X1 i_0_0_264 (.ZN (n_0_352), .A1 (n_0_0_138), .A2 (n_0_0_75));
NOR2_X1 i_0_0_263 (.ZN (n_0_351), .A1 (n_0_0_137), .A2 (n_0_0_75));
NOR2_X1 i_0_0_262 (.ZN (n_0_350), .A1 (n_0_0_136), .A2 (n_0_0_75));
NOR2_X1 i_0_0_261 (.ZN (n_0_349), .A1 (n_0_0_135), .A2 (n_0_0_75));
NOR2_X1 i_0_0_260 (.ZN (n_0_348), .A1 (n_0_0_134), .A2 (n_0_0_75));
NOR2_X1 i_0_0_259 (.ZN (n_0_347), .A1 (n_0_0_133), .A2 (n_0_0_75));
NOR2_X1 i_0_0_258 (.ZN (n_0_346), .A1 (n_0_0_132), .A2 (n_0_0_75));
NOR2_X1 i_0_0_257 (.ZN (n_0_345), .A1 (n_0_0_131), .A2 (n_0_0_75));
NOR2_X1 i_0_0_256 (.ZN (n_0_344), .A1 (n_0_0_130), .A2 (n_0_0_75));
NOR2_X1 i_0_0_255 (.ZN (n_0_343), .A1 (n_0_0_129), .A2 (n_0_0_75));
NOR2_X1 i_0_0_254 (.ZN (n_0_342), .A1 (n_0_0_128), .A2 (n_0_0_75));
NOR2_X1 i_0_0_253 (.ZN (n_0_341), .A1 (n_0_0_127), .A2 (n_0_0_75));
NOR2_X1 i_0_0_252 (.ZN (n_0_340), .A1 (n_0_0_126), .A2 (n_0_0_75));
NOR2_X1 i_0_0_251 (.ZN (n_0_339), .A1 (n_0_0_125), .A2 (n_0_0_75));
NOR2_X1 i_0_0_250 (.ZN (n_0_338), .A1 (n_0_0_124), .A2 (n_0_0_75));
NOR2_X1 i_0_0_249 (.ZN (n_0_337), .A1 (n_0_0_123), .A2 (n_0_0_75));
NOR2_X1 i_0_0_248 (.ZN (n_0_336), .A1 (n_0_0_122), .A2 (n_0_0_75));
NOR2_X1 i_0_0_247 (.ZN (n_0_335), .A1 (n_0_0_121), .A2 (n_0_0_75));
NOR2_X1 i_0_0_246 (.ZN (n_0_334), .A1 (n_0_0_120), .A2 (n_0_0_75));
NOR2_X1 i_0_0_245 (.ZN (n_0_333), .A1 (n_0_0_119), .A2 (n_0_0_75));
NOR2_X1 i_0_0_244 (.ZN (n_0_332), .A1 (n_0_0_118), .A2 (n_0_0_75));
NOR2_X1 i_0_0_243 (.ZN (n_0_331), .A1 (n_0_0_117), .A2 (n_0_0_75));
NOR2_X1 i_0_0_242 (.ZN (n_0_330), .A1 (n_0_0_116), .A2 (n_0_0_75));
NOR2_X1 i_0_0_241 (.ZN (n_0_329), .A1 (n_0_0_115), .A2 (n_0_0_75));
NOR2_X1 i_0_0_240 (.ZN (n_0_328), .A1 (n_0_0_114), .A2 (n_0_0_75));
NOR2_X1 i_0_0_239 (.ZN (n_0_327), .A1 (n_0_0_113), .A2 (n_0_0_75));
NOR2_X1 i_0_0_238 (.ZN (n_0_326), .A1 (n_0_0_112), .A2 (n_0_0_75));
NOR2_X1 i_0_0_237 (.ZN (n_0_325), .A1 (n_0_0_111), .A2 (n_0_0_75));
NOR2_X1 i_0_0_236 (.ZN (n_0_324), .A1 (n_0_0_110), .A2 (n_0_0_75));
NOR2_X1 i_0_0_235 (.ZN (n_0_323), .A1 (n_0_0_109), .A2 (n_0_0_75));
AND2_X1 i_0_0_234 (.ZN (n_0_322), .A1 (\Accumulator[30] ), .A2 (hfn_ipo_n30));
AND2_X1 i_0_0_233 (.ZN (n_0_321), .A1 (\Accumulator[29] ), .A2 (hfn_ipo_n30));
AND2_X1 i_0_0_232 (.ZN (n_0_320), .A1 (\Accumulator[28] ), .A2 (hfn_ipo_n30));
AND2_X1 i_0_0_231 (.ZN (n_0_319), .A1 (\Accumulator[27] ), .A2 (hfn_ipo_n30));
AND2_X1 i_0_0_230 (.ZN (n_0_318), .A1 (\Accumulator[26] ), .A2 (hfn_ipo_n30));
AND2_X1 i_0_0_229 (.ZN (n_0_317), .A1 (\Accumulator[25] ), .A2 (hfn_ipo_n30));
AND2_X1 i_0_0_228 (.ZN (n_0_316), .A1 (\Accumulator[24] ), .A2 (hfn_ipo_n30));
AND2_X1 i_0_0_227 (.ZN (n_0_315), .A1 (\Accumulator[23] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_226 (.ZN (n_0_314), .A1 (\Accumulator[22] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_225 (.ZN (n_0_313), .A1 (\Accumulator[21] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_224 (.ZN (n_0_312), .A1 (\Accumulator[20] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_223 (.ZN (n_0_311), .A1 (\Accumulator[19] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_222 (.ZN (n_0_310), .A1 (\Accumulator[18] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_221 (.ZN (n_0_309), .A1 (\Accumulator[17] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_220 (.ZN (n_0_308), .A1 (\Accumulator[16] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_219 (.ZN (n_0_307), .A1 (\Accumulator[15] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_218 (.ZN (n_0_306), .A1 (\Accumulator[14] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_217 (.ZN (n_0_305), .A1 (\Accumulator[13] ), .A2 (n_0_0_144));
AND2_X1 i_0_0_216 (.ZN (n_0_304), .A1 (\Accumulator[12] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_215 (.ZN (n_0_303), .A1 (\Accumulator[11] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_214 (.ZN (n_0_302), .A1 (\Accumulator[10] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_213 (.ZN (n_0_301), .A1 (\Accumulator[9] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_212 (.ZN (n_0_300), .A1 (\Accumulator[8] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_211 (.ZN (n_0_299), .A1 (\Accumulator[7] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_210 (.ZN (n_0_298), .A1 (\Accumulator[6] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_209 (.ZN (n_0_297), .A1 (\Accumulator[5] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_208 (.ZN (n_0_296), .A1 (\Accumulator[4] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_207 (.ZN (n_0_295), .A1 (\Accumulator[3] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_206 (.ZN (n_0_294), .A1 (\Accumulator[2] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_205 (.ZN (n_0_293), .A1 (\Accumulator[1] ), .A2 (hfn_ipo_n31));
AND2_X1 i_0_0_204 (.ZN (n_0_292), .A1 (\Accumulator[0] ), .A2 (hfn_ipo_n29));
AND2_X1 i_0_0_203 (.ZN (n_0_291), .A1 (n_0_0_157), .A2 (n_0_63));
NOR2_X1 i_0_0_202 (.ZN (n_0_290), .A1 (hfn_ipo_n23), .A2 (n_0_0_107));
NOR2_X1 i_0_0_201 (.ZN (n_0_289), .A1 (hfn_ipo_n23), .A2 (n_0_0_105));
NOR2_X1 i_0_0_200 (.ZN (CLOCK_slh__n293), .A1 (hfn_ipo_n23), .A2 (n_0_0_104));
NOR2_X1 i_0_0_199 (.ZN (n_0_287), .A1 (hfn_ipo_n23), .A2 (n_0_0_103));
NOR2_X1 i_0_0_198 (.ZN (CLOCK_slh__n299), .A1 (hfn_ipo_n23), .A2 (n_0_0_102));
NOR2_X1 i_0_0_197 (.ZN (CLOCK_slh__n295), .A1 (hfn_ipo_n23), .A2 (n_0_0_101));
NOR2_X1 i_0_0_196 (.ZN (CLOCK_slh__n267), .A1 (hfn_ipo_n23), .A2 (n_0_0_100));
NOR2_X1 i_0_0_195 (.ZN (n_0_283), .A1 (hfn_ipo_n23), .A2 (n_0_0_99));
NOR2_X1 i_0_0_194 (.ZN (n_0_282), .A1 (hfn_ipo_n23), .A2 (n_0_0_98));
NOR2_X1 i_0_0_193 (.ZN (n_0_281), .A1 (hfn_ipo_n23), .A2 (n_0_0_97));
NOR2_X1 i_0_0_192 (.ZN (CLOCK_slh__n277), .A1 (hfn_ipo_n23), .A2 (n_0_0_96));
NOR2_X1 i_0_0_191 (.ZN (CLOCK_slh__n283), .A1 (hfn_ipo_n23), .A2 (n_0_0_95));
NOR2_X1 i_0_0_190 (.ZN (CLOCK_slh__n245), .A1 (hfn_ipo_n23), .A2 (n_0_0_94));
NOR2_X1 i_0_0_189 (.ZN (CLOCK_slh__n249), .A1 (hfn_ipo_n23), .A2 (n_0_0_93));
NOR2_X1 i_0_0_188 (.ZN (CLOCK_slh__n261), .A1 (hfn_ipo_n23), .A2 (n_0_0_92));
NOR2_X1 i_0_0_187 (.ZN (CLOCK_slh__n269), .A1 (hfn_ipo_n23), .A2 (n_0_0_91));
NOR2_X1 i_0_0_186 (.ZN (CLOCK_slh__n253), .A1 (hfn_ipo_n23), .A2 (n_0_0_90));
NOR2_X1 i_0_0_185 (.ZN (CLOCK_slh__n265), .A1 (hfn_ipo_n23), .A2 (n_0_0_89));
NOR2_X1 i_0_0_184 (.ZN (CLOCK_slh__n279), .A1 (hfn_ipo_n23), .A2 (n_0_0_88));
NOR2_X1 i_0_0_183 (.ZN (CLOCK_slh__n300), .A1 (hfn_ipo_n23), .A2 (n_0_0_87));
NOR2_X1 i_0_0_182 (.ZN (CLOCK_slh__n275), .A1 (hfn_ipo_n23), .A2 (n_0_0_86));
NOR2_X1 i_0_0_181 (.ZN (CLOCK_slh__n285), .A1 (hfn_ipo_n23), .A2 (n_0_0_85));
NOR2_X1 i_0_0_180 (.ZN (CLOCK_slh__n289), .A1 (hfn_ipo_n23), .A2 (n_0_0_84));
NOR2_X1 i_0_0_179 (.ZN (CLOCK_slh__n287), .A1 (hfn_ipo_n23), .A2 (n_0_0_83));
NOR2_X1 i_0_0_178 (.ZN (CLOCK_slh__n281), .A1 (hfn_ipo_n23), .A2 (n_0_0_82));
NOR2_X1 i_0_0_177 (.ZN (CLOCK_slh__n263), .A1 (hfn_ipo_n23), .A2 (n_0_0_81));
NOR2_X1 i_0_0_176 (.ZN (CLOCK_slh__n241), .A1 (hfn_ipo_n23), .A2 (n_0_0_80));
NOR2_X1 i_0_0_175 (.ZN (CLOCK_slh__n257), .A1 (hfn_ipo_n23), .A2 (n_0_0_79));
NOR2_X1 i_0_0_174 (.ZN (CLOCK_slh__n291), .A1 (hfn_ipo_n23), .A2 (n_0_0_78));
NOR2_X1 i_0_0_173 (.ZN (CLOCK_slh__n297), .A1 (hfn_ipo_n23), .A2 (n_0_0_77));
NOR2_X1 i_0_0_172 (.ZN (CLOCK_slh__n271), .A1 (hfn_ipo_n23), .A2 (n_0_0_76));
AND2_X1 i_0_0_171 (.ZN (n_0_259), .A1 (n_0_0_157), .A2 (n_0_94));
AND2_X1 i_0_0_170 (.ZN (n_0_258), .A1 (n_0_0_157), .A2 (n_0_93));
AND2_X1 i_0_0_169 (.ZN (n_0_257), .A1 (n_0_0_157), .A2 (n_0_92));
AND2_X1 i_0_0_168 (.ZN (n_0_256), .A1 (n_0_0_157), .A2 (n_0_91));
AND2_X1 i_0_0_167 (.ZN (n_0_255), .A1 (n_0_0_157), .A2 (n_0_90));
AND2_X1 i_0_0_166 (.ZN (n_0_254), .A1 (n_0_0_157), .A2 (n_0_89));
AND2_X1 i_0_0_165 (.ZN (n_0_253), .A1 (n_0_0_157), .A2 (n_0_88));
AND2_X1 i_0_0_164 (.ZN (n_0_252), .A1 (n_0_0_157), .A2 (n_0_87));
AND2_X1 i_0_0_163 (.ZN (n_0_251), .A1 (n_0_0_157), .A2 (n_0_86));
AND2_X1 i_0_0_162 (.ZN (n_0_250), .A1 (n_0_0_157), .A2 (n_0_85));
AND2_X1 i_0_0_161 (.ZN (n_0_249), .A1 (n_0_0_157), .A2 (n_0_84));
AND2_X1 i_0_0_160 (.ZN (n_0_248), .A1 (n_0_0_157), .A2 (n_0_83));
AND2_X1 i_0_0_159 (.ZN (n_0_247), .A1 (n_0_0_157), .A2 (n_0_82));
AND2_X1 i_0_0_158 (.ZN (n_0_246), .A1 (n_0_0_157), .A2 (n_0_81));
AND2_X1 i_0_0_157 (.ZN (n_0_245), .A1 (n_0_0_157), .A2 (n_0_80));
AND2_X1 i_0_0_156 (.ZN (n_0_244), .A1 (n_0_0_157), .A2 (n_0_79));
AND2_X1 i_0_0_155 (.ZN (n_0_243), .A1 (n_0_0_157), .A2 (n_0_78));
AND2_X1 i_0_0_154 (.ZN (n_0_242), .A1 (n_0_0_157), .A2 (n_0_77));
AND2_X1 i_0_0_153 (.ZN (n_0_241), .A1 (n_0_0_157), .A2 (n_0_76));
AND2_X1 i_0_0_152 (.ZN (n_0_240), .A1 (n_0_0_157), .A2 (n_0_75));
AND2_X1 i_0_0_151 (.ZN (n_0_239), .A1 (n_0_0_157), .A2 (n_0_74));
AND2_X1 i_0_0_150 (.ZN (n_0_238), .A1 (n_0_0_157), .A2 (n_0_73));
AND2_X1 i_0_0_149 (.ZN (n_0_237), .A1 (n_0_0_157), .A2 (n_0_72));
AND2_X1 i_0_0_148 (.ZN (n_0_236), .A1 (n_0_0_157), .A2 (n_0_71));
AND2_X1 i_0_0_147 (.ZN (n_0_235), .A1 (n_0_0_157), .A2 (n_0_70));
AND2_X1 i_0_0_146 (.ZN (n_0_234), .A1 (n_0_0_157), .A2 (n_0_69));
AND2_X1 i_0_0_145 (.ZN (n_0_233), .A1 (n_0_0_157), .A2 (n_0_68));
AND2_X1 i_0_0_144 (.ZN (n_0_232), .A1 (n_0_0_157), .A2 (n_0_67));
AND2_X1 i_0_0_143 (.ZN (n_0_231), .A1 (n_0_0_157), .A2 (n_0_66));
AND2_X1 i_0_0_142 (.ZN (n_0_230), .A1 (n_0_0_157), .A2 (n_0_65));
AND2_X1 i_0_0_141 (.ZN (n_0_229), .A1 (n_0_0_157), .A2 (n_0_64));
AND2_X1 i_0_0_139 (.ZN (n_0_228), .A1 (n_0_157), .A2 (hfn_ipo_n28));
AOI22_X1 i_0_0_131 (.ZN (n_0_0_69), .A1 (n_0_153), .A2 (hfn_ipo_n28), .B1 (n_0_91), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_130 (.ZN (n_0_224), .A (n_0_0_69));
AOI22_X1 i_0_0_129 (.ZN (n_0_0_68), .A1 (n_0_152), .A2 (hfn_ipo_n28), .B1 (n_0_90), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_128 (.ZN (n_0_223), .A (n_0_0_68));
AOI22_X1 i_0_0_127 (.ZN (n_0_0_67), .A1 (n_0_151), .A2 (hfn_ipo_n28), .B1 (n_0_89), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_126 (.ZN (n_0_222), .A (n_0_0_67));
AOI22_X1 i_0_0_125 (.ZN (n_0_0_66), .A1 (n_0_150), .A2 (hfn_ipo_n28), .B1 (n_0_88), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_124 (.ZN (n_0_221), .A (n_0_0_66));
AOI22_X1 i_0_0_123 (.ZN (n_0_0_65), .A1 (n_0_149), .A2 (hfn_ipo_n28), .B1 (n_0_87), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_122 (.ZN (n_0_220), .A (n_0_0_65));
AOI22_X1 i_0_0_121 (.ZN (n_0_0_64), .A1 (n_0_148), .A2 (hfn_ipo_n28), .B1 (n_0_86), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_120 (.ZN (n_0_219), .A (n_0_0_64));
AOI22_X1 i_0_0_119 (.ZN (n_0_0_63), .A1 (n_0_147), .A2 (hfn_ipo_n28), .B1 (n_0_85), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_118 (.ZN (n_0_218), .A (n_0_0_63));
AOI22_X1 i_0_0_117 (.ZN (n_0_0_62), .A1 (n_0_146), .A2 (hfn_ipo_n28), .B1 (n_0_84), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_116 (.ZN (n_0_217), .A (n_0_0_62));
AOI22_X1 i_0_0_115 (.ZN (n_0_0_61), .A1 (n_0_145), .A2 (hfn_ipo_n28), .B1 (n_0_83), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_114 (.ZN (n_0_216), .A (n_0_0_61));
AOI22_X1 i_0_0_113 (.ZN (n_0_0_60), .A1 (n_0_144), .A2 (hfn_ipo_n28), .B1 (n_0_82), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_112 (.ZN (n_0_215), .A (n_0_0_60));
AOI22_X1 i_0_0_111 (.ZN (n_0_0_59), .A1 (n_0_143), .A2 (hfn_ipo_n28), .B1 (n_0_81), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_110 (.ZN (n_0_214), .A (n_0_0_59));
AOI22_X1 i_0_0_109 (.ZN (n_0_0_58), .A1 (n_0_142), .A2 (hfn_ipo_n28), .B1 (n_0_80), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_108 (.ZN (n_0_213), .A (n_0_0_58));
AOI22_X1 i_0_0_107 (.ZN (n_0_0_57), .A1 (n_0_141), .A2 (hfn_ipo_n28), .B1 (n_0_79), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_106 (.ZN (n_0_212), .A (n_0_0_57));
AOI22_X1 i_0_0_105 (.ZN (n_0_0_56), .A1 (n_0_140), .A2 (hfn_ipo_n28), .B1 (n_0_78), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_104 (.ZN (n_0_211), .A (n_0_0_56));
AOI22_X1 i_0_0_103 (.ZN (n_0_0_55), .A1 (n_0_139), .A2 (hfn_ipo_n28), .B1 (n_0_77), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_102 (.ZN (n_0_210), .A (n_0_0_55));
AOI22_X1 i_0_0_101 (.ZN (n_0_0_54), .A1 (n_0_138), .A2 (hfn_ipo_n28), .B1 (n_0_76), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_100 (.ZN (n_0_209), .A (n_0_0_54));
AOI22_X1 i_0_0_99 (.ZN (n_0_0_53), .A1 (n_0_137), .A2 (hfn_ipo_n27), .B1 (n_0_75), .B2 (hfn_ipo_n26));
INV_X1 i_0_0_98 (.ZN (n_0_208), .A (n_0_0_53));
AOI22_X1 i_0_0_97 (.ZN (n_0_0_52), .A1 (n_0_136), .A2 (hfn_ipo_n27), .B1 (n_0_74), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_96 (.ZN (n_0_207), .A (n_0_0_52));
AOI22_X1 i_0_0_95 (.ZN (n_0_0_51), .A1 (n_0_135), .A2 (hfn_ipo_n27), .B1 (n_0_73), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_94 (.ZN (n_0_206), .A (n_0_0_51));
AOI22_X1 i_0_0_93 (.ZN (n_0_0_50), .A1 (n_0_134), .A2 (hfn_ipo_n27), .B1 (n_0_72), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_92 (.ZN (n_0_205), .A (n_0_0_50));
AOI22_X1 i_0_0_91 (.ZN (n_0_0_49), .A1 (n_0_133), .A2 (hfn_ipo_n27), .B1 (n_0_71), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_90 (.ZN (n_0_204), .A (n_0_0_49));
AOI22_X1 i_0_0_89 (.ZN (n_0_0_48), .A1 (n_0_132), .A2 (hfn_ipo_n27), .B1 (n_0_70), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_88 (.ZN (n_0_203), .A (n_0_0_48));
AOI22_X1 i_0_0_87 (.ZN (n_0_0_47), .A1 (n_0_131), .A2 (hfn_ipo_n27), .B1 (n_0_69), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_86 (.ZN (n_0_202), .A (n_0_0_47));
AOI22_X1 i_0_0_85 (.ZN (n_0_0_46), .A1 (n_0_130), .A2 (hfn_ipo_n27), .B1 (n_0_68), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_84 (.ZN (n_0_201), .A (n_0_0_46));
AOI22_X1 i_0_0_83 (.ZN (n_0_0_45), .A1 (n_0_129), .A2 (hfn_ipo_n27), .B1 (n_0_67), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_82 (.ZN (n_0_200), .A (n_0_0_45));
AOI22_X1 i_0_0_81 (.ZN (n_0_0_44), .A1 (n_0_128), .A2 (hfn_ipo_n27), .B1 (n_0_66), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_80 (.ZN (n_0_199), .A (n_0_0_44));
AOI22_X1 i_0_0_79 (.ZN (n_0_0_43), .A1 (n_0_127), .A2 (hfn_ipo_n27), .B1 (n_0_65), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_78 (.ZN (n_0_198), .A (n_0_0_43));
AOI22_X1 i_0_0_77 (.ZN (n_0_0_42), .A1 (n_0_126), .A2 (hfn_ipo_n27), .B1 (n_0_64), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_76 (.ZN (n_0_197), .A (n_0_0_42));
AOI22_X1 i_0_0_75 (.ZN (n_0_0_41), .A1 (n_0_125), .A2 (hfn_ipo_n27), .B1 (n_0_63), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_74 (.ZN (n_0_196), .A (n_0_0_41));
AOI22_X1 i_0_0_73 (.ZN (n_0_0_40), .A1 (n_0_124), .A2 (hfn_ipo_n27), .B1 (n_0_385), .B2 (hfn_ipo_n25));
INV_X1 i_0_0_72 (.ZN (n_0_195), .A (n_0_0_40));
AOI22_X1 i_0_0_71 (.ZN (n_0_0_39), .A1 (n_0_384), .A2 (hfn_ipo_n25), .B1 (n_0_123), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_70 (.ZN (n_0_194), .A (n_0_0_39));
AOI22_X1 i_0_0_69 (.ZN (n_0_0_38), .A1 (n_0_383), .A2 (hfn_ipo_n25), .B1 (n_0_122), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_68 (.ZN (n_0_193), .A (n_0_0_38));
AOI22_X1 i_0_0_67 (.ZN (n_0_0_37), .A1 (n_0_382), .A2 (hfn_ipo_n25), .B1 (n_0_121), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_66 (.ZN (n_0_192), .A (n_0_0_37));
AOI22_X1 i_0_0_65 (.ZN (n_0_0_36), .A1 (n_0_381), .A2 (hfn_ipo_n25), .B1 (n_0_120), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_64 (.ZN (n_0_191), .A (n_0_0_36));
AOI22_X1 i_0_0_63 (.ZN (n_0_0_35), .A1 (n_0_380), .A2 (hfn_ipo_n25), .B1 (n_0_119), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_62 (.ZN (n_0_190), .A (n_0_0_35));
AOI22_X1 i_0_0_61 (.ZN (n_0_0_34), .A1 (n_0_379), .A2 (hfn_ipo_n25), .B1 (n_0_118), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_60 (.ZN (n_0_189), .A (n_0_0_34));
AOI22_X1 i_0_0_59 (.ZN (n_0_0_33), .A1 (n_0_378), .A2 (hfn_ipo_n25), .B1 (n_0_117), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_58 (.ZN (n_0_188), .A (n_0_0_33));
AOI22_X1 i_0_0_57 (.ZN (n_0_0_32), .A1 (n_0_377), .A2 (hfn_ipo_n26), .B1 (n_0_116), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_56 (.ZN (n_0_187), .A (n_0_0_32));
AOI22_X1 i_0_0_55 (.ZN (n_0_0_31), .A1 (n_0_376), .A2 (hfn_ipo_n26), .B1 (n_0_115), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_54 (.ZN (n_0_186), .A (n_0_0_31));
AOI22_X1 i_0_0_53 (.ZN (n_0_0_30), .A1 (n_0_375), .A2 (hfn_ipo_n26), .B1 (n_0_114), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_52 (.ZN (n_0_185), .A (n_0_0_30));
AOI22_X1 i_0_0_51 (.ZN (n_0_0_29), .A1 (n_0_374), .A2 (hfn_ipo_n26), .B1 (n_0_113), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_50 (.ZN (n_0_184), .A (n_0_0_29));
AOI22_X1 i_0_0_49 (.ZN (n_0_0_28), .A1 (n_0_373), .A2 (hfn_ipo_n26), .B1 (n_0_112), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_48 (.ZN (n_0_183), .A (n_0_0_28));
AOI22_X1 i_0_0_47 (.ZN (n_0_0_27), .A1 (n_0_372), .A2 (hfn_ipo_n26), .B1 (n_0_111), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_46 (.ZN (n_0_182), .A (n_0_0_27));
AOI22_X1 i_0_0_45 (.ZN (n_0_0_26), .A1 (n_0_371), .A2 (hfn_ipo_n26), .B1 (n_0_110), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_44 (.ZN (n_0_181), .A (n_0_0_26));
AOI22_X1 i_0_0_43 (.ZN (n_0_0_25), .A1 (n_0_370), .A2 (hfn_ipo_n26), .B1 (n_0_109), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_42 (.ZN (n_0_180), .A (n_0_0_25));
AOI22_X1 i_0_0_41 (.ZN (n_0_0_24), .A1 (n_0_369), .A2 (hfn_ipo_n26), .B1 (n_0_108), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_40 (.ZN (n_0_179), .A (n_0_0_24));
AOI22_X1 i_0_0_39 (.ZN (n_0_0_23), .A1 (n_0_368), .A2 (hfn_ipo_n26), .B1 (n_0_107), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_38 (.ZN (n_0_178), .A (n_0_0_23));
AOI22_X1 i_0_0_37 (.ZN (n_0_0_22), .A1 (n_0_367), .A2 (hfn_ipo_n26), .B1 (n_0_106), .B2 (hfn_ipo_n28));
INV_X1 i_0_0_36 (.ZN (n_0_177), .A (n_0_0_22));
AOI22_X1 i_0_0_35 (.ZN (n_0_0_21), .A1 (n_0_366), .A2 (hfn_ipo_n25), .B1 (n_0_105), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_34 (.ZN (n_0_176), .A (n_0_0_21));
AOI22_X1 i_0_0_33 (.ZN (n_0_0_20), .A1 (n_0_365), .A2 (hfn_ipo_n25), .B1 (n_0_104), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_32 (.ZN (n_0_175), .A (n_0_0_20));
AOI22_X1 i_0_0_31 (.ZN (n_0_0_19), .A1 (n_0_364), .A2 (hfn_ipo_n25), .B1 (n_0_103), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_30 (.ZN (n_0_174), .A (n_0_0_19));
AOI22_X1 i_0_0_29 (.ZN (n_0_0_18), .A1 (n_0_363), .A2 (hfn_ipo_n25), .B1 (n_0_102), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_28 (.ZN (n_0_173), .A (n_0_0_18));
AOI22_X1 i_0_0_27 (.ZN (n_0_0_17), .A1 (n_0_362), .A2 (hfn_ipo_n25), .B1 (n_0_101), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_26 (.ZN (n_0_172), .A (n_0_0_17));
AOI22_X1 i_0_0_25 (.ZN (n_0_0_16), .A1 (n_0_361), .A2 (hfn_ipo_n25), .B1 (n_0_100), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_24 (.ZN (n_0_171), .A (n_0_0_16));
AOI22_X1 i_0_0_23 (.ZN (n_0_0_15), .A1 (n_0_360), .A2 (hfn_ipo_n25), .B1 (n_0_99), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_22 (.ZN (n_0_170), .A (n_0_0_15));
AOI22_X1 i_0_0_21 (.ZN (n_0_0_14), .A1 (n_0_359), .A2 (hfn_ipo_n25), .B1 (n_0_98), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_20 (.ZN (n_0_169), .A (n_0_0_14));
AOI22_X1 i_0_0_19 (.ZN (n_0_0_13), .A1 (n_0_358), .A2 (hfn_ipo_n25), .B1 (n_0_97), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_18 (.ZN (n_0_168), .A (n_0_0_13));
AOI22_X1 i_0_0_17 (.ZN (n_0_0_12), .A1 (n_0_357), .A2 (hfn_ipo_n25), .B1 (n_0_96), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_16 (.ZN (n_0_167), .A (n_0_0_12));
AOI22_X1 i_0_0_15 (.ZN (n_0_0_11), .A1 (n_0_356), .A2 (hfn_ipo_n25), .B1 (n_0_95), .B2 (hfn_ipo_n27));
INV_X1 i_0_0_14 (.ZN (n_0_166), .A (n_0_0_11));
AOI221_X1 i_0_0_13 (.ZN (n_0_0_10), .A (hfn_ipo_n30), .B1 (drc_ipo_n98), .B2 (n_0_0_154)
    , .C1 (n_0_0_155), .C2 (drc_ipo_n66));
AOI211_X1 i_0_0_12 (.ZN (n_0_165), .A (n_0_0_10), .B (hfn_ipo_n23), .C1 (n_0_0_153), .C2 (hfn_ipo_n30));
AOI221_X1 i_0_0_11 (.ZN (n_0_164), .A (n_0_418), .B1 (n_0_0_156), .B2 (n_0_0_152)
    , .C1 (\counter[6] ), .C2 (n_0_0_4));
AND2_X1 i_0_0_10 (.ZN (n_0_163), .A1 (n_0_0_9), .A2 (n_0_0_147));
AND2_X1 i_0_0_9 (.ZN (n_0_162), .A1 (n_0_0_8), .A2 (n_0_0_147));
AND2_X1 i_0_0_8 (.ZN (n_0_161), .A1 (n_0_0_7), .A2 (n_0_0_147));
AND2_X1 i_0_0_7 (.ZN (n_0_160), .A1 (n_0_0_6), .A2 (n_0_0_147));
AND2_X1 i_0_0_6 (.ZN (n_0_159), .A1 (n_0_0_5), .A2 (n_0_0_147));
NOR2_X1 i_0_0_5 (.ZN (n_0_158), .A1 (hfn_ipo_n23), .A2 (\counter[0] ));
HA_X1 i_0_0_4 (.CO (n_0_0_4), .S (n_0_0_9), .A (\counter[5] ), .B (n_0_0_3));
HA_X1 i_0_0_3 (.CO (n_0_0_3), .S (n_0_0_8), .A (\counter[4] ), .B (n_0_0_2));
HA_X1 i_0_0_2 (.CO (n_0_0_2), .S (n_0_0_7), .A (\counter[3] ), .B (n_0_0_1));
HA_X1 i_0_0_1 (.CO (n_0_0_1), .S (n_0_0_6), .A (\counter[2] ), .B (n_0_0_0));
HA_X1 i_0_0_0 (.CO (n_0_0_0), .S (n_0_0_5), .A (\counter[1] ), .B (\counter[0] ));
datapath__0_9 i_0_11 (.p_1 ({n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, 
    n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, 
    n_0_142, n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, 
    n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, 
    n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, 
    n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, 
    n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, 
    n_0_97, n_0_96, n_0_95, uc_4}), .p_0 ({uc_3, n_0_94, n_0_93, n_0_92, n_0_91, 
    n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, 
    n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, 
    n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_385, n_0_384, 
    n_0_383, n_0_382, n_0_381, n_0_380, n_0_379, n_0_378, n_0_377, n_0_376, n_0_375, 
    n_0_374, n_0_373, n_0_372, n_0_371, n_0_370, n_0_369, n_0_368, n_0_367, n_0_366, 
    n_0_365, n_0_364, n_0_363, n_0_362, n_0_361, n_0_360, n_0_359, n_0_358, n_0_357, 
    n_0_356, n_0_355}));
datapath__0_6 i_0_8 (.Accumulator1 ({n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, 
    n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, 
    n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, 
    n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63}), .Accumulator ({uc_2, n_0_322, 
    n_0_321, n_0_320, n_0_319, n_0_318, n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, 
    n_0_312, n_0_311, n_0_310, n_0_309, n_0_308, n_0_307, n_0_306, n_0_305, n_0_304, 
    n_0_303, n_0_302, n_0_301, n_0_300, n_0_299, n_0_298, n_0_297, n_0_296, n_0_295, 
    n_0_294, n_0_293, n_0_292}), .p_0 ({n_0_354, n_0_353, n_0_352, n_0_351, n_0_350, 
    n_0_349, n_0_348, n_0_347, n_0_346, n_0_345, n_0_344, n_0_343, n_0_342, n_0_341, 
    n_0_340, n_0_339, n_0_338, n_0_337, n_0_336, n_0_335, n_0_334, n_0_333, n_0_332, 
    n_0_331, n_0_330, n_0_329, n_0_328, n_0_327, n_0_326, n_0_325, n_0_324, n_0_323}));
datapath__0_2 i_0_4 (.p_0 ({n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, 
    n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, 
    n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, 
    n_0_35, n_0_34, n_0_33, n_0_32, uc_1}), .b ({drc_ipo_n66, drc_ipo_n65, drc_ipo_n64, 
    drc_ipo_n63, drc_ipo_n62, drc_ipo_n61, drc_ipo_n60, drc_ipo_n59, drc_ipo_n58, 
    drc_ipo_n57, drc_ipo_n56, drc_ipo_n55, drc_ipo_n54, drc_ipo_n53, drc_ipo_n52, 
    drc_ipo_n51, drc_ipo_n50, drc_ipo_n49, drc_ipo_n48, drc_ipo_n47, drc_ipo_n46, 
    drc_ipo_n45, drc_ipo_n44, drc_ipo_n43, drc_ipo_n42, drc_ipo_n41, drc_ipo_n40, 
    drc_ipo_n39, drc_ipo_n38, drc_ipo_n37, drc_ipo_n36, drc_ipo_n35}));
datapath i_0_1 (.p_0 ({n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, 
    n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, 
    n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, 
    n_0_2, n_0_1, uc_0}), .a ({drc_ipo_n98, drc_ipo_n97, drc_ipo_n96, drc_ipo_n95, 
    drc_ipo_n94, drc_ipo_n93, drc_ipo_n92, drc_ipo_n91, drc_ipo_n90, drc_ipo_n89, 
    drc_ipo_n88, drc_ipo_n87, drc_ipo_n86, drc_ipo_n85, drc_ipo_n84, drc_ipo_n83, 
    drc_ipo_n82, drc_ipo_n81, drc_ipo_n80, drc_ipo_n79, drc_ipo_n78, drc_ipo_n77, 
    drc_ipo_n76, drc_ipo_n75, drc_ipo_n74, drc_ipo_n73, drc_ipo_n72, drc_ipo_n71, 
    drc_ipo_n70, drc_ipo_n69, drc_ipo_n68, drc_ipo_n67}));
DFF_X1 \c_reg[0]  (.Q (c[0]), .CK (CTS_n_tid1_120), .D (n_0_260));
DFF_X1 \c_reg[1]  (.Q (c[1]), .CK (CTS_n_tid1_120), .D (n_0_166));
DFF_X1 \c_reg[2]  (.Q (c[2]), .CK (CTS_n_tid1_120), .D (n_0_167));
DFF_X1 \c_reg[3]  (.Q (c[3]), .CK (CTS_n_tid1_120), .D (n_0_168));
DFF_X1 \c_reg[4]  (.Q (c[4]), .CK (CTS_n_tid1_120), .D (n_0_169));
DFF_X1 \c_reg[5]  (.Q (c[5]), .CK (CTS_n_tid1_120), .D (n_0_170));
DFF_X1 \c_reg[6]  (.Q (c[6]), .CK (CTS_n_tid1_120), .D (n_0_171));
DFF_X1 \c_reg[7]  (.Q (c[7]), .CK (CTS_n_tid1_120), .D (n_0_172));
DFF_X1 \c_reg[8]  (.Q (c[8]), .CK (CTS_n_tid1_120), .D (n_0_173));
DFF_X1 \c_reg[9]  (.Q (c[9]), .CK (CTS_n_tid1_120), .D (n_0_174));
DFF_X1 \c_reg[10]  (.Q (c[10]), .CK (CTS_n_tid1_120), .D (n_0_175));
DFF_X1 \c_reg[11]  (.Q (c[11]), .CK (CTS_n_tid1_120), .D (n_0_176));
DFF_X1 \c_reg[12]  (.Q (c[12]), .CK (CTS_n_tid1_120), .D (n_0_177));
DFF_X1 \c_reg[13]  (.Q (c[13]), .CK (CTS_n_tid1_120), .D (n_0_178));
DFF_X1 \c_reg[14]  (.Q (c[14]), .CK (CTS_n_tid1_120), .D (n_0_179));
DFF_X1 \c_reg[15]  (.Q (c[15]), .CK (CTS_n_tid1_120), .D (n_0_180));
DFF_X1 \c_reg[16]  (.Q (c[16]), .CK (CTS_n_tid1_120), .D (n_0_181));
DFF_X1 \c_reg[17]  (.Q (c[17]), .CK (CTS_n_tid1_120), .D (n_0_182));
DFF_X1 \c_reg[18]  (.Q (c[18]), .CK (CTS_n_tid1_120), .D (n_0_183));
DFF_X1 \c_reg[19]  (.Q (c[19]), .CK (CTS_n_tid1_120), .D (n_0_184));
DFF_X1 \c_reg[20]  (.Q (c[20]), .CK (CTS_n_tid1_120), .D (n_0_185));
DFF_X1 \c_reg[21]  (.Q (c[21]), .CK (CTS_n_tid1_120), .D (n_0_186));
DFF_X1 \c_reg[22]  (.Q (c[22]), .CK (CTS_n_tid1_120), .D (n_0_187));
DFF_X1 \c_reg[23]  (.Q (c[23]), .CK (CTS_n_tid1_120), .D (n_0_188));
DFF_X1 \c_reg[24]  (.Q (c[24]), .CK (CTS_n_tid1_120), .D (n_0_189));
DFF_X1 \c_reg[25]  (.Q (c[25]), .CK (CTS_n_tid1_120), .D (n_0_190));
DFF_X1 \c_reg[26]  (.Q (c[26]), .CK (CTS_n_tid1_120), .D (n_0_191));
DFF_X1 \c_reg[27]  (.Q (c[27]), .CK (CTS_n_tid1_120), .D (n_0_192));
DFF_X1 \c_reg[28]  (.Q (c[28]), .CK (CTS_n_tid1_120), .D (n_0_193));
DFF_X1 \c_reg[29]  (.Q (c[29]), .CK (CTS_n_tid1_120), .D (n_0_194));
DFF_X1 \c_reg[30]  (.Q (c[30]), .CK (CTS_n_tid1_120), .D (n_0_195));
DFF_X1 \c_reg[31]  (.Q (c[31]), .CK (CTS_n_tid1_120), .D (n_0_196));
DFF_X1 \c_reg[32]  (.Q (c[32]), .CK (CTS_n_tid1_120), .D (n_0_197));
DFF_X1 \c_reg[33]  (.Q (c[33]), .CK (CTS_n_tid1_120), .D (n_0_198));
DFF_X1 \c_reg[34]  (.Q (c[34]), .CK (CTS_n_tid1_120), .D (n_0_199));
DFF_X1 \c_reg[35]  (.Q (c[35]), .CK (CTS_n_tid1_120), .D (n_0_200));
DFF_X1 \c_reg[36]  (.Q (c[36]), .CK (CTS_n_tid1_120), .D (n_0_201));
DFF_X1 \c_reg[37]  (.Q (c[37]), .CK (CTS_n_tid1_120), .D (n_0_202));
DFF_X1 \c_reg[38]  (.Q (c[38]), .CK (CTS_n_tid1_120), .D (n_0_203));
DFF_X1 \c_reg[39]  (.Q (c[39]), .CK (CTS_n_tid1_120), .D (n_0_204));
DFF_X1 \c_reg[40]  (.Q (c[40]), .CK (CTS_n_tid1_120), .D (n_0_205));
DFF_X1 \c_reg[41]  (.Q (c[41]), .CK (CTS_n_tid1_120), .D (n_0_206));
DFF_X1 \c_reg[42]  (.Q (c[42]), .CK (CTS_n_tid1_120), .D (n_0_207));
DFF_X1 \c_reg[43]  (.Q (c[43]), .CK (CTS_n_tid1_120), .D (n_0_208));
DFF_X1 \c_reg[44]  (.Q (c[44]), .CK (CTS_n_tid1_120), .D (n_0_209));
DFF_X1 \c_reg[45]  (.Q (c[45]), .CK (CTS_n_tid1_120), .D (n_0_210));
DFF_X1 \c_reg[46]  (.Q (c[46]), .CK (CTS_n_tid1_120), .D (n_0_211));
DFF_X1 \c_reg[47]  (.Q (c[47]), .CK (CTS_n_tid1_120), .D (n_0_212));
DFF_X1 \c_reg[48]  (.Q (c[48]), .CK (CTS_n_tid1_120), .D (n_0_213));
DFF_X1 \c_reg[49]  (.Q (c[49]), .CK (CTS_n_tid1_120), .D (n_0_214));
DFF_X1 \c_reg[50]  (.Q (c[50]), .CK (CTS_n_tid1_120), .D (n_0_215));
DFF_X1 \c_reg[51]  (.Q (c[51]), .CK (CTS_n_tid1_120), .D (n_0_216));
DFF_X1 \c_reg[52]  (.Q (c[52]), .CK (CTS_n_tid1_120), .D (n_0_217));
DFF_X1 \c_reg[53]  (.Q (c[53]), .CK (CTS_n_tid1_120), .D (n_0_218));
DFF_X1 \c_reg[54]  (.Q (c[54]), .CK (CTS_n_tid1_120), .D (n_0_219));
DFF_X1 \c_reg[55]  (.Q (c[55]), .CK (CTS_n_tid1_120), .D (n_0_220));
DFF_X1 \c_reg[56]  (.Q (c[56]), .CK (CTS_n_tid1_120), .D (n_0_221));
DFF_X1 \c_reg[57]  (.Q (c[57]), .CK (CTS_n_tid1_120), .D (n_0_222));
DFF_X1 \c_reg[58]  (.Q (c[58]), .CK (CTS_n_tid1_120), .D (n_0_223));
DFF_X1 \c_reg[59]  (.Q (c[59]), .CK (CTS_n_tid1_120), .D (n_0_224));
DFF_X1 \c_reg[60]  (.Q (c[60]), .CK (CTS_n_tid1_120), .D (n_0_225));
DFF_X1 \c_reg[61]  (.Q (c[61]), .CK (CTS_n_tid1_120), .D (n_0_226));
DFF_X1 \c_reg[62]  (.Q (c[62]), .CK (CTS_n_tid1_120), .D (n_0_227));
DFF_X1 \c_reg[63]  (.Q (c[63]), .CK (CTS_n_tid1_120), .D (n_0_228));
CLKGATETST_X8 clk_gate_c_reg (.GCK (CTS_n_tid1_121), .CK (CTS_n_tid0_170), .E (n_0_418), .SE (1'b0 ));
BUF_X4 hfn_ipo_c23 (.Z (hfn_ipo_n23), .A (drc_ipo_n99));
BUF_X4 hfn_ipo_c24 (.Z (hfn_ipo_n24), .A (drc_ipo_n99));
CLKBUF_X2 hfn_ipo_c26 (.Z (hfn_ipo_n26), .A (n_0_0_73));
CLKBUF_X2 hfn_ipo_c27 (.Z (hfn_ipo_n27), .A (n_0_0_74));
CLKBUF_X2 hfn_ipo_c28 (.Z (hfn_ipo_n28), .A (n_0_0_74));
CLKBUF_X2 hfn_ipo_c29 (.Z (hfn_ipo_n29), .A (n_0_0_144));
CLKBUF_X2 hfn_ipo_c30 (.Z (hfn_ipo_n30), .A (n_0_0_144));
BUF_X1 hfn_ipo_c31 (.Z (hfn_ipo_n31), .A (n_0_0_144));
CLKBUF_X2 CTS_L2_c_tid0_150 (.Z (CTS_n_tid0_168), .A (CTS_n_tid0_170));
CLKBUF_X3 CTS_L3_c_tid1_121 (.Z (CTS_n_tid1_120), .A (CTS_n_tid1_121));
CLKBUF_X2 hfn_ipo_c25 (.Z (hfn_ipo_n25), .A (n_0_0_73));
CLKBUF_X2 CTS_L2_c_tid0_151 (.Z (CTS_n_tid0_169), .A (CTS_n_tid0_170));
CLKBUF_X1 drc_ipo_c35 (.Z (drc_ipo_n35), .A (b[0]));
CLKBUF_X1 drc_ipo_c36 (.Z (drc_ipo_n36), .A (b[1]));
CLKBUF_X1 drc_ipo_c37 (.Z (drc_ipo_n37), .A (b[2]));
CLKBUF_X1 drc_ipo_c38 (.Z (drc_ipo_n38), .A (b[3]));
CLKBUF_X1 drc_ipo_c39 (.Z (drc_ipo_n39), .A (b[4]));
CLKBUF_X1 drc_ipo_c40 (.Z (drc_ipo_n40), .A (b[5]));
CLKBUF_X1 drc_ipo_c41 (.Z (drc_ipo_n41), .A (b[6]));
CLKBUF_X1 drc_ipo_c42 (.Z (drc_ipo_n42), .A (b[7]));
CLKBUF_X1 drc_ipo_c43 (.Z (drc_ipo_n43), .A (b[8]));
CLKBUF_X1 drc_ipo_c44 (.Z (drc_ipo_n44), .A (b[9]));
CLKBUF_X1 drc_ipo_c45 (.Z (drc_ipo_n45), .A (b[10]));
CLKBUF_X1 drc_ipo_c46 (.Z (drc_ipo_n46), .A (b[11]));
CLKBUF_X1 drc_ipo_c47 (.Z (drc_ipo_n47), .A (b[12]));
CLKBUF_X1 drc_ipo_c48 (.Z (drc_ipo_n48), .A (b[13]));
CLKBUF_X1 drc_ipo_c49 (.Z (drc_ipo_n49), .A (b[14]));
CLKBUF_X1 drc_ipo_c50 (.Z (drc_ipo_n50), .A (b[15]));
CLKBUF_X1 drc_ipo_c51 (.Z (drc_ipo_n51), .A (b[16]));
CLKBUF_X1 drc_ipo_c52 (.Z (drc_ipo_n52), .A (b[17]));
CLKBUF_X1 drc_ipo_c53 (.Z (drc_ipo_n53), .A (b[18]));
CLKBUF_X1 drc_ipo_c54 (.Z (drc_ipo_n54), .A (b[19]));
CLKBUF_X1 drc_ipo_c55 (.Z (drc_ipo_n55), .A (b[20]));
CLKBUF_X1 drc_ipo_c56 (.Z (drc_ipo_n56), .A (b[21]));
CLKBUF_X1 drc_ipo_c57 (.Z (drc_ipo_n57), .A (b[22]));
CLKBUF_X1 drc_ipo_c58 (.Z (drc_ipo_n58), .A (b[23]));
CLKBUF_X1 drc_ipo_c59 (.Z (drc_ipo_n59), .A (b[24]));
CLKBUF_X1 drc_ipo_c60 (.Z (drc_ipo_n60), .A (b[25]));
CLKBUF_X1 drc_ipo_c61 (.Z (drc_ipo_n61), .A (b[26]));
CLKBUF_X1 drc_ipo_c62 (.Z (drc_ipo_n62), .A (b[27]));
CLKBUF_X1 drc_ipo_c63 (.Z (drc_ipo_n63), .A (b[28]));
CLKBUF_X1 drc_ipo_c64 (.Z (drc_ipo_n64), .A (b[29]));
CLKBUF_X1 drc_ipo_c65 (.Z (drc_ipo_n65), .A (b[30]));
CLKBUF_X1 drc_ipo_c66 (.Z (drc_ipo_n66), .A (b[31]));
CLKBUF_X1 drc_ipo_c67 (.Z (drc_ipo_n67), .A (a[0]));
CLKBUF_X1 drc_ipo_c68 (.Z (drc_ipo_n68), .A (a[1]));
CLKBUF_X1 drc_ipo_c69 (.Z (drc_ipo_n69), .A (a[2]));
CLKBUF_X1 drc_ipo_c70 (.Z (drc_ipo_n70), .A (a[3]));
CLKBUF_X1 drc_ipo_c71 (.Z (drc_ipo_n71), .A (a[4]));
CLKBUF_X1 drc_ipo_c72 (.Z (drc_ipo_n72), .A (a[5]));
CLKBUF_X1 drc_ipo_c73 (.Z (drc_ipo_n73), .A (a[6]));
CLKBUF_X1 drc_ipo_c74 (.Z (drc_ipo_n74), .A (a[7]));
CLKBUF_X1 drc_ipo_c75 (.Z (drc_ipo_n75), .A (a[8]));
CLKBUF_X1 drc_ipo_c76 (.Z (drc_ipo_n76), .A (a[9]));
CLKBUF_X1 drc_ipo_c77 (.Z (drc_ipo_n77), .A (a[10]));
CLKBUF_X1 drc_ipo_c78 (.Z (drc_ipo_n78), .A (a[11]));
CLKBUF_X1 drc_ipo_c79 (.Z (drc_ipo_n79), .A (a[12]));
CLKBUF_X1 drc_ipo_c80 (.Z (drc_ipo_n80), .A (a[13]));
CLKBUF_X1 drc_ipo_c81 (.Z (drc_ipo_n81), .A (a[14]));
CLKBUF_X1 drc_ipo_c82 (.Z (drc_ipo_n82), .A (a[15]));
CLKBUF_X1 drc_ipo_c83 (.Z (drc_ipo_n83), .A (a[16]));
CLKBUF_X1 drc_ipo_c84 (.Z (drc_ipo_n84), .A (a[17]));
CLKBUF_X1 drc_ipo_c85 (.Z (drc_ipo_n85), .A (a[18]));
CLKBUF_X1 drc_ipo_c86 (.Z (drc_ipo_n86), .A (a[19]));
CLKBUF_X1 drc_ipo_c87 (.Z (drc_ipo_n87), .A (a[20]));
CLKBUF_X1 drc_ipo_c88 (.Z (drc_ipo_n88), .A (a[21]));
CLKBUF_X1 drc_ipo_c89 (.Z (drc_ipo_n89), .A (a[22]));
CLKBUF_X1 drc_ipo_c90 (.Z (drc_ipo_n90), .A (a[23]));
CLKBUF_X1 drc_ipo_c91 (.Z (drc_ipo_n91), .A (a[24]));
CLKBUF_X1 drc_ipo_c92 (.Z (drc_ipo_n92), .A (a[25]));
CLKBUF_X1 drc_ipo_c93 (.Z (drc_ipo_n93), .A (a[26]));
CLKBUF_X1 drc_ipo_c94 (.Z (drc_ipo_n94), .A (a[27]));
CLKBUF_X1 drc_ipo_c95 (.Z (drc_ipo_n95), .A (a[28]));
CLKBUF_X1 drc_ipo_c96 (.Z (drc_ipo_n96), .A (a[29]));
CLKBUF_X1 drc_ipo_c97 (.Z (drc_ipo_n97), .A (a[30]));
CLKBUF_X1 drc_ipo_c98 (.Z (drc_ipo_n98), .A (a[31]));
BUF_X4 drc_ipo_c99 (.Z (drc_ipo_n99), .A (rst));
CLKBUF_X1 CTS_L1_c_tid0_152 (.Z (CTS_n_tid0_170), .A (clk));
CLKBUF_X1 CLOCK_slh__c177 (.Z (CLOCK_slh__n242), .A (CLOCK_slh__n241));
CLKBUF_X1 CLOCK_slh__c178 (.Z (n_0_264), .A (CLOCK_slh__n242));
CLKBUF_X1 CLOCK_slh__c181 (.Z (CLOCK_slh__n246), .A (CLOCK_slh__n245));
CLKBUF_X1 CLOCK_slh__c182 (.Z (n_0_278), .A (CLOCK_slh__n246));
CLKBUF_X1 CLOCK_slh__c185 (.Z (CLOCK_slh__n250), .A (CLOCK_slh__n249));
CLKBUF_X1 CLOCK_slh__c186 (.Z (n_0_277), .A (CLOCK_slh__n250));
CLKBUF_X1 CLOCK_slh__c189 (.Z (CLOCK_slh__n254), .A (CLOCK_slh__n253));
CLKBUF_X1 CLOCK_slh__c190 (.Z (n_0_274), .A (CLOCK_slh__n254));
CLKBUF_X1 CLOCK_slh__c193 (.Z (CLOCK_slh__n258), .A (CLOCK_slh__n257));
CLKBUF_X1 CLOCK_slh__c194 (.Z (n_0_263), .A (CLOCK_slh__n258));
CLKBUF_X1 CLOCK_slh__c197 (.Z (n_0_276), .A (CLOCK_slh__n261));
CLKBUF_X1 CLOCK_slh__c199 (.Z (n_0_265), .A (CLOCK_slh__n263));
CLKBUF_X1 CLOCK_slh__c201 (.Z (n_0_273), .A (CLOCK_slh__n265));
CLKBUF_X1 CLOCK_slh__c203 (.Z (n_0_284), .A (CLOCK_slh__n267));
CLKBUF_X1 CLOCK_slh__c205 (.Z (n_0_275), .A (CLOCK_slh__n269));
CLKBUF_X1 CLOCK_slh__c207 (.Z (n_0_260), .A (CLOCK_slh__n271));
CLKBUF_X1 CLOCK_slh__c209 (.Z (n_0_386), .A (CLOCK_slh__n273));
CLKBUF_X1 CLOCK_slh__c211 (.Z (n_0_270), .A (CLOCK_slh__n275));
CLKBUF_X1 CLOCK_slh__c213 (.Z (n_0_280), .A (CLOCK_slh__n277));
CLKBUF_X1 CLOCK_slh__c215 (.Z (n_0_272), .A (CLOCK_slh__n279));
CLKBUF_X1 CLOCK_slh__c217 (.Z (n_0_266), .A (CLOCK_slh__n281));
CLKBUF_X1 CLOCK_slh__c219 (.Z (n_0_279), .A (CLOCK_slh__n283));
CLKBUF_X1 CLOCK_slh__c221 (.Z (n_0_269), .A (CLOCK_slh__n285));
CLKBUF_X1 CLOCK_slh__c223 (.Z (n_0_267), .A (CLOCK_slh__n287));
CLKBUF_X1 CLOCK_slh__c225 (.Z (n_0_268), .A (CLOCK_slh__n289));
CLKBUF_X1 CLOCK_slh__c227 (.Z (n_0_262), .A (CLOCK_slh__n291));
CLKBUF_X1 CLOCK_slh__c229 (.Z (n_0_288), .A (CLOCK_slh__n293));
CLKBUF_X1 CLOCK_slh__c231 (.Z (n_0_285), .A (CLOCK_slh__n295));
CLKBUF_X1 CLOCK_slh__c233 (.Z (n_0_261), .A (CLOCK_slh__n297));
CLKBUF_X1 CLOCK_slh__c235 (.Z (n_0_286), .A (CLOCK_slh__n299));
CLKBUF_X1 CLOCK_slh__c236 (.Z (n_0_271), .A (CLOCK_slh__n300));

endmodule //seq_multiplier


