
// 	Tue Jan  3 14:18:07 2023
//	vlsi
//	localhost.localdomain

module datapath (p_0, Accumulator, Accumulator1);

output [23:0] Accumulator1;
input [23:0] Accumulator;
input [23:0] p_0;
wire n_0;
wire n_98;
wire n_1;
wire n_97;
wire n_96;
wire n_2;
wire n_100;
wire n_94;
wire n_3;
wire n_93;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_90;
wire n_81;
wire n_11;
wire n_5;
wire n_91;
wire n_85;
wire n_8;
wire n_88;
wire n_86;
wire n_92;
wire n_83;
wire n_79;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_76;
wire n_67;
wire n_19;
wire n_13;
wire n_77;
wire n_71;
wire n_16;
wire n_74;
wire n_72;
wire n_78;
wire n_69;
wire n_65;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_62;
wire n_53;
wire n_27;
wire n_21;
wire n_63;
wire n_57;
wire n_24;
wire n_60;
wire n_58;
wire n_64;
wire n_55;
wire n_51;
wire n_34;
wire n_33;
wire n_31;
wire n_29;
wire n_28;
wire n_108;
wire n_32;
wire n_103;
wire n_35;
wire n_30;
wire n_107;
wire n_49;
wire n_105;
wire n_109;
wire n_47;
wire n_39;
wire n_37;
wire n_36;
wire n_112;
wire n_45;
wire n_43;
wire n_40;
wire n_38;
wire n_110;
wire n_111;
wire n_115;
wire n_114;
wire n_113;
wire n_41;
wire n_42;
wire n_44;
wire n_46;
wire n_102;
wire n_50;
wire n_48;
wire n_106;
wire n_52;
wire n_56;
wire n_59;
wire n_54;
wire n_61;
wire n_66;
wire n_70;
wire n_73;
wire n_68;
wire n_75;
wire n_80;
wire n_84;
wire n_87;
wire n_82;
wire n_89;
wire n_101;
wire n_95;
wire n_99;
wire n_104;


INV_X1 i_139 (.ZN (n_115), .A (p_0[20]));
INV_X1 i_138 (.ZN (n_114), .A (Accumulator[20]));
NOR2_X1 i_137 (.ZN (n_113), .A1 (p_0[22]), .A2 (Accumulator[22]));
NOR2_X1 i_136 (.ZN (n_112), .A1 (p_0[20]), .A2 (Accumulator[20]));
INV_X1 i_135 (.ZN (n_111), .A (n_112));
OAI21_X1 i_134 (.ZN (n_110), .A (n_111), .B1 (p_0[21]), .B2 (Accumulator[21]));
NOR2_X1 i_133 (.ZN (n_109), .A1 (p_0[19]), .A2 (Accumulator[19]));
NOR2_X1 i_132 (.ZN (n_108), .A1 (p_0[17]), .A2 (Accumulator[17]));
OAI22_X1 i_131 (.ZN (n_107), .A1 (p_0[17]), .A2 (Accumulator[17]), .B1 (p_0[18]), .B2 (Accumulator[18]));
OR2_X1 i_130 (.ZN (n_106), .A1 (n_109), .A2 (n_107));
NAND2_X1 i_129 (.ZN (n_105), .A1 (p_0[16]), .A2 (Accumulator[16]));
AOI22_X1 i_128 (.ZN (n_104), .A1 (p_0[16]), .A2 (Accumulator[16]), .B1 (p_0[17]), .B2 (Accumulator[17]));
NAND2_X1 i_127 (.ZN (n_103), .A1 (p_0[18]), .A2 (Accumulator[18]));
OAI22_X1 i_126 (.ZN (n_102), .A1 (n_106), .A2 (n_104), .B1 (n_109), .B2 (n_103));
AND2_X1 i_125 (.ZN (n_101), .A1 (p_0[3]), .A2 (Accumulator[3]));
NAND2_X1 i_124 (.ZN (n_100), .A1 (p_0[2]), .A2 (Accumulator[2]));
NOR2_X1 i_123 (.ZN (n_99), .A1 (p_0[1]), .A2 (Accumulator[1]));
NAND2_X1 i_122 (.ZN (n_98), .A1 (p_0[0]), .A2 (Accumulator[0]));
NAND2_X1 i_121 (.ZN (n_97), .A1 (p_0[1]), .A2 (Accumulator[1]));
AOI21_X1 i_120 (.ZN (n_96), .A (n_99), .B1 (n_98), .B2 (n_97));
OAI21_X1 i_119 (.ZN (n_95), .A (n_96), .B1 (p_0[2]), .B2 (Accumulator[2]));
NAND2_X1 i_118 (.ZN (n_94), .A1 (n_100), .A2 (n_95));
OAI22_X1 i_117 (.ZN (n_93), .A1 (p_0[3]), .A2 (Accumulator[3]), .B1 (n_101), .B2 (n_94));
NOR2_X1 i_116 (.ZN (n_92), .A1 (p_0[7]), .A2 (Accumulator[7]));
NOR2_X1 i_115 (.ZN (n_91), .A1 (p_0[5]), .A2 (Accumulator[5]));
NOR2_X1 i_114 (.ZN (n_90), .A1 (p_0[6]), .A2 (Accumulator[6]));
OR3_X1 i_113 (.ZN (n_89), .A1 (n_92), .A2 (n_90), .A3 (n_91));
NOR2_X1 i_112 (.ZN (n_88), .A1 (p_0[4]), .A2 (Accumulator[4]));
NOR3_X1 i_111 (.ZN (n_87), .A1 (n_89), .A2 (n_88), .A3 (n_93));
NAND2_X1 i_110 (.ZN (n_86), .A1 (p_0[4]), .A2 (Accumulator[4]));
NAND2_X1 i_109 (.ZN (n_85), .A1 (p_0[5]), .A2 (Accumulator[5]));
AOI21_X1 i_108 (.ZN (n_84), .A (n_89), .B1 (n_86), .B2 (n_85));
AND2_X1 i_107 (.ZN (n_83), .A1 (p_0[7]), .A2 (Accumulator[7]));
NAND2_X1 i_106 (.ZN (n_82), .A1 (p_0[6]), .A2 (Accumulator[6]));
INV_X1 i_105 (.ZN (n_81), .A (n_82));
NOR2_X1 i_104 (.ZN (n_80), .A1 (n_92), .A2 (n_82));
NOR4_X1 i_103 (.ZN (n_79), .A1 (n_83), .A2 (n_80), .A3 (n_84), .A4 (n_87));
NOR2_X1 i_102 (.ZN (n_78), .A1 (p_0[11]), .A2 (Accumulator[11]));
NOR2_X1 i_101 (.ZN (n_77), .A1 (p_0[9]), .A2 (Accumulator[9]));
NOR2_X1 i_100 (.ZN (n_76), .A1 (p_0[10]), .A2 (Accumulator[10]));
OR3_X1 i_99 (.ZN (n_75), .A1 (n_78), .A2 (n_76), .A3 (n_77));
NOR2_X1 i_98 (.ZN (n_74), .A1 (p_0[8]), .A2 (Accumulator[8]));
NOR3_X1 i_97 (.ZN (n_73), .A1 (n_75), .A2 (n_74), .A3 (n_79));
NAND2_X1 i_96 (.ZN (n_72), .A1 (p_0[8]), .A2 (Accumulator[8]));
NAND2_X1 i_95 (.ZN (n_71), .A1 (p_0[9]), .A2 (Accumulator[9]));
AOI21_X1 i_94 (.ZN (n_70), .A (n_75), .B1 (n_72), .B2 (n_71));
AND2_X1 i_93 (.ZN (n_69), .A1 (p_0[11]), .A2 (Accumulator[11]));
NAND2_X1 i_92 (.ZN (n_68), .A1 (p_0[10]), .A2 (Accumulator[10]));
INV_X1 i_91 (.ZN (n_67), .A (n_68));
NOR2_X1 i_90 (.ZN (n_66), .A1 (n_78), .A2 (n_68));
NOR4_X1 i_89 (.ZN (n_65), .A1 (n_69), .A2 (n_66), .A3 (n_70), .A4 (n_73));
NOR2_X1 i_88 (.ZN (n_64), .A1 (p_0[15]), .A2 (Accumulator[15]));
NOR2_X1 i_87 (.ZN (n_63), .A1 (p_0[13]), .A2 (Accumulator[13]));
NOR2_X1 i_86 (.ZN (n_62), .A1 (p_0[14]), .A2 (Accumulator[14]));
OR3_X1 i_85 (.ZN (n_61), .A1 (n_64), .A2 (n_62), .A3 (n_63));
NOR2_X1 i_84 (.ZN (n_60), .A1 (p_0[12]), .A2 (Accumulator[12]));
NOR3_X1 i_83 (.ZN (n_59), .A1 (n_61), .A2 (n_60), .A3 (n_65));
NAND2_X1 i_82 (.ZN (n_58), .A1 (p_0[12]), .A2 (Accumulator[12]));
NAND2_X1 i_81 (.ZN (n_57), .A1 (p_0[13]), .A2 (Accumulator[13]));
AOI21_X1 i_80 (.ZN (n_56), .A (n_61), .B1 (n_58), .B2 (n_57));
AND2_X1 i_79 (.ZN (n_55), .A1 (p_0[15]), .A2 (Accumulator[15]));
NAND2_X1 i_78 (.ZN (n_54), .A1 (p_0[14]), .A2 (Accumulator[14]));
INV_X1 i_77 (.ZN (n_53), .A (n_54));
NOR2_X1 i_76 (.ZN (n_52), .A1 (n_64), .A2 (n_54));
NOR4_X1 i_75 (.ZN (n_51), .A1 (n_55), .A2 (n_52), .A3 (n_56), .A4 (n_59));
INV_X1 i_74 (.ZN (n_50), .A (n_51));
NOR2_X1 i_73 (.ZN (n_49), .A1 (p_0[16]), .A2 (Accumulator[16]));
NOR2_X1 i_72 (.ZN (n_48), .A1 (n_106), .A2 (n_49));
AOI221_X1 i_71 (.ZN (n_47), .A (n_102), .B1 (p_0[19]), .B2 (Accumulator[19]), .C1 (n_50), .C2 (n_48));
OAI21_X1 i_70 (.ZN (n_46), .A (n_47), .B1 (n_115), .B2 (n_114));
INV_X1 i_69 (.ZN (n_45), .A (n_46));
NOR3_X1 i_68 (.ZN (n_44), .A1 (n_113), .A2 (n_110), .A3 (n_45));
NAND2_X1 i_67 (.ZN (n_43), .A1 (p_0[21]), .A2 (Accumulator[21]));
NOR2_X1 i_66 (.ZN (n_42), .A1 (n_113), .A2 (n_43));
AOI211_X1 i_65 (.ZN (n_41), .A (n_42), .B (n_44), .C1 (p_0[22]), .C2 (Accumulator[22]));
XNOR2_X1 i_64 (.ZN (Accumulator1[23]), .A (p_0[23]), .B (n_41));
AOI21_X1 i_63 (.ZN (n_40), .A (n_113), .B1 (p_0[22]), .B2 (Accumulator[22]));
OAI21_X1 i_62 (.ZN (n_39), .A (n_111), .B1 (n_115), .B2 (n_114));
OAI21_X1 i_61 (.ZN (n_38), .A (n_43), .B1 (n_110), .B2 (n_45));
XOR2_X1 i_60 (.Z (Accumulator1[22]), .A (n_40), .B (n_38));
OAI21_X1 i_59 (.ZN (n_37), .A (n_43), .B1 (p_0[21]), .B2 (Accumulator[21]));
NOR2_X1 i_58 (.ZN (n_36), .A1 (n_112), .A2 (n_45));
XNOR2_X1 i_57 (.ZN (Accumulator1[21]), .A (n_37), .B (n_36));
XOR2_X1 i_56 (.Z (Accumulator1[20]), .A (n_47), .B (n_39));
AOI21_X1 i_55 (.ZN (n_35), .A (n_109), .B1 (p_0[19]), .B2 (Accumulator[19]));
OAI21_X1 i_54 (.ZN (n_34), .A (n_105), .B1 (p_0[16]), .B2 (Accumulator[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_49), .B1 (n_105), .B2 (n_51));
AOI21_X1 i_52 (.ZN (n_32), .A (n_33), .B1 (p_0[17]), .B2 (Accumulator[17]));
AOI21_X1 i_51 (.ZN (n_31), .A (n_108), .B1 (p_0[17]), .B2 (Accumulator[17]));
OAI21_X1 i_50 (.ZN (n_30), .A (n_103), .B1 (n_107), .B2 (n_32));
XOR2_X1 i_49 (.Z (Accumulator1[19]), .A (n_35), .B (n_30));
OAI21_X1 i_48 (.ZN (n_29), .A (n_103), .B1 (p_0[18]), .B2 (Accumulator[18]));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_108), .A2 (n_32));
XNOR2_X1 i_46 (.ZN (Accumulator1[18]), .A (n_29), .B (n_28));
XOR2_X1 i_45 (.Z (Accumulator1[17]), .A (n_33), .B (n_31));
XOR2_X1 i_44 (.Z (Accumulator1[16]), .A (n_51), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_64), .A2 (n_55));
OAI21_X1 i_42 (.ZN (n_26), .A (n_58), .B1 (p_0[12]), .B2 (Accumulator[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_60), .B1 (n_65), .B2 (n_58));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_63), .B1 (n_57), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_63), .B1 (p_0[13]), .B2 (Accumulator[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (p_0[14]), .A2 (Accumulator[14]), .B1 (n_53), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (Accumulator1[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_62), .A2 (n_53));
XOR2_X1 i_34 (.Z (Accumulator1[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (Accumulator1[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (Accumulator1[12]), .A (n_65), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_78), .A2 (n_69));
AOI21_X1 i_30 (.ZN (n_18), .A (n_74), .B1 (p_0[8]), .B2 (Accumulator[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_74), .B1 (n_79), .B2 (n_72));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_77), .B1 (n_71), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_77), .B1 (p_0[9]), .B2 (Accumulator[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (p_0[10]), .A2 (Accumulator[10]), .B1 (n_67), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (Accumulator1[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_76), .A2 (n_67));
XOR2_X1 i_22 (.Z (Accumulator1[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (Accumulator1[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (Accumulator1[8]), .A (n_79), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_92), .A2 (n_83));
OAI21_X1 i_18 (.ZN (n_10), .A (n_86), .B1 (p_0[4]), .B2 (Accumulator[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_88), .B1 (n_93), .B2 (n_86));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_91), .B1 (n_85), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_91), .B1 (p_0[5]), .B2 (Accumulator[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (p_0[6]), .A2 (Accumulator[6]), .B1 (n_81), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (Accumulator1[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_90), .A2 (n_81));
XOR2_X1 i_10 (.Z (Accumulator1[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (Accumulator1[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (Accumulator1[4]), .A (n_93), .B (n_10));
XOR2_X1 i_7 (.Z (n_3), .A (p_0[3]), .B (Accumulator[3]));
XOR2_X1 i_6 (.Z (Accumulator1[3]), .A (n_94), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_100), .B1 (p_0[2]), .B2 (Accumulator[2]));
XNOR2_X1 i_4 (.ZN (Accumulator1[2]), .A (n_96), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_97), .B1 (p_0[1]), .B2 (Accumulator[1]));
XOR2_X1 i_2 (.Z (Accumulator1[1]), .A (n_98), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_98), .B1 (p_0[0]), .B2 (Accumulator[0]));
INV_X1 i_0 (.ZN (Accumulator1[0]), .A (n_0));

endmodule //datapath

module unsigned_seq_multiplier (clk, rst, start_s, a, b, c);

output [47:0] c;
input [23:0] a;
input [23:0] b;
input clk;
input rst;
input start_s;
wire \A_r[22] ;
wire \A_r[21] ;
wire \A_r[20] ;
wire \A_r[19] ;
wire \A_r[18] ;
wire \A_r[17] ;
wire \A_r[16] ;
wire \A_r[15] ;
wire \A_r[14] ;
wire \A_r[13] ;
wire \A_r[12] ;
wire \A_r[11] ;
wire \A_r[10] ;
wire \A_r[9] ;
wire \A_r[8] ;
wire \A_r[7] ;
wire \A_r[6] ;
wire \A_r[5] ;
wire \A_r[4] ;
wire \A_r[3] ;
wire \A_r[2] ;
wire \A_r[1] ;
wire \A_r[0] ;
wire n_1_0;
wire n_1_1;
wire n_1_2;
wire n_1_3;
wire n_1_4;
wire n_1_5;
wire n_1_6;
wire n_1_7;
wire n_1_8;
wire n_1_9;
wire n_1_10;
wire n_1_11;
wire n_1_12;
wire n_1_13;
wire n_1_14;
wire n_1_15;
wire n_1_16;
wire n_1_17;
wire n_1_18;
wire n_1_19;
wire n_1_20;
wire n_1_21;
wire n_1_22;
wire n_1_23;
wire n_1_24;
wire n_1_25;
wire n_1_26;
wire n_95;
wire n_24;
wire n_0;
wire n_94;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire uc_0;
wire n_118;
wire n_117;
wire n_116;
wire n_115;
wire n_114;
wire n_113;
wire n_112;
wire n_111;
wire n_110;
wire n_109;
wire n_108;
wire n_107;
wire n_106;
wire n_105;
wire n_104;
wire n_103;
wire n_102;
wire n_101;
wire n_100;
wire n_99;
wire n_98;
wire n_97;
wire n_96;
wire n_72;
wire n_120;
wire n_47;
wire n_1;
wire n_46;
wire n_2;
wire n_45;
wire n_3;
wire n_44;
wire n_4;
wire n_43;
wire n_5;
wire n_42;
wire n_6;
wire n_41;
wire n_7;
wire n_40;
wire n_8;
wire n_39;
wire n_9;
wire n_38;
wire n_10;
wire n_37;
wire n_11;
wire n_36;
wire n_12;
wire n_35;
wire n_13;
wire n_34;
wire n_14;
wire n_33;
wire n_15;
wire n_32;
wire n_16;
wire n_31;
wire n_17;
wire n_30;
wire n_18;
wire n_29;
wire n_19;
wire n_28;
wire n_20;
wire n_27;
wire n_21;
wire n_26;
wire n_22;
wire n_25;
wire n_23;
wire n_142;
wire n_141;
wire n_140;
wire n_139;
wire n_138;
wire n_137;
wire n_136;
wire n_135;
wire n_134;
wire n_133;
wire n_132;
wire n_131;
wire n_130;
wire n_129;
wire n_128;
wire n_127;
wire n_126;
wire n_125;
wire n_124;
wire n_123;
wire n_122;
wire n_121;
wire n_119;


INV_X1 i_1_119 (.ZN (n_1_26), .A (start_s));
MUX2_X1 i_1_118 (.Z (n_142), .A (\A_r[22] ), .B (a[22]), .S (start_s));
MUX2_X1 i_1_117 (.Z (n_141), .A (\A_r[21] ), .B (a[21]), .S (start_s));
MUX2_X1 i_1_116 (.Z (n_140), .A (\A_r[20] ), .B (a[20]), .S (start_s));
MUX2_X1 i_1_115 (.Z (n_139), .A (\A_r[19] ), .B (a[19]), .S (start_s));
MUX2_X1 i_1_114 (.Z (n_138), .A (\A_r[18] ), .B (a[18]), .S (start_s));
MUX2_X1 i_1_113 (.Z (n_137), .A (\A_r[17] ), .B (a[17]), .S (start_s));
MUX2_X1 i_1_112 (.Z (n_136), .A (\A_r[16] ), .B (a[16]), .S (start_s));
MUX2_X1 i_1_111 (.Z (n_135), .A (\A_r[15] ), .B (a[15]), .S (start_s));
MUX2_X1 i_1_110 (.Z (n_134), .A (\A_r[14] ), .B (a[14]), .S (start_s));
MUX2_X1 i_1_109 (.Z (n_133), .A (\A_r[13] ), .B (a[13]), .S (start_s));
MUX2_X1 i_1_108 (.Z (n_132), .A (\A_r[12] ), .B (a[12]), .S (start_s));
MUX2_X1 i_1_107 (.Z (n_131), .A (\A_r[11] ), .B (a[11]), .S (start_s));
MUX2_X1 i_1_106 (.Z (n_130), .A (\A_r[10] ), .B (a[10]), .S (start_s));
MUX2_X1 i_1_105 (.Z (n_129), .A (\A_r[9] ), .B (a[9]), .S (start_s));
MUX2_X1 i_1_104 (.Z (n_128), .A (\A_r[8] ), .B (a[8]), .S (start_s));
MUX2_X1 i_1_103 (.Z (n_127), .A (\A_r[7] ), .B (a[7]), .S (start_s));
MUX2_X1 i_1_102 (.Z (n_126), .A (\A_r[6] ), .B (a[6]), .S (start_s));
MUX2_X1 i_1_101 (.Z (n_125), .A (\A_r[5] ), .B (a[5]), .S (start_s));
MUX2_X1 i_1_100 (.Z (n_124), .A (\A_r[4] ), .B (a[4]), .S (start_s));
MUX2_X1 i_1_99 (.Z (n_123), .A (\A_r[3] ), .B (a[3]), .S (start_s));
MUX2_X1 i_1_98 (.Z (n_122), .A (\A_r[2] ), .B (a[2]), .S (start_s));
MUX2_X1 i_1_97 (.Z (n_121), .A (\A_r[1] ), .B (a[1]), .S (start_s));
MUX2_X1 i_1_96 (.Z (n_119), .A (\A_r[0] ), .B (a[0]), .S (start_s));
AND2_X1 i_1_95 (.ZN (n_118), .A1 (n_1_26), .A2 (n_0));
AND2_X1 i_1_94 (.ZN (n_117), .A1 (n_1_26), .A2 (c[45]));
AND2_X1 i_1_93 (.ZN (n_116), .A1 (n_1_26), .A2 (c[44]));
AND2_X1 i_1_92 (.ZN (n_115), .A1 (n_1_26), .A2 (c[43]));
AND2_X1 i_1_91 (.ZN (n_114), .A1 (n_1_26), .A2 (c[42]));
AND2_X1 i_1_90 (.ZN (n_113), .A1 (n_1_26), .A2 (c[41]));
AND2_X1 i_1_89 (.ZN (n_112), .A1 (n_1_26), .A2 (c[40]));
AND2_X1 i_1_88 (.ZN (n_111), .A1 (n_1_26), .A2 (c[39]));
AND2_X1 i_1_87 (.ZN (n_110), .A1 (n_1_26), .A2 (c[38]));
AND2_X1 i_1_86 (.ZN (n_109), .A1 (n_1_26), .A2 (c[37]));
AND2_X1 i_1_85 (.ZN (n_108), .A1 (n_1_26), .A2 (c[36]));
AND2_X1 i_1_84 (.ZN (n_107), .A1 (n_1_26), .A2 (c[35]));
AND2_X1 i_1_83 (.ZN (n_106), .A1 (n_1_26), .A2 (c[34]));
AND2_X1 i_1_82 (.ZN (n_105), .A1 (n_1_26), .A2 (c[33]));
AND2_X1 i_1_81 (.ZN (n_104), .A1 (n_1_26), .A2 (c[32]));
AND2_X1 i_1_80 (.ZN (n_103), .A1 (n_1_26), .A2 (c[31]));
AND2_X1 i_1_79 (.ZN (n_102), .A1 (n_1_26), .A2 (c[30]));
AND2_X1 i_1_78 (.ZN (n_101), .A1 (n_1_26), .A2 (c[29]));
AND2_X1 i_1_77 (.ZN (n_100), .A1 (n_1_26), .A2 (c[28]));
AND2_X1 i_1_76 (.ZN (n_99), .A1 (n_1_26), .A2 (c[27]));
AND2_X1 i_1_75 (.ZN (n_98), .A1 (n_1_26), .A2 (c[26]));
AND2_X1 i_1_74 (.ZN (n_97), .A1 (n_1_26), .A2 (c[25]));
AND2_X1 i_1_73 (.ZN (n_96), .A1 (n_1_26), .A2 (c[24]));
NOR2_X1 i_1_72 (.ZN (n_1_25), .A1 (n_1_0), .A2 (n_1_1));
INV_X1 i_1_71 (.ZN (n_71), .A (n_1_25));
INV_X1 i_1_70 (.ZN (n_70), .A (n_1_24));
AOI22_X1 i_1_69 (.ZN (n_1_24), .A1 (a[22]), .A2 (n_1_0), .B1 (\A_r[22] ), .B2 (n_1_1));
INV_X1 i_1_68 (.ZN (n_69), .A (n_1_23));
AOI22_X1 i_1_67 (.ZN (n_1_23), .A1 (a[21]), .A2 (n_1_0), .B1 (\A_r[21] ), .B2 (n_1_1));
INV_X1 i_1_66 (.ZN (n_68), .A (n_1_22));
AOI22_X1 i_1_65 (.ZN (n_1_22), .A1 (a[20]), .A2 (n_1_0), .B1 (\A_r[20] ), .B2 (n_1_1));
INV_X1 i_1_64 (.ZN (n_67), .A (n_1_21));
AOI22_X1 i_1_63 (.ZN (n_1_21), .A1 (a[19]), .A2 (n_1_0), .B1 (\A_r[19] ), .B2 (n_1_1));
INV_X1 i_1_62 (.ZN (n_66), .A (n_1_20));
AOI22_X1 i_1_61 (.ZN (n_1_20), .A1 (a[18]), .A2 (n_1_0), .B1 (\A_r[18] ), .B2 (n_1_1));
INV_X1 i_1_60 (.ZN (n_65), .A (n_1_19));
AOI22_X1 i_1_59 (.ZN (n_1_19), .A1 (a[17]), .A2 (n_1_0), .B1 (\A_r[17] ), .B2 (n_1_1));
INV_X1 i_1_58 (.ZN (n_64), .A (n_1_18));
AOI22_X1 i_1_57 (.ZN (n_1_18), .A1 (a[16]), .A2 (n_1_0), .B1 (\A_r[16] ), .B2 (n_1_1));
INV_X1 i_1_56 (.ZN (n_63), .A (n_1_17));
AOI22_X1 i_1_55 (.ZN (n_1_17), .A1 (a[15]), .A2 (n_1_0), .B1 (\A_r[15] ), .B2 (n_1_1));
INV_X1 i_1_54 (.ZN (n_62), .A (n_1_16));
AOI22_X1 i_1_53 (.ZN (n_1_16), .A1 (a[14]), .A2 (n_1_0), .B1 (\A_r[14] ), .B2 (n_1_1));
INV_X1 i_1_52 (.ZN (n_61), .A (n_1_15));
AOI22_X1 i_1_51 (.ZN (n_1_15), .A1 (a[13]), .A2 (n_1_0), .B1 (\A_r[13] ), .B2 (n_1_1));
INV_X1 i_1_50 (.ZN (n_60), .A (n_1_14));
AOI22_X1 i_1_49 (.ZN (n_1_14), .A1 (a[12]), .A2 (n_1_0), .B1 (\A_r[12] ), .B2 (n_1_1));
INV_X1 i_1_48 (.ZN (n_59), .A (n_1_13));
AOI22_X1 i_1_47 (.ZN (n_1_13), .A1 (a[11]), .A2 (n_1_0), .B1 (\A_r[11] ), .B2 (n_1_1));
INV_X1 i_1_46 (.ZN (n_58), .A (n_1_12));
AOI22_X1 i_1_45 (.ZN (n_1_12), .A1 (a[10]), .A2 (n_1_0), .B1 (\A_r[10] ), .B2 (n_1_1));
INV_X1 i_1_44 (.ZN (n_57), .A (n_1_11));
AOI22_X1 i_1_43 (.ZN (n_1_11), .A1 (a[9]), .A2 (n_1_0), .B1 (\A_r[9] ), .B2 (n_1_1));
INV_X1 i_1_42 (.ZN (n_56), .A (n_1_10));
AOI22_X1 i_1_41 (.ZN (n_1_10), .A1 (a[8]), .A2 (n_1_0), .B1 (\A_r[8] ), .B2 (n_1_1));
INV_X1 i_1_40 (.ZN (n_55), .A (n_1_9));
AOI22_X1 i_1_39 (.ZN (n_1_9), .A1 (a[7]), .A2 (n_1_0), .B1 (\A_r[7] ), .B2 (n_1_1));
INV_X1 i_1_38 (.ZN (n_54), .A (n_1_8));
AOI22_X1 i_1_37 (.ZN (n_1_8), .A1 (a[6]), .A2 (n_1_0), .B1 (\A_r[6] ), .B2 (n_1_1));
INV_X1 i_1_36 (.ZN (n_53), .A (n_1_7));
AOI22_X1 i_1_35 (.ZN (n_1_7), .A1 (a[5]), .A2 (n_1_0), .B1 (\A_r[5] ), .B2 (n_1_1));
INV_X1 i_1_34 (.ZN (n_52), .A (n_1_6));
AOI22_X1 i_1_33 (.ZN (n_1_6), .A1 (a[4]), .A2 (n_1_0), .B1 (\A_r[4] ), .B2 (n_1_1));
INV_X1 i_1_32 (.ZN (n_51), .A (n_1_5));
AOI22_X1 i_1_31 (.ZN (n_1_5), .A1 (a[3]), .A2 (n_1_0), .B1 (\A_r[3] ), .B2 (n_1_1));
INV_X1 i_1_30 (.ZN (n_50), .A (n_1_4));
AOI22_X1 i_1_29 (.ZN (n_1_4), .A1 (a[2]), .A2 (n_1_0), .B1 (\A_r[2] ), .B2 (n_1_1));
INV_X1 i_1_28 (.ZN (n_49), .A (n_1_3));
AOI22_X1 i_1_27 (.ZN (n_1_3), .A1 (a[1]), .A2 (n_1_0), .B1 (\A_r[1] ), .B2 (n_1_1));
INV_X1 i_1_26 (.ZN (n_48), .A (n_1_2));
AOI22_X1 i_1_25 (.ZN (n_1_2), .A1 (a[0]), .A2 (n_1_0), .B1 (\A_r[0] ), .B2 (n_1_1));
AND2_X1 i_1_24 (.ZN (n_1_1), .A1 (n_1_26), .A2 (n_23));
AND2_X1 i_1_23 (.ZN (n_1_0), .A1 (start_s), .A2 (b[0]));
OR2_X1 i_1_22 (.ZN (n_47), .A1 (start_s), .A2 (c[23]));
MUX2_X1 i_1_21 (.Z (n_46), .A (n_1), .B (b[22]), .S (start_s));
MUX2_X1 i_1_20 (.Z (n_45), .A (n_2), .B (b[21]), .S (start_s));
MUX2_X1 i_1_19 (.Z (n_44), .A (n_3), .B (b[20]), .S (start_s));
MUX2_X1 i_1_18 (.Z (n_43), .A (n_4), .B (b[19]), .S (start_s));
MUX2_X1 i_1_17 (.Z (n_42), .A (n_5), .B (b[18]), .S (start_s));
MUX2_X1 i_1_16 (.Z (n_41), .A (n_6), .B (b[17]), .S (start_s));
MUX2_X1 i_1_15 (.Z (n_40), .A (n_7), .B (b[16]), .S (start_s));
MUX2_X1 i_1_14 (.Z (n_39), .A (n_8), .B (b[15]), .S (start_s));
MUX2_X1 i_1_13 (.Z (n_38), .A (n_9), .B (b[14]), .S (start_s));
MUX2_X1 i_1_12 (.Z (n_37), .A (n_10), .B (b[13]), .S (start_s));
MUX2_X1 i_1_11 (.Z (n_36), .A (n_11), .B (b[12]), .S (start_s));
MUX2_X1 i_1_10 (.Z (n_35), .A (n_12), .B (b[11]), .S (start_s));
MUX2_X1 i_1_9 (.Z (n_34), .A (n_13), .B (b[10]), .S (start_s));
MUX2_X1 i_1_8 (.Z (n_33), .A (n_14), .B (b[9]), .S (start_s));
MUX2_X1 i_1_7 (.Z (n_32), .A (n_15), .B (b[8]), .S (start_s));
MUX2_X1 i_1_6 (.Z (n_31), .A (n_16), .B (b[7]), .S (start_s));
MUX2_X1 i_1_5 (.Z (n_30), .A (n_17), .B (b[6]), .S (start_s));
MUX2_X1 i_1_4 (.Z (n_29), .A (n_18), .B (b[5]), .S (start_s));
MUX2_X1 i_1_3 (.Z (n_28), .A (n_19), .B (b[4]), .S (start_s));
MUX2_X1 i_1_2 (.Z (n_27), .A (n_20), .B (b[3]), .S (start_s));
MUX2_X1 i_1_1 (.Z (n_26), .A (n_21), .B (b[2]), .S (start_s));
MUX2_X1 i_1_0 (.Z (n_25), .A (n_22), .B (b[1]), .S (start_s));
CLKGATETST_X1 clk_gate_B_r_reg (.GCK (n_120), .CK (clk), .E (n_24), .SE (1'b0 ));
INV_X4 i_0_0 (.ZN (n_24), .A (rst));
DFF_X1 \A_r_reg[0]  (.Q (\A_r[0] ), .CK (n_120), .D (n_119));
DFF_X1 \A_r_reg[1]  (.Q (\A_r[1] ), .CK (n_120), .D (n_121));
DFF_X1 \A_r_reg[2]  (.Q (\A_r[2] ), .CK (n_120), .D (n_122));
DFF_X1 \A_r_reg[3]  (.Q (\A_r[3] ), .CK (n_120), .D (n_123));
DFF_X1 \A_r_reg[4]  (.Q (\A_r[4] ), .CK (n_120), .D (n_124));
DFF_X1 \A_r_reg[5]  (.Q (\A_r[5] ), .CK (n_120), .D (n_125));
DFF_X1 \A_r_reg[6]  (.Q (\A_r[6] ), .CK (n_120), .D (n_126));
DFF_X1 \A_r_reg[7]  (.Q (\A_r[7] ), .CK (n_120), .D (n_127));
DFF_X1 \A_r_reg[8]  (.Q (\A_r[8] ), .CK (n_120), .D (n_128));
DFF_X1 \A_r_reg[9]  (.Q (\A_r[9] ), .CK (n_120), .D (n_129));
DFF_X1 \A_r_reg[10]  (.Q (\A_r[10] ), .CK (n_120), .D (n_130));
DFF_X1 \A_r_reg[11]  (.Q (\A_r[11] ), .CK (n_120), .D (n_131));
DFF_X1 \A_r_reg[12]  (.Q (\A_r[12] ), .CK (n_120), .D (n_132));
DFF_X1 \A_r_reg[13]  (.Q (\A_r[13] ), .CK (n_120), .D (n_133));
DFF_X1 \A_r_reg[14]  (.Q (\A_r[14] ), .CK (n_120), .D (n_134));
DFF_X1 \A_r_reg[15]  (.Q (\A_r[15] ), .CK (n_120), .D (n_135));
DFF_X1 \A_r_reg[16]  (.Q (\A_r[16] ), .CK (n_120), .D (n_136));
DFF_X1 \A_r_reg[17]  (.Q (\A_r[17] ), .CK (n_120), .D (n_137));
DFF_X1 \A_r_reg[18]  (.Q (\A_r[18] ), .CK (n_120), .D (n_138));
DFF_X1 \A_r_reg[19]  (.Q (\A_r[19] ), .CK (n_120), .D (n_139));
DFF_X1 \A_r_reg[20]  (.Q (\A_r[20] ), .CK (n_120), .D (n_140));
DFF_X1 \A_r_reg[21]  (.Q (\A_r[21] ), .CK (n_120), .D (n_141));
DFF_X1 \A_r_reg[22]  (.Q (\A_r[22] ), .CK (n_120), .D (n_142));
DFF_X1 \B_r_reg[0]  (.Q (n_23), .CK (n_120), .D (n_25));
DFF_X1 \B_r_reg[1]  (.Q (n_22), .CK (n_120), .D (n_26));
DFF_X1 \B_r_reg[2]  (.Q (n_21), .CK (n_120), .D (n_27));
DFF_X1 \B_r_reg[3]  (.Q (n_20), .CK (n_120), .D (n_28));
DFF_X1 \B_r_reg[4]  (.Q (n_19), .CK (n_120), .D (n_29));
DFF_X1 \B_r_reg[5]  (.Q (n_18), .CK (n_120), .D (n_30));
DFF_X1 \B_r_reg[6]  (.Q (n_17), .CK (n_120), .D (n_31));
DFF_X1 \B_r_reg[7]  (.Q (n_16), .CK (n_120), .D (n_32));
DFF_X1 \B_r_reg[8]  (.Q (n_15), .CK (n_120), .D (n_33));
DFF_X1 \B_r_reg[9]  (.Q (n_14), .CK (n_120), .D (n_34));
DFF_X1 \B_r_reg[10]  (.Q (n_13), .CK (n_120), .D (n_35));
DFF_X1 \B_r_reg[11]  (.Q (n_12), .CK (n_120), .D (n_36));
DFF_X1 \B_r_reg[12]  (.Q (n_11), .CK (n_120), .D (n_37));
DFF_X1 \B_r_reg[13]  (.Q (n_10), .CK (n_120), .D (n_38));
DFF_X1 \B_r_reg[14]  (.Q (n_9), .CK (n_120), .D (n_39));
DFF_X1 \B_r_reg[15]  (.Q (n_8), .CK (n_120), .D (n_40));
DFF_X1 \B_r_reg[16]  (.Q (n_7), .CK (n_120), .D (n_41));
DFF_X1 \B_r_reg[17]  (.Q (n_6), .CK (n_120), .D (n_42));
DFF_X1 \B_r_reg[18]  (.Q (n_5), .CK (n_120), .D (n_43));
DFF_X1 \B_r_reg[19]  (.Q (n_4), .CK (n_120), .D (n_44));
DFF_X1 \B_r_reg[20]  (.Q (n_3), .CK (n_120), .D (n_45));
DFF_X1 \B_r_reg[21]  (.Q (n_2), .CK (n_120), .D (n_46));
DFF_X1 \B_r_reg[22]  (.Q (n_1), .CK (n_120), .D (n_47));
DFF_X1 \B_r_reg[23]  (.Q (c[23]), .CK (n_120), .D (n_72));
datapath i_4 (.Accumulator1 ({n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, 
    n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72}), .Accumulator ({uc_0, n_118, n_117, n_116, n_115, n_114, n_113, 
    n_112, n_111, n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, 
    n_101, n_100, n_99, n_98, n_97, n_96}), .p_0 ({n_71, n_70, n_69, n_68, n_67, 
    n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
    n_53, n_52, n_51, n_50, n_49, n_48}));
DFFR_X1 \Accumulator_reg[0]  (.Q (c[24]), .CK (clk), .D (n_73), .RN (n_24));
DFFR_X1 \Accumulator_reg[1]  (.Q (c[25]), .CK (clk), .D (n_74), .RN (n_24));
DFFR_X1 \Accumulator_reg[2]  (.Q (c[26]), .CK (clk), .D (n_75), .RN (n_24));
DFFR_X1 \Accumulator_reg[3]  (.Q (c[27]), .CK (clk), .D (n_76), .RN (n_24));
DFFR_X1 \Accumulator_reg[4]  (.Q (c[28]), .CK (clk), .D (n_77), .RN (n_24));
DFFR_X1 \Accumulator_reg[5]  (.Q (c[29]), .CK (clk), .D (n_78), .RN (n_24));
DFFR_X1 \Accumulator_reg[6]  (.Q (c[30]), .CK (clk), .D (n_79), .RN (n_24));
DFFR_X1 \Accumulator_reg[7]  (.Q (c[31]), .CK (clk), .D (n_80), .RN (n_24));
DFFR_X1 \Accumulator_reg[8]  (.Q (c[32]), .CK (clk), .D (n_81), .RN (n_24));
DFFR_X1 \Accumulator_reg[9]  (.Q (c[33]), .CK (clk), .D (n_82), .RN (n_24));
DFFR_X1 \Accumulator_reg[10]  (.Q (c[34]), .CK (clk), .D (n_83), .RN (n_24));
DFFR_X1 \Accumulator_reg[11]  (.Q (c[35]), .CK (clk), .D (n_84), .RN (n_24));
DFFR_X1 \Accumulator_reg[12]  (.Q (c[36]), .CK (clk), .D (n_85), .RN (n_24));
DFFR_X1 \Accumulator_reg[13]  (.Q (c[37]), .CK (clk), .D (n_86), .RN (n_24));
DFFR_X1 \Accumulator_reg[14]  (.Q (c[38]), .CK (clk), .D (n_87), .RN (n_24));
DFFR_X1 \Accumulator_reg[15]  (.Q (c[39]), .CK (clk), .D (n_88), .RN (n_24));
DFFR_X1 \Accumulator_reg[16]  (.Q (c[40]), .CK (clk), .D (n_89), .RN (n_24));
DFFR_X1 \Accumulator_reg[17]  (.Q (c[41]), .CK (clk), .D (n_90), .RN (n_24));
DFFR_X1 \Accumulator_reg[18]  (.Q (c[42]), .CK (clk), .D (n_91), .RN (n_24));
DFFR_X1 \Accumulator_reg[19]  (.Q (c[43]), .CK (clk), .D (n_92), .RN (n_24));
DFFR_X1 \Accumulator_reg[20]  (.Q (c[44]), .CK (clk), .D (n_93), .RN (n_24));
DFFR_X1 \Accumulator_reg[21]  (.Q (c[45]), .CK (clk), .D (n_94), .RN (n_24));
DFFR_X1 \Accumulator_reg[22]  (.Q (n_0), .CK (clk), .D (n_95), .RN (n_24));

endmodule //unsigned_seq_multiplier

module fp_mul (clk, rst, a_s, b_s, c_out, overflow);

output [31:0] c_out;
output overflow;
input [31:0] a_s;
input [31:0] b_s;
input clk;
input rst;
wire sph_n82;
wire sph_n232;
wire sph_n217;
wire sph_n102;
wire sph_n227;
wire sph_n157;
wire sph_n242;
wire sph_n147;
wire sph_n77;
wire sph_n292;
wire sph_n262;
wire sph_n187;
wire sph_n162;
wire sph_n152;
wire sph_n92;
wire sph_n12;
wire sph_n37;
wire sph_n307;
wire sph_n302;
wire sph_n312;
wire sph_n22;
wire sph_n112;
wire sph_n252;
wire sph_n267;
wire sph_n277;
wire sph_n297;
wire sph_n222;
wire sph_n237;
wire sph_n282;
wire sph_n127;
wire sph_n47;
wire sph_n32;
wire sph_n322;
wire sph_n87;
wire sph_n17;
wire sph_n62;
wire sph_n122;
wire sph_n57;
wire sph_n287;
wire sph_n107;
wire sph_n27;
wire sph_n317;
wire sph_n42;
wire sph_n72;
wire sph_n67;
wire sph_n132;
wire sph_n257;
wire sph_n212;
wire sph_n142;
wire sph_n117;
wire sph_n7;
wire sph_n52;
wire sph_n172;
wire sph_n197;
wire sph_n207;
wire sph_n177;
wire sph_n247;
wire sph_n137;
wire sph_n97;
wire sph_n202;
wire sph_n272;
wire sph_n192;
wire sph_n167;
wire sph_n182;
wire sps__n1;
wire \res_mant[23] ;
wire \res_mant[22] ;
wire \res_mant[21] ;
wire \res_mant[20] ;
wire \res_mant[19] ;
wire \res_mant[18] ;
wire \res_mant[17] ;
wire \res_mant[16] ;
wire \res_mant[15] ;
wire \res_mant[14] ;
wire \res_mant[13] ;
wire \res_mant[12] ;
wire \res_mant[11] ;
wire \res_mant[10] ;
wire \res_mant[9] ;
wire \res_mant[8] ;
wire \res_mant[7] ;
wire \res_mant[6] ;
wire \res_mant[5] ;
wire \res_mant[4] ;
wire \res_mant[3] ;
wire \res_mant[2] ;
wire \res_mant[1] ;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire mul_start;
wire n_0_41;
wire b;
wire a;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire \counter[4] ;
wire \counter[3] ;
wire \counter[2] ;
wire \counter[1] ;
wire \counter[0] ;
wire n_0_50;
wire n_0_40;
wire n_0_0_12;
wire n_0_0_2;
wire n_0_0_13;
wire n_0_0_3;
wire n_0_0_14;
wire n_0_0_4;
wire n_0_0_15;
wire n_0_0_5;
wire n_0_0_16;
wire n_0_0_6;
wire n_0_0_17;
wire n_0_0_7;
wire n_0_0_18;
wire n_0_0_8;
wire n_0_0_19;
wire n_0_0_0;
wire n_0_0_20;
wire n_0_0_1;
wire n_0_0_21;
wire n_0_0_9;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_0_22;
wire n_0_0_10;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_0_23;
wire n_0_90;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_98;
wire n_0_0_34;
wire start;
wire n_0_97;
wire n_0_0_11;
wire n_0_96;
wire n_0_0_33;
wire n_0_0_35;
wire n_0_99;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_0_38;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;


INV_X1 i_0_0_70 (.ZN (n_0_0_38), .A (rst));
OR2_X1 i_0_0_69 (.ZN (n_0_0_37), .A1 (\counter[2] ), .A2 (\counter[1] ));
NAND3_X1 i_0_0_68 (.ZN (n_0_0_36), .A1 (\counter[4] ), .A2 (\counter[3] ), .A3 (\counter[0] ));
OAI21_X1 i_0_0_67 (.ZN (n_0_99), .A (n_0_0_38), .B1 (n_0_0_37), .B2 (n_0_0_36));
INV_X1 i_0_0_66 (.ZN (n_0_0_35), .A (n_0_99));
NOR2_X1 i_0_0_65 (.ZN (n_0_0_33), .A1 (\counter[4] ), .A2 (n_0_0_9));
AOI211_X1 i_0_0_64 (.ZN (n_0_96), .A (n_0_0_33), .B (n_0_99), .C1 (\counter[4] ), .C2 (n_0_0_9));
INV_X1 i_0_0_63 (.ZN (n_0_0_11), .A (n_0_42));
INV_X1 i_0_0_62 (.ZN (n_0_97), .A (rst));
NOR4_X1 i_0_0_61 (.ZN (start), .A1 (n_0_0_37), .A2 (\counter[0] ), .A3 (\counter[3] ), .A4 (\counter[4] ));
OAI21_X1 i_0_0_60 (.ZN (n_0_0_34), .A (n_0_97), .B1 (n_0_0_11), .B2 (n_0_0_8));
AOI21_X1 i_0_0_59 (.ZN (n_0_98), .A (n_0_0_34), .B1 (n_0_0_8), .B2 (n_0_0_11));
AND2_X1 i_0_0_58 (.ZN (n_0_95), .A1 (n_0_0_21), .A2 (n_0_0_35));
AND2_X1 i_0_0_57 (.ZN (n_0_94), .A1 (n_0_0_20), .A2 (n_0_0_35));
AND2_X1 i_0_0_56 (.ZN (n_0_93), .A1 (n_0_0_19), .A2 (n_0_0_35));
NOR2_X1 i_0_0_55 (.ZN (n_0_92), .A1 (rst), .A2 (\counter[0] ));
AND2_X1 i_0_0_54 (.ZN (n_0_91), .A1 (start), .A2 (n_0_97));
NOR4_X1 i_0_0_53 (.ZN (n_0_0_32), .A1 (n_0_55), .A2 (n_0_56), .A3 (n_0_57), .A4 (n_0_58));
NOR4_X1 i_0_0_52 (.ZN (n_0_0_31), .A1 (n_0_51), .A2 (n_0_52), .A3 (n_0_53), .A4 (n_0_54));
NAND2_X1 i_0_0_51 (.ZN (n_0_0_30), .A1 (n_0_0_32), .A2 (n_0_0_31));
NOR4_X1 i_0_0_50 (.ZN (n_0_0_29), .A1 (n_0_46), .A2 (n_0_47), .A3 (n_0_48), .A4 (n_0_49));
NOR4_X1 i_0_0_49 (.ZN (n_0_0_28), .A1 (n_0_42), .A2 (n_0_43), .A3 (n_0_44), .A4 (n_0_45));
NAND2_X1 i_0_0_48 (.ZN (n_0_0_27), .A1 (n_0_0_29), .A2 (n_0_0_28));
NAND2_X1 i_0_0_47 (.ZN (n_0_0_26), .A1 (n_0_0_30), .A2 (n_0_0_27));
NAND3_X1 i_0_0_46 (.ZN (n_0_0_25), .A1 (n_0_0_30), .A2 (n_0_0_27), .A3 (b));
XNOR2_X1 i_0_0_45 (.ZN (n_0_0_24), .A (a), .B (n_0_0_25));
AND2_X1 i_0_0_44 (.ZN (n_0_90), .A1 (n_0_0_24), .A2 (n_0_97));
NOR2_X2 i_0_0_43 (.ZN (n_0_0_23), .A1 (n_0_0_26), .A2 (rst));
AND2_X1 i_0_0_42 (.ZN (n_0_89), .A1 (n_0_0_18), .A2 (n_0_0_23));
AND2_X1 i_0_0_41 (.ZN (n_0_88), .A1 (n_0_0_17), .A2 (n_0_0_23));
AND2_X1 i_0_0_40 (.ZN (n_0_87), .A1 (n_0_0_16), .A2 (n_0_0_23));
AND2_X1 i_0_0_39 (.ZN (n_0_86), .A1 (n_0_0_15), .A2 (n_0_0_23));
AND2_X1 i_0_0_38 (.ZN (n_0_85), .A1 (n_0_0_14), .A2 (n_0_0_23));
AND2_X1 i_0_0_37 (.ZN (n_0_84), .A1 (n_0_0_13), .A2 (n_0_0_23));
AND2_X1 i_0_0_36 (.ZN (n_0_83), .A1 (n_0_0_12), .A2 (n_0_0_23));
OR2_X1 i_0_0_35 (.ZN (n_0_0_10), .A1 (n_0_49), .A2 (n_0_58));
NAND2_X1 i_0_0_34 (.ZN (n_0_0_22), .A1 (n_0_49), .A2 (n_0_58));
AOI211_X1 i_0_0_33 (.ZN (n_0_82), .A (rst), .B (n_0_0_26), .C1 (n_0_0_10), .C2 (n_0_0_22));
AND2_X1 i_0_0_32 (.ZN (n_0_81), .A1 (\res_mant[23] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_31 (.ZN (n_0_80), .A1 (\res_mant[22] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_30 (.ZN (n_0_79), .A1 (\res_mant[21] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_29 (.ZN (n_0_78), .A1 (\res_mant[20] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_28 (.ZN (n_0_77), .A1 (\res_mant[19] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_27 (.ZN (n_0_76), .A1 (\res_mant[18] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_26 (.ZN (n_0_75), .A1 (\res_mant[17] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_25 (.ZN (n_0_74), .A1 (\res_mant[16] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_24 (.ZN (n_0_73), .A1 (\res_mant[15] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_23 (.ZN (n_0_72), .A1 (\res_mant[14] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_22 (.ZN (n_0_71), .A1 (\res_mant[13] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_21 (.ZN (n_0_70), .A1 (\res_mant[12] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_20 (.ZN (n_0_69), .A1 (\res_mant[11] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_19 (.ZN (n_0_68), .A1 (\res_mant[10] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_18 (.ZN (n_0_67), .A1 (\res_mant[9] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_17 (.ZN (n_0_66), .A1 (\res_mant[8] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_16 (.ZN (n_0_65), .A1 (\res_mant[7] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_15 (.ZN (n_0_64), .A1 (\res_mant[6] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_14 (.ZN (n_0_63), .A1 (\res_mant[5] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_13 (.ZN (n_0_62), .A1 (\res_mant[4] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_12 (.ZN (n_0_61), .A1 (\res_mant[3] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_11 (.ZN (n_0_60), .A1 (\res_mant[2] ), .A2 (n_0_0_23));
AND2_X1 i_0_0_10 (.ZN (n_0_59), .A1 (\res_mant[1] ), .A2 (n_0_0_23));
HA_X1 i_0_0_9 (.CO (n_0_0_9), .S (n_0_0_21), .A (\counter[3] ), .B (n_0_0_1));
HA_X1 i_0_0_8 (.CO (n_0_0_1), .S (n_0_0_20), .A (\counter[2] ), .B (n_0_0_0));
HA_X1 i_0_0_7 (.CO (n_0_0_0), .S (n_0_0_19), .A (\counter[1] ), .B (\counter[0] ));
FA_X1 i_0_0_6 (.CO (n_0_0_8), .S (n_0_0_18), .A (n_0_51), .B (n_0_0_11), .CI (n_0_0_7));
FA_X1 i_0_0_5 (.CO (n_0_0_7), .S (n_0_0_17), .A (n_0_43), .B (n_0_52), .CI (n_0_0_6));
FA_X1 i_0_0_4 (.CO (n_0_0_6), .S (n_0_0_16), .A (n_0_44), .B (n_0_53), .CI (n_0_0_5));
FA_X1 i_0_0_3 (.CO (n_0_0_5), .S (n_0_0_15), .A (n_0_45), .B (n_0_54), .CI (n_0_0_4));
FA_X1 i_0_0_2 (.CO (n_0_0_4), .S (n_0_0_14), .A (n_0_46), .B (n_0_55), .CI (n_0_0_3));
FA_X1 i_0_0_1 (.CO (n_0_0_3), .S (n_0_0_13), .A (n_0_47), .B (n_0_56), .CI (n_0_0_2));
FA_X1 i_0_0_0 (.CO (n_0_0_2), .S (n_0_0_12), .A (n_0_48), .B (n_0_57), .CI (n_0_0_10));
CLKGATETST_X1 clk_gate_b_reg__1 (.GCK (n_0_40), .CK (clk), .E (n_0_91), .SE (1'b0 ));
CLKGATETST_X1 clk_gate_overflow_reg (.GCK (n_0_50), .CK (clk), .E (n_0_99), .SE (1'b0 ));
DFF_X1 \counter_reg[0]  (.Q (\counter[0] ), .CK (clk), .D (n_0_92));
DFF_X1 \counter_reg[1]  (.Q (\counter[1] ), .CK (clk), .D (n_0_93));
DFF_X1 \counter_reg[2]  (.Q (\counter[2] ), .CK (clk), .D (n_0_94));
DFF_X1 \counter_reg[3]  (.Q (\counter[3] ), .CK (clk), .D (n_0_95));
DFF_X1 \counter_reg[4]  (.Q (\counter[4] ), .CK (clk), .D (n_0_96));
DFF_X1 \a_reg[23]  (.Q (n_0_58), .CK (n_0_40), .D (sph_n77));
DFF_X1 \a_reg[24]  (.Q (n_0_57), .CK (n_0_40), .D (sph_n147));
DFF_X1 \a_reg[25]  (.Q (n_0_56), .CK (n_0_40), .D (sph_n242));
DFF_X1 \a_reg[26]  (.Q (n_0_55), .CK (n_0_40), .D (sph_n157));
DFF_X1 \a_reg[27]  (.Q (n_0_54), .CK (n_0_40), .D (sph_n227));
DFF_X1 \a_reg[28]  (.Q (n_0_53), .CK (n_0_40), .D (sph_n102));
DFF_X1 \a_reg[29]  (.Q (n_0_52), .CK (n_0_40), .D (sph_n217));
DFF_X1 \a_reg[30]  (.Q (n_0_51), .CK (n_0_40), .D (sph_n232));
DFF_X1 \b_reg[23]  (.Q (n_0_49), .CK (n_0_40), .D (sph_n27));
DFF_X1 \b_reg[24]  (.Q (n_0_48), .CK (n_0_40), .D (sph_n107));
DFF_X1 \b_reg[25]  (.Q (n_0_47), .CK (n_0_40), .D (sph_n287));
DFF_X1 \b_reg[26]  (.Q (n_0_46), .CK (n_0_40), .D (sph_n57));
DFF_X1 \b_reg[27]  (.Q (n_0_45), .CK (n_0_40), .D (sph_n122));
DFF_X1 \b_reg[28]  (.Q (n_0_44), .CK (n_0_40), .D (sph_n62));
DFF_X1 \b_reg[29]  (.Q (n_0_43), .CK (n_0_40), .D (sph_n17));
DFF_X1 \b_reg[30]  (.Q (n_0_42), .CK (n_0_40), .D (sph_n87));
DFF_X1 \a_reg[31]  (.Q (a), .CK (n_0_40), .D (sph_n82));
DFF_X1 \b_reg[31]  (.Q (b), .CK (n_0_40), .D (sph_n322));
MUX2_X1 mul_start_reg_enable_mux_0 (.Z (n_0_41), .A (mul_start), .B (start), .S (n_0_97));
DFF_X1 mul_start_reg (.Q (sps__n1), .CK (clk), .D (n_0_41));
DFF_X1 \a_reg[0]  (.Q (n_0_39), .CK (n_0_40), .D (sph_n32));
DFF_X1 \a_reg[1]  (.Q (n_0_38), .CK (n_0_40), .D (sph_n47));
DFF_X1 \a_reg[2]  (.Q (n_0_37), .CK (n_0_40), .D (sph_n127));
DFF_X1 \a_reg[3]  (.Q (n_0_36), .CK (n_0_40), .D (sph_n282));
DFF_X1 \a_reg[4]  (.Q (n_0_35), .CK (n_0_40), .D (sph_n237));
DFF_X1 \a_reg[5]  (.Q (n_0_34), .CK (n_0_40), .D (sph_n222));
DFF_X1 \a_reg[6]  (.Q (n_0_33), .CK (n_0_40), .D (sph_n297));
DFF_X1 \a_reg[7]  (.Q (n_0_32), .CK (n_0_40), .D (sph_n277));
DFF_X1 \a_reg[8]  (.Q (n_0_31), .CK (n_0_40), .D (sph_n267));
DFF_X1 \a_reg[9]  (.Q (n_0_30), .CK (n_0_40), .D (sph_n252));
DFF_X1 \a_reg[10]  (.Q (n_0_29), .CK (n_0_40), .D (sph_n112));
DFF_X1 \a_reg[11]  (.Q (n_0_28), .CK (n_0_40), .D (sph_n22));
DFF_X1 \a_reg[12]  (.Q (n_0_27), .CK (n_0_40), .D (sph_n312));
DFF_X1 \a_reg[13]  (.Q (n_0_26), .CK (n_0_40), .D (sph_n302));
DFF_X1 \a_reg[14]  (.Q (n_0_25), .CK (n_0_40), .D (sph_n307));
DFF_X1 \a_reg[15]  (.Q (n_0_24), .CK (n_0_40), .D (sph_n37));
DFF_X1 \a_reg[16]  (.Q (n_0_23), .CK (n_0_40), .D (sph_n12));
DFF_X1 \a_reg[17]  (.Q (n_0_22), .CK (n_0_40), .D (sph_n92));
DFF_X1 \a_reg[18]  (.Q (n_0_21), .CK (n_0_40), .D (sph_n152));
DFF_X1 \a_reg[19]  (.Q (n_0_20), .CK (n_0_40), .D (sph_n162));
DFF_X1 \a_reg[20]  (.Q (n_0_19), .CK (n_0_40), .D (sph_n187));
DFF_X1 \a_reg[21]  (.Q (n_0_18), .CK (n_0_40), .D (sph_n262));
DFF_X1 \a_reg[22]  (.Q (n_0_17), .CK (n_0_40), .D (sph_n292));
DFF_X1 \b_reg[0]  (.Q (n_0_16), .CK (n_0_40), .D (sph_n182));
DFF_X1 \b_reg[1]  (.Q (n_0_15), .CK (n_0_40), .D (sph_n167));
DFF_X1 \b_reg[2]  (.Q (n_0_14), .CK (n_0_40), .D (sph_n192));
DFF_X1 \b_reg[3]  (.Q (n_0_13), .CK (n_0_40), .D (sph_n272));
DFF_X1 \b_reg[4]  (.Q (n_0_12), .CK (n_0_40), .D (sph_n202));
DFF_X1 \b_reg[5]  (.Q (n_0_11), .CK (n_0_40), .D (sph_n97));
DFF_X1 \b_reg[6]  (.Q (n_0_10), .CK (n_0_40), .D (sph_n137));
DFF_X1 \b_reg[7]  (.Q (n_0_9), .CK (n_0_40), .D (sph_n247));
DFF_X1 \b_reg[8]  (.Q (n_0_8), .CK (n_0_40), .D (sph_n177));
DFF_X1 \b_reg[9]  (.Q (n_0_7), .CK (n_0_40), .D (sph_n207));
DFF_X1 \b_reg[10]  (.Q (n_0_6), .CK (n_0_40), .D (sph_n197));
DFF_X1 \b_reg[11]  (.Q (n_0_5), .CK (n_0_40), .D (sph_n172));
DFF_X1 \b_reg[12]  (.Q (n_0_4), .CK (n_0_40), .D (sph_n52));
DFF_X1 \b_reg[13]  (.Q (n_0_3), .CK (n_0_40), .D (sph_n7));
DFF_X1 \b_reg[14]  (.Q (n_0_2), .CK (n_0_40), .D (sph_n117));
DFF_X1 \b_reg[15]  (.Q (n_0_1), .CK (n_0_40), .D (sph_n142));
DFF_X1 \b_reg[16]  (.Q (n_0_0), .CK (n_0_40), .D (sph_n212));
DFF_X1 \b_reg[17]  (.Q (n_0_105), .CK (n_0_40), .D (sph_n257));
DFF_X1 \b_reg[18]  (.Q (n_0_104), .CK (n_0_40), .D (sph_n132));
DFF_X1 \b_reg[19]  (.Q (n_0_103), .CK (n_0_40), .D (sph_n67));
DFF_X1 \b_reg[20]  (.Q (n_0_102), .CK (n_0_40), .D (sph_n72));
DFF_X1 \b_reg[21]  (.Q (n_0_101), .CK (n_0_40), .D (sph_n42));
DFF_X1 \b_reg[22]  (.Q (n_0_100), .CK (n_0_40), .D (sph_n317));
DFF_X1 \c_out_reg[0]  (.Q (c_out[0]), .CK (n_0_50), .D (n_0_59));
DFF_X1 \c_out_reg[1]  (.Q (c_out[1]), .CK (n_0_50), .D (n_0_60));
DFF_X1 \c_out_reg[2]  (.Q (c_out[2]), .CK (n_0_50), .D (n_0_61));
DFF_X1 \c_out_reg[3]  (.Q (c_out[3]), .CK (n_0_50), .D (n_0_62));
DFF_X1 \c_out_reg[4]  (.Q (c_out[4]), .CK (n_0_50), .D (n_0_63));
DFF_X1 \c_out_reg[5]  (.Q (c_out[5]), .CK (n_0_50), .D (n_0_64));
DFF_X1 \c_out_reg[6]  (.Q (c_out[6]), .CK (n_0_50), .D (n_0_65));
DFF_X1 \c_out_reg[7]  (.Q (c_out[7]), .CK (n_0_50), .D (n_0_66));
DFF_X1 \c_out_reg[8]  (.Q (c_out[8]), .CK (n_0_50), .D (n_0_67));
DFF_X1 \c_out_reg[9]  (.Q (c_out[9]), .CK (n_0_50), .D (n_0_68));
DFF_X1 \c_out_reg[10]  (.Q (c_out[10]), .CK (n_0_50), .D (n_0_69));
DFF_X1 \c_out_reg[11]  (.Q (c_out[11]), .CK (n_0_50), .D (n_0_70));
DFF_X1 \c_out_reg[12]  (.Q (c_out[12]), .CK (n_0_50), .D (n_0_71));
DFF_X1 \c_out_reg[13]  (.Q (c_out[13]), .CK (n_0_50), .D (n_0_72));
DFF_X1 \c_out_reg[14]  (.Q (c_out[14]), .CK (n_0_50), .D (n_0_73));
DFF_X1 \c_out_reg[15]  (.Q (c_out[15]), .CK (n_0_50), .D (n_0_74));
DFF_X1 \c_out_reg[16]  (.Q (c_out[16]), .CK (n_0_50), .D (n_0_75));
DFF_X1 \c_out_reg[17]  (.Q (c_out[17]), .CK (n_0_50), .D (n_0_76));
DFF_X1 \c_out_reg[18]  (.Q (c_out[18]), .CK (n_0_50), .D (n_0_77));
DFF_X1 \c_out_reg[19]  (.Q (c_out[19]), .CK (n_0_50), .D (n_0_78));
DFF_X1 \c_out_reg[20]  (.Q (c_out[20]), .CK (n_0_50), .D (n_0_79));
DFF_X1 \c_out_reg[21]  (.Q (c_out[21]), .CK (n_0_50), .D (n_0_80));
DFF_X1 \c_out_reg[22]  (.Q (c_out[22]), .CK (n_0_50), .D (n_0_81));
DFF_X1 \c_out_reg[23]  (.Q (c_out[23]), .CK (n_0_50), .D (n_0_82));
DFF_X1 \c_out_reg[24]  (.Q (c_out[24]), .CK (n_0_50), .D (n_0_83));
DFF_X1 \c_out_reg[25]  (.Q (c_out[25]), .CK (n_0_50), .D (n_0_84));
DFF_X1 \c_out_reg[26]  (.Q (c_out[26]), .CK (n_0_50), .D (n_0_85));
DFF_X1 \c_out_reg[27]  (.Q (c_out[27]), .CK (n_0_50), .D (n_0_86));
DFF_X1 \c_out_reg[28]  (.Q (c_out[28]), .CK (n_0_50), .D (n_0_87));
DFF_X1 \c_out_reg[29]  (.Q (c_out[29]), .CK (n_0_50), .D (n_0_88));
DFF_X1 \c_out_reg[30]  (.Q (c_out[30]), .CK (n_0_50), .D (n_0_89));
DFF_X1 \c_out_reg[31]  (.Q (c_out[31]), .CK (n_0_50), .D (n_0_90));
DFF_X1 overflow_reg (.Q (overflow), .CK (n_0_50), .D (n_0_98));
unsigned_seq_multiplier unsigned_seq_multiplier_dut (.c ({uc_2, uc_3, \res_mant[23] , 
    \res_mant[22] , \res_mant[21] , \res_mant[20] , \res_mant[19] , \res_mant[18] , 
    \res_mant[17] , \res_mant[16] , \res_mant[15] , \res_mant[14] , \res_mant[13] , 
    \res_mant[12] , \res_mant[11] , \res_mant[10] , \res_mant[9] , \res_mant[8] , 
    \res_mant[7] , \res_mant[6] , \res_mant[5] , \res_mant[4] , \res_mant[3] , \res_mant[2] , 
    \res_mant[1] , uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, 
    uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, 
    uc_25, uc_26}), .a ({uc_0, n_0_17, n_0_18, n_0_19, n_0_20, n_0_21, n_0_22, n_0_23, 
    n_0_24, n_0_25, n_0_26, n_0_27, n_0_28, n_0_29, n_0_30, n_0_31, n_0_32, n_0_33, 
    n_0_34, n_0_35, n_0_36, n_0_37, n_0_38, n_0_39}), .b ({uc_1, n_0_100, n_0_101, 
    n_0_102, n_0_103, n_0_104, n_0_105, n_0_0, n_0_1, n_0_2, n_0_3, n_0_4, n_0_5, 
    n_0_6, n_0_7, n_0_8, n_0_9, n_0_10, n_0_11, n_0_12, n_0_13, n_0_14, n_0_15, n_0_16})
    , .clk (clk), .rst (rst), .start_s (mul_start));
BUF_X8 sps__L1_c1_c1 (.Z (mul_start), .A (sps__n1));
CLKBUF_X1 sph__c3 (.Z (sph_n7), .A (b_s[13]));
CLKBUF_X1 sph__c5 (.Z (sph_n12), .A (a_s[16]));
CLKBUF_X1 sph__c7 (.Z (sph_n17), .A (b_s[29]));
CLKBUF_X1 sph__c9 (.Z (sph_n22), .A (a_s[11]));
CLKBUF_X1 sph__c11 (.Z (sph_n27), .A (b_s[23]));
CLKBUF_X1 sph__c13 (.Z (sph_n32), .A (a_s[0]));
CLKBUF_X1 sph__c15 (.Z (sph_n37), .A (a_s[15]));
CLKBUF_X1 sph__c17 (.Z (sph_n42), .A (b_s[21]));
CLKBUF_X1 sph__c19 (.Z (sph_n47), .A (a_s[1]));
CLKBUF_X1 sph__c21 (.Z (sph_n52), .A (b_s[12]));
CLKBUF_X1 sph__c23 (.Z (sph_n57), .A (b_s[26]));
CLKBUF_X1 sph__c25 (.Z (sph_n62), .A (b_s[28]));
CLKBUF_X1 sph__c27 (.Z (sph_n67), .A (b_s[19]));
CLKBUF_X1 sph__c29 (.Z (sph_n72), .A (b_s[20]));
CLKBUF_X1 sph__c31 (.Z (sph_n77), .A (a_s[23]));
CLKBUF_X1 sph__c33 (.Z (sph_n82), .A (a_s[31]));
CLKBUF_X1 sph__c35 (.Z (sph_n87), .A (b_s[30]));
CLKBUF_X1 sph__c37 (.Z (sph_n92), .A (a_s[17]));
CLKBUF_X1 sph__c39 (.Z (sph_n97), .A (b_s[5]));
CLKBUF_X1 sph__c41 (.Z (sph_n102), .A (a_s[28]));
CLKBUF_X1 sph__c43 (.Z (sph_n107), .A (b_s[24]));
CLKBUF_X1 sph__c45 (.Z (sph_n112), .A (a_s[10]));
CLKBUF_X1 sph__c47 (.Z (sph_n117), .A (b_s[14]));
CLKBUF_X1 sph__c49 (.Z (sph_n122), .A (b_s[27]));
CLKBUF_X1 sph__c51 (.Z (sph_n127), .A (a_s[2]));
CLKBUF_X1 sph__c53 (.Z (sph_n132), .A (b_s[18]));
CLKBUF_X1 sph__c55 (.Z (sph_n137), .A (b_s[6]));
CLKBUF_X1 sph__c57 (.Z (sph_n142), .A (b_s[15]));
CLKBUF_X1 sph__c59 (.Z (sph_n147), .A (a_s[24]));
CLKBUF_X1 sph__c61 (.Z (sph_n152), .A (a_s[18]));
CLKBUF_X1 sph__c63 (.Z (sph_n157), .A (a_s[26]));
CLKBUF_X1 sph__c65 (.Z (sph_n162), .A (a_s[19]));
CLKBUF_X1 sph__c67 (.Z (sph_n167), .A (b_s[1]));
CLKBUF_X1 sph__c69 (.Z (sph_n172), .A (b_s[11]));
CLKBUF_X1 sph__c71 (.Z (sph_n177), .A (b_s[8]));
CLKBUF_X1 sph__c73 (.Z (sph_n182), .A (b_s[0]));
CLKBUF_X1 sph__c75 (.Z (sph_n187), .A (a_s[20]));
CLKBUF_X1 sph__c77 (.Z (sph_n192), .A (b_s[2]));
CLKBUF_X1 sph__c79 (.Z (sph_n197), .A (b_s[10]));
CLKBUF_X1 sph__c81 (.Z (sph_n202), .A (b_s[4]));
CLKBUF_X1 sph__c83 (.Z (sph_n207), .A (b_s[9]));
CLKBUF_X1 sph__c85 (.Z (sph_n212), .A (b_s[16]));
CLKBUF_X1 sph__c87 (.Z (sph_n217), .A (a_s[29]));
CLKBUF_X1 sph__c89 (.Z (sph_n222), .A (a_s[5]));
CLKBUF_X1 sph__c91 (.Z (sph_n227), .A (a_s[27]));
CLKBUF_X1 sph__c93 (.Z (sph_n232), .A (a_s[30]));
CLKBUF_X1 sph__c95 (.Z (sph_n237), .A (a_s[4]));
CLKBUF_X1 sph__c97 (.Z (sph_n242), .A (a_s[25]));
CLKBUF_X1 sph__c99 (.Z (sph_n247), .A (b_s[7]));
CLKBUF_X1 sph__c101 (.Z (sph_n252), .A (a_s[9]));
CLKBUF_X1 sph__c103 (.Z (sph_n257), .A (b_s[17]));
CLKBUF_X1 sph__c105 (.Z (sph_n262), .A (a_s[21]));
CLKBUF_X1 sph__c107 (.Z (sph_n267), .A (a_s[8]));
CLKBUF_X1 sph__c109 (.Z (sph_n272), .A (b_s[3]));
CLKBUF_X1 sph__c111 (.Z (sph_n277), .A (a_s[7]));
CLKBUF_X1 sph__c113 (.Z (sph_n282), .A (a_s[3]));
CLKBUF_X1 sph__c115 (.Z (sph_n287), .A (b_s[25]));
CLKBUF_X1 sph__c117 (.Z (sph_n292), .A (a_s[22]));
CLKBUF_X1 sph__c119 (.Z (sph_n297), .A (a_s[6]));
CLKBUF_X1 sph__c121 (.Z (sph_n302), .A (a_s[13]));
CLKBUF_X1 sph__c123 (.Z (sph_n307), .A (a_s[14]));
CLKBUF_X1 sph__c125 (.Z (sph_n312), .A (a_s[12]));
CLKBUF_X1 sph__c127 (.Z (sph_n317), .A (b_s[22]));
CLKBUF_X1 sph__c129 (.Z (sph_n322), .A (b_s[31]));

endmodule //fp_mul


