/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 23:22:53 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1544719207 */

module datapath(p_0, p_1, Accumulator);
   input [63:0]p_0;
   input [63:0]p_1;
   output [63:0]Accumulator;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(Accumulator[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(Accumulator[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(Accumulator[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(Accumulator[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(Accumulator[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(Accumulator[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(Accumulator[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(Accumulator[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(Accumulator[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(Accumulator[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(Accumulator[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(
      Accumulator[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(
      Accumulator[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(
      Accumulator[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(
      Accumulator[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(
      Accumulator[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(
      Accumulator[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(
      Accumulator[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(
      Accumulator[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(
      Accumulator[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(
      Accumulator[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(
      Accumulator[21]));
   FA_X1 i_22 (.A(p_0[22]), .B(p_1[22]), .CI(n_21), .CO(n_22), .S(
      Accumulator[22]));
   FA_X1 i_23 (.A(p_0[23]), .B(p_1[23]), .CI(n_22), .CO(n_23), .S(
      Accumulator[23]));
   FA_X1 i_24 (.A(p_0[24]), .B(p_1[24]), .CI(n_23), .CO(n_24), .S(
      Accumulator[24]));
   FA_X1 i_25 (.A(p_0[25]), .B(p_1[25]), .CI(n_24), .CO(n_25), .S(
      Accumulator[25]));
   FA_X1 i_26 (.A(p_0[26]), .B(p_1[26]), .CI(n_25), .CO(n_26), .S(
      Accumulator[26]));
   FA_X1 i_27 (.A(p_0[27]), .B(p_1[27]), .CI(n_26), .CO(n_27), .S(
      Accumulator[27]));
   FA_X1 i_28 (.A(p_0[28]), .B(p_1[28]), .CI(n_27), .CO(n_28), .S(
      Accumulator[28]));
   FA_X1 i_29 (.A(p_0[29]), .B(p_1[29]), .CI(n_28), .CO(n_29), .S(
      Accumulator[29]));
   FA_X1 i_30 (.A(p_0[30]), .B(p_1[30]), .CI(n_29), .CO(n_30), .S(
      Accumulator[30]));
   FA_X1 i_31 (.A(p_0[31]), .B(p_1[31]), .CI(n_30), .CO(n_31), .S(
      Accumulator[31]));
   FA_X1 i_32 (.A(p_0[32]), .B(p_1[32]), .CI(n_31), .CO(n_32), .S(
      Accumulator[32]));
   FA_X1 i_33 (.A(p_0[33]), .B(p_1[33]), .CI(n_32), .CO(n_33), .S(
      Accumulator[33]));
   FA_X1 i_34 (.A(p_0[34]), .B(p_1[34]), .CI(n_33), .CO(n_34), .S(
      Accumulator[34]));
   FA_X1 i_35 (.A(p_0[35]), .B(p_1[35]), .CI(n_34), .CO(n_35), .S(
      Accumulator[35]));
   FA_X1 i_36 (.A(p_0[36]), .B(p_1[36]), .CI(n_35), .CO(n_36), .S(
      Accumulator[36]));
   FA_X1 i_37 (.A(p_0[37]), .B(p_1[37]), .CI(n_36), .CO(n_37), .S(
      Accumulator[37]));
   FA_X1 i_38 (.A(p_0[38]), .B(p_1[38]), .CI(n_37), .CO(n_38), .S(
      Accumulator[38]));
   FA_X1 i_39 (.A(p_0[39]), .B(p_1[39]), .CI(n_38), .CO(n_39), .S(
      Accumulator[39]));
   FA_X1 i_40 (.A(p_0[40]), .B(p_1[40]), .CI(n_39), .CO(n_40), .S(
      Accumulator[40]));
   FA_X1 i_41 (.A(p_0[41]), .B(p_1[41]), .CI(n_40), .CO(n_41), .S(
      Accumulator[41]));
   FA_X1 i_42 (.A(p_0[42]), .B(p_1[42]), .CI(n_41), .CO(n_42), .S(
      Accumulator[42]));
   FA_X1 i_43 (.A(p_0[43]), .B(p_1[43]), .CI(n_42), .CO(n_43), .S(
      Accumulator[43]));
   FA_X1 i_44 (.A(p_0[44]), .B(p_1[44]), .CI(n_43), .CO(n_44), .S(
      Accumulator[44]));
   FA_X1 i_45 (.A(p_0[45]), .B(p_1[45]), .CI(n_44), .CO(n_45), .S(
      Accumulator[45]));
   FA_X1 i_46 (.A(p_0[46]), .B(p_1[46]), .CI(n_45), .CO(n_46), .S(
      Accumulator[46]));
   FA_X1 i_47 (.A(p_0[47]), .B(p_1[47]), .CI(n_46), .CO(n_47), .S(
      Accumulator[47]));
   FA_X1 i_48 (.A(p_0[48]), .B(p_1[48]), .CI(n_47), .CO(n_48), .S(
      Accumulator[48]));
   FA_X1 i_49 (.A(p_0[49]), .B(p_1[49]), .CI(n_48), .CO(n_49), .S(
      Accumulator[49]));
   FA_X1 i_50 (.A(p_0[50]), .B(p_1[50]), .CI(n_49), .CO(n_50), .S(
      Accumulator[50]));
   FA_X1 i_51 (.A(p_0[51]), .B(p_1[51]), .CI(n_50), .CO(n_51), .S(
      Accumulator[51]));
   FA_X1 i_52 (.A(p_0[52]), .B(p_1[52]), .CI(n_51), .CO(n_52), .S(
      Accumulator[52]));
   FA_X1 i_53 (.A(p_0[53]), .B(p_1[53]), .CI(n_52), .CO(n_53), .S(
      Accumulator[53]));
   FA_X1 i_54 (.A(p_0[54]), .B(p_1[54]), .CI(n_53), .CO(n_54), .S(
      Accumulator[54]));
   FA_X1 i_55 (.A(p_0[55]), .B(p_1[55]), .CI(n_54), .CO(n_55), .S(
      Accumulator[55]));
   FA_X1 i_56 (.A(p_0[56]), .B(p_1[56]), .CI(n_55), .CO(n_56), .S(
      Accumulator[56]));
   FA_X1 i_57 (.A(p_0[57]), .B(p_1[57]), .CI(n_56), .CO(n_57), .S(
      Accumulator[57]));
   FA_X1 i_58 (.A(p_0[58]), .B(p_1[58]), .CI(n_57), .CO(n_58), .S(
      Accumulator[58]));
   FA_X1 i_59 (.A(p_0[59]), .B(p_1[59]), .CI(n_58), .CO(n_59), .S(
      Accumulator[59]));
   FA_X1 i_60 (.A(p_0[60]), .B(p_1[60]), .CI(n_59), .CO(n_60), .S(
      Accumulator[60]));
   FA_X1 i_61 (.A(p_0[61]), .B(p_1[61]), .CI(n_60), .CO(n_61), .S(
      Accumulator[61]));
   FA_X1 i_62 (.A(p_0[62]), .B(p_1[62]), .CI(n_61), .CO(n_62), .S(
      Accumulator[62]));
   XNOR2_X1 i_63 (.A(p_0[63]), .B(p_1[63]), .ZN(n_63));
   XNOR2_X1 i_64 (.A(n_63), .B(n_62), .ZN(Accumulator[63]));
endmodule

module seq_multiplier_v2(clk, rst, a, b, c);
   input clk;
   input rst;
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   wire n_0_0;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire [7:0]counter;
   wire [63:0]B;
   wire [63:0]Q;
   wire [63:0]Accumulator;
   wire n_0_1;
   wire n_0_0_6;
   wire n_0_0_0;
   wire n_0_0_7;
   wire n_0_0_1;
   wire n_0_0_8;
   wire n_0_0_2;
   wire n_0_0_9;
   wire n_0_0_3;
   wire n_0_0_10;
   wire n_0_0_4;
   wire n_0_0_11;
   wire n_0_0_5;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_3;
   wire n_0_195;
   wire n_0_4;
   wire n_0_0_12;
   wire n_0_5;
   wire n_0_0_13;
   wire n_0_6;
   wire n_0_0_14;
   wire n_0_7;
   wire n_0_0_15;
   wire n_0_8;
   wire n_0_0_16;
   wire n_0_9;
   wire n_0_0_17;
   wire n_0_10;
   wire n_0_0_18;
   wire n_0_11;
   wire n_0_0_19;
   wire n_0_12;
   wire n_0_0_20;
   wire n_0_13;
   wire n_0_0_21;
   wire n_0_14;
   wire n_0_0_22;
   wire n_0_15;
   wire n_0_0_23;
   wire n_0_16;
   wire n_0_0_24;
   wire n_0_17;
   wire n_0_0_25;
   wire n_0_18;
   wire n_0_0_26;
   wire n_0_19;
   wire n_0_0_27;
   wire n_0_20;
   wire n_0_0_28;
   wire n_0_21;
   wire n_0_0_29;
   wire n_0_22;
   wire n_0_0_30;
   wire n_0_23;
   wire n_0_0_31;
   wire n_0_24;
   wire n_0_0_32;
   wire n_0_25;
   wire n_0_0_33;
   wire n_0_26;
   wire n_0_0_34;
   wire n_0_27;
   wire n_0_0_35;
   wire n_0_28;
   wire n_0_0_36;
   wire n_0_29;
   wire n_0_0_37;
   wire n_0_30;
   wire n_0_0_38;
   wire n_0_31;
   wire n_0_0_39;
   wire n_0_32;
   wire n_0_0_40;
   wire n_0_33;
   wire n_0_0_41;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_2;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_289;
   wire n_0_290;
   wire n_0_0_87;

   CLKGATETST_X1 clk_gate_c_reg (.CK(clk), .E(n_0_2), .SE(1'b0), .GCK(n_0_0));
   DFFR_X1 \c_reg[63]  (.D(n_0_194), .RN(n_0_289), .CK(n_0_0), .Q(c[63]), .QN());
   DFFR_X1 \c_reg[62]  (.D(n_0_193), .RN(n_0_289), .CK(n_0_0), .Q(c[62]), .QN());
   DFFR_X1 \c_reg[61]  (.D(n_0_192), .RN(n_0_289), .CK(n_0_0), .Q(c[61]), .QN());
   DFFR_X1 \c_reg[60]  (.D(n_0_191), .RN(n_0_289), .CK(n_0_0), .Q(c[60]), .QN());
   DFFR_X1 \c_reg[59]  (.D(n_0_190), .RN(n_0_289), .CK(n_0_0), .Q(c[59]), .QN());
   DFFR_X1 \c_reg[58]  (.D(n_0_189), .RN(n_0_289), .CK(n_0_0), .Q(c[58]), .QN());
   DFFR_X1 \c_reg[57]  (.D(n_0_188), .RN(n_0_289), .CK(n_0_0), .Q(c[57]), .QN());
   DFFR_X1 \c_reg[56]  (.D(n_0_187), .RN(n_0_289), .CK(n_0_0), .Q(c[56]), .QN());
   DFFR_X1 \c_reg[55]  (.D(n_0_186), .RN(n_0_289), .CK(n_0_0), .Q(c[55]), .QN());
   DFFR_X1 \c_reg[54]  (.D(n_0_185), .RN(n_0_289), .CK(n_0_0), .Q(c[54]), .QN());
   DFFR_X1 \c_reg[53]  (.D(n_0_184), .RN(n_0_289), .CK(n_0_0), .Q(c[53]), .QN());
   DFFR_X1 \c_reg[52]  (.D(n_0_183), .RN(n_0_289), .CK(n_0_0), .Q(c[52]), .QN());
   DFFR_X1 \c_reg[51]  (.D(n_0_182), .RN(n_0_289), .CK(n_0_0), .Q(c[51]), .QN());
   DFFR_X1 \c_reg[50]  (.D(n_0_181), .RN(n_0_289), .CK(n_0_0), .Q(c[50]), .QN());
   DFFR_X1 \c_reg[49]  (.D(n_0_180), .RN(n_0_289), .CK(n_0_0), .Q(c[49]), .QN());
   DFFR_X1 \c_reg[48]  (.D(n_0_179), .RN(n_0_289), .CK(n_0_0), .Q(c[48]), .QN());
   DFFR_X1 \c_reg[47]  (.D(n_0_178), .RN(n_0_289), .CK(n_0_0), .Q(c[47]), .QN());
   DFFR_X1 \c_reg[46]  (.D(n_0_177), .RN(n_0_289), .CK(n_0_0), .Q(c[46]), .QN());
   DFFR_X1 \c_reg[45]  (.D(n_0_176), .RN(n_0_289), .CK(n_0_0), .Q(c[45]), .QN());
   DFFR_X1 \c_reg[44]  (.D(n_0_175), .RN(n_0_289), .CK(n_0_0), .Q(c[44]), .QN());
   DFFR_X1 \c_reg[43]  (.D(n_0_174), .RN(n_0_289), .CK(n_0_0), .Q(c[43]), .QN());
   DFFR_X1 \c_reg[42]  (.D(n_0_173), .RN(n_0_289), .CK(n_0_0), .Q(c[42]), .QN());
   DFFR_X1 \c_reg[41]  (.D(n_0_172), .RN(n_0_289), .CK(n_0_0), .Q(c[41]), .QN());
   DFFR_X1 \c_reg[40]  (.D(n_0_171), .RN(n_0_289), .CK(n_0_0), .Q(c[40]), .QN());
   DFFR_X1 \c_reg[39]  (.D(n_0_170), .RN(n_0_289), .CK(n_0_0), .Q(c[39]), .QN());
   DFFR_X1 \c_reg[38]  (.D(n_0_169), .RN(n_0_289), .CK(n_0_0), .Q(c[38]), .QN());
   DFFR_X1 \c_reg[37]  (.D(n_0_168), .RN(n_0_289), .CK(n_0_0), .Q(c[37]), .QN());
   DFFR_X1 \c_reg[36]  (.D(n_0_167), .RN(n_0_289), .CK(n_0_0), .Q(c[36]), .QN());
   DFFR_X1 \c_reg[35]  (.D(n_0_166), .RN(n_0_289), .CK(n_0_0), .Q(c[35]), .QN());
   DFFR_X1 \c_reg[34]  (.D(n_0_165), .RN(n_0_289), .CK(n_0_0), .Q(c[34]), .QN());
   DFFR_X1 \c_reg[33]  (.D(n_0_164), .RN(n_0_289), .CK(n_0_0), .Q(c[33]), .QN());
   DFFR_X1 \c_reg[32]  (.D(n_0_163), .RN(n_0_289), .CK(n_0_0), .Q(c[32]), .QN());
   DFFR_X1 \c_reg[31]  (.D(n_0_162), .RN(n_0_289), .CK(n_0_0), .Q(c[31]), .QN());
   DFFR_X1 \c_reg[30]  (.D(n_0_161), .RN(n_0_289), .CK(n_0_0), .Q(c[30]), .QN());
   DFFR_X1 \c_reg[29]  (.D(n_0_160), .RN(n_0_289), .CK(n_0_0), .Q(c[29]), .QN());
   DFFR_X1 \c_reg[28]  (.D(n_0_159), .RN(n_0_289), .CK(n_0_0), .Q(c[28]), .QN());
   DFFR_X1 \c_reg[27]  (.D(n_0_158), .RN(n_0_289), .CK(n_0_0), .Q(c[27]), .QN());
   DFFR_X1 \c_reg[26]  (.D(n_0_157), .RN(n_0_289), .CK(n_0_0), .Q(c[26]), .QN());
   DFFR_X1 \c_reg[25]  (.D(n_0_156), .RN(n_0_289), .CK(n_0_0), .Q(c[25]), .QN());
   DFFR_X1 \c_reg[24]  (.D(n_0_155), .RN(n_0_289), .CK(n_0_0), .Q(c[24]), .QN());
   DFFR_X1 \c_reg[23]  (.D(n_0_154), .RN(n_0_289), .CK(n_0_0), .Q(c[23]), .QN());
   DFFR_X1 \c_reg[22]  (.D(n_0_153), .RN(n_0_289), .CK(n_0_0), .Q(c[22]), .QN());
   DFFR_X1 \c_reg[21]  (.D(n_0_152), .RN(n_0_289), .CK(n_0_0), .Q(c[21]), .QN());
   DFFR_X1 \c_reg[20]  (.D(n_0_151), .RN(n_0_289), .CK(n_0_0), .Q(c[20]), .QN());
   DFFR_X1 \c_reg[19]  (.D(n_0_150), .RN(n_0_289), .CK(n_0_0), .Q(c[19]), .QN());
   DFFR_X1 \c_reg[18]  (.D(n_0_149), .RN(n_0_289), .CK(n_0_0), .Q(c[18]), .QN());
   DFFR_X1 \c_reg[17]  (.D(n_0_148), .RN(n_0_289), .CK(n_0_0), .Q(c[17]), .QN());
   DFFR_X1 \c_reg[16]  (.D(n_0_147), .RN(n_0_289), .CK(n_0_0), .Q(c[16]), .QN());
   DFFR_X1 \c_reg[15]  (.D(n_0_146), .RN(n_0_289), .CK(n_0_0), .Q(c[15]), .QN());
   DFFR_X1 \c_reg[14]  (.D(n_0_145), .RN(n_0_289), .CK(n_0_0), .Q(c[14]), .QN());
   DFFR_X1 \c_reg[13]  (.D(n_0_144), .RN(n_0_289), .CK(n_0_0), .Q(c[13]), .QN());
   DFFR_X1 \c_reg[12]  (.D(n_0_143), .RN(n_0_289), .CK(n_0_0), .Q(c[12]), .QN());
   DFFR_X1 \c_reg[11]  (.D(n_0_142), .RN(n_0_289), .CK(n_0_0), .Q(c[11]), .QN());
   DFFR_X1 \c_reg[10]  (.D(n_0_141), .RN(n_0_289), .CK(n_0_0), .Q(c[10]), .QN());
   DFFR_X1 \c_reg[9]  (.D(n_0_140), .RN(n_0_289), .CK(n_0_0), .Q(c[9]), .QN());
   DFFR_X1 \c_reg[8]  (.D(n_0_139), .RN(n_0_289), .CK(n_0_0), .Q(c[8]), .QN());
   DFFR_X1 \c_reg[7]  (.D(n_0_138), .RN(n_0_289), .CK(n_0_0), .Q(c[7]), .QN());
   DFFR_X1 \c_reg[6]  (.D(n_0_137), .RN(n_0_289), .CK(n_0_0), .Q(c[6]), .QN());
   DFFR_X1 \c_reg[5]  (.D(n_0_136), .RN(n_0_289), .CK(n_0_0), .Q(c[5]), .QN());
   DFFR_X1 \c_reg[4]  (.D(n_0_135), .RN(n_0_289), .CK(n_0_0), .Q(c[4]), .QN());
   DFFR_X1 \c_reg[3]  (.D(n_0_134), .RN(n_0_289), .CK(n_0_0), .Q(c[3]), .QN());
   DFFR_X1 \c_reg[2]  (.D(n_0_133), .RN(n_0_289), .CK(n_0_0), .Q(c[2]), .QN());
   DFFR_X1 \c_reg[1]  (.D(n_0_132), .RN(n_0_289), .CK(n_0_0), .Q(c[1]), .QN());
   DFFR_X1 \c_reg[0]  (.D(n_0_131), .RN(n_0_289), .CK(n_0_0), .Q(c[0]), .QN());
   datapath i_0_4 (.p_0({n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, 
      n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, 
      n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, 
      n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, 
      n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, 
      n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, 
      n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, 
      n_0_4, n_0_3}), .p_1({n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, 
      n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, 
      n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, 
      n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, 
      n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, 
      n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, 
      n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, 
      n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67}), .Accumulator({
      n_0_194, n_0_193, n_0_192, n_0_191, n_0_190, n_0_189, n_0_188, n_0_187, 
      n_0_186, n_0_185, n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, 
      n_0_178, n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, 
      n_0_170, n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, 
      n_0_162, n_0_161, n_0_160, n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, 
      n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, 
      n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, n_0_141, n_0_140, n_0_139, 
      n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, n_0_133, n_0_132, n_0_131}));
   DFFR_X1 \counter_reg[7]  (.D(n_0_297), .RN(n_0_289), .CK(clk), .Q(counter[7]), 
      .QN());
   DFFR_X1 \counter_reg[6]  (.D(n_0_296), .RN(n_0_289), .CK(clk), .Q(counter[6]), 
      .QN());
   DFFR_X1 \counter_reg[5]  (.D(n_0_295), .RN(n_0_289), .CK(clk), .Q(counter[5]), 
      .QN());
   DFFR_X1 \counter_reg[4]  (.D(n_0_294), .RN(n_0_289), .CK(clk), .Q(counter[4]), 
      .QN());
   DFFR_X1 \counter_reg[3]  (.D(n_0_293), .RN(n_0_289), .CK(clk), .Q(counter[3]), 
      .QN());
   DFFR_X1 \counter_reg[2]  (.D(n_0_292), .RN(n_0_289), .CK(clk), .Q(counter[2]), 
      .QN());
   DFFR_X1 \counter_reg[1]  (.D(n_0_291), .RN(n_0_289), .CK(clk), .Q(counter[1]), 
      .QN());
   DFFR_X1 \counter_reg[0]  (.D(n_0_290), .RN(n_0_289), .CK(clk), .Q(counter[0]), 
      .QN());
   DFF_X1 \B_reg[63]  (.D(n_0_257), .CK(n_0_1), .Q(B[63]), .QN());
   DFF_X1 \B_reg[62]  (.D(n_0_256), .CK(n_0_1), .Q(B[62]), .QN());
   DFF_X1 \B_reg[61]  (.D(n_0_255), .CK(n_0_1), .Q(B[61]), .QN());
   DFF_X1 \B_reg[60]  (.D(n_0_254), .CK(n_0_1), .Q(B[60]), .QN());
   DFF_X1 \B_reg[59]  (.D(n_0_253), .CK(n_0_1), .Q(B[59]), .QN());
   DFF_X1 \B_reg[58]  (.D(n_0_252), .CK(n_0_1), .Q(B[58]), .QN());
   DFF_X1 \B_reg[57]  (.D(n_0_251), .CK(n_0_1), .Q(B[57]), .QN());
   DFF_X1 \B_reg[56]  (.D(n_0_250), .CK(n_0_1), .Q(B[56]), .QN());
   DFF_X1 \B_reg[55]  (.D(n_0_249), .CK(n_0_1), .Q(B[55]), .QN());
   DFF_X1 \B_reg[54]  (.D(n_0_248), .CK(n_0_1), .Q(B[54]), .QN());
   DFF_X1 \B_reg[53]  (.D(n_0_247), .CK(n_0_1), .Q(B[53]), .QN());
   DFF_X1 \B_reg[52]  (.D(n_0_246), .CK(n_0_1), .Q(B[52]), .QN());
   DFF_X1 \B_reg[51]  (.D(n_0_245), .CK(n_0_1), .Q(B[51]), .QN());
   DFF_X1 \B_reg[50]  (.D(n_0_244), .CK(n_0_1), .Q(B[50]), .QN());
   DFF_X1 \B_reg[49]  (.D(n_0_243), .CK(n_0_1), .Q(B[49]), .QN());
   DFF_X1 \B_reg[48]  (.D(n_0_242), .CK(n_0_1), .Q(B[48]), .QN());
   DFF_X1 \B_reg[47]  (.D(n_0_241), .CK(n_0_1), .Q(B[47]), .QN());
   DFF_X1 \B_reg[46]  (.D(n_0_240), .CK(n_0_1), .Q(B[46]), .QN());
   DFF_X1 \B_reg[45]  (.D(n_0_239), .CK(n_0_1), .Q(B[45]), .QN());
   DFF_X1 \B_reg[44]  (.D(n_0_238), .CK(n_0_1), .Q(B[44]), .QN());
   DFF_X1 \B_reg[43]  (.D(n_0_237), .CK(n_0_1), .Q(B[43]), .QN());
   DFF_X1 \B_reg[42]  (.D(n_0_236), .CK(n_0_1), .Q(B[42]), .QN());
   DFF_X1 \B_reg[41]  (.D(n_0_235), .CK(n_0_1), .Q(B[41]), .QN());
   DFF_X1 \B_reg[40]  (.D(n_0_234), .CK(n_0_1), .Q(B[40]), .QN());
   DFF_X1 \B_reg[39]  (.D(n_0_233), .CK(n_0_1), .Q(B[39]), .QN());
   DFF_X1 \B_reg[38]  (.D(n_0_232), .CK(n_0_1), .Q(B[38]), .QN());
   DFF_X1 \B_reg[37]  (.D(n_0_231), .CK(n_0_1), .Q(B[37]), .QN());
   DFF_X1 \B_reg[36]  (.D(n_0_230), .CK(n_0_1), .Q(B[36]), .QN());
   DFF_X1 \B_reg[35]  (.D(n_0_229), .CK(n_0_1), .Q(B[35]), .QN());
   DFF_X1 \B_reg[34]  (.D(n_0_228), .CK(n_0_1), .Q(B[34]), .QN());
   DFF_X1 \B_reg[33]  (.D(n_0_227), .CK(n_0_1), .Q(B[33]), .QN());
   DFF_X1 \B_reg[32]  (.D(n_0_226), .CK(n_0_1), .Q(B[32]), .QN());
   DFF_X1 \B_reg[31]  (.D(n_0_225), .CK(n_0_1), .Q(B[31]), .QN());
   DFF_X1 \B_reg[30]  (.D(n_0_224), .CK(n_0_1), .Q(B[30]), .QN());
   DFF_X1 \B_reg[29]  (.D(n_0_223), .CK(n_0_1), .Q(B[29]), .QN());
   DFF_X1 \B_reg[28]  (.D(n_0_222), .CK(n_0_1), .Q(B[28]), .QN());
   DFF_X1 \B_reg[27]  (.D(n_0_221), .CK(n_0_1), .Q(B[27]), .QN());
   DFF_X1 \B_reg[26]  (.D(n_0_220), .CK(n_0_1), .Q(B[26]), .QN());
   DFF_X1 \B_reg[25]  (.D(n_0_219), .CK(n_0_1), .Q(B[25]), .QN());
   DFF_X1 \B_reg[24]  (.D(n_0_218), .CK(n_0_1), .Q(B[24]), .QN());
   DFF_X1 \B_reg[23]  (.D(n_0_217), .CK(n_0_1), .Q(B[23]), .QN());
   DFF_X1 \B_reg[22]  (.D(n_0_216), .CK(n_0_1), .Q(B[22]), .QN());
   DFF_X1 \B_reg[21]  (.D(n_0_215), .CK(n_0_1), .Q(B[21]), .QN());
   DFF_X1 \B_reg[20]  (.D(n_0_214), .CK(n_0_1), .Q(B[20]), .QN());
   DFF_X1 \B_reg[19]  (.D(n_0_213), .CK(n_0_1), .Q(B[19]), .QN());
   DFF_X1 \B_reg[18]  (.D(n_0_212), .CK(n_0_1), .Q(B[18]), .QN());
   DFF_X1 \B_reg[17]  (.D(n_0_211), .CK(n_0_1), .Q(B[17]), .QN());
   DFF_X1 \B_reg[16]  (.D(n_0_210), .CK(n_0_1), .Q(B[16]), .QN());
   DFF_X1 \B_reg[15]  (.D(n_0_209), .CK(n_0_1), .Q(B[15]), .QN());
   DFF_X1 \B_reg[14]  (.D(n_0_208), .CK(n_0_1), .Q(B[14]), .QN());
   DFF_X1 \B_reg[13]  (.D(n_0_207), .CK(n_0_1), .Q(B[13]), .QN());
   DFF_X1 \B_reg[12]  (.D(n_0_206), .CK(n_0_1), .Q(B[12]), .QN());
   DFF_X1 \B_reg[11]  (.D(n_0_205), .CK(n_0_1), .Q(B[11]), .QN());
   DFF_X1 \B_reg[10]  (.D(n_0_204), .CK(n_0_1), .Q(B[10]), .QN());
   DFF_X1 \B_reg[9]  (.D(n_0_203), .CK(n_0_1), .Q(B[9]), .QN());
   DFF_X1 \B_reg[8]  (.D(n_0_202), .CK(n_0_1), .Q(B[8]), .QN());
   DFF_X1 \B_reg[7]  (.D(n_0_201), .CK(n_0_1), .Q(B[7]), .QN());
   DFF_X1 \B_reg[6]  (.D(n_0_200), .CK(n_0_1), .Q(B[6]), .QN());
   DFF_X1 \B_reg[5]  (.D(n_0_199), .CK(n_0_1), .Q(B[5]), .QN());
   DFF_X1 \B_reg[4]  (.D(n_0_198), .CK(n_0_1), .Q(B[4]), .QN());
   DFF_X1 \B_reg[3]  (.D(n_0_197), .CK(n_0_1), .Q(B[3]), .QN());
   DFF_X1 \B_reg[2]  (.D(n_0_196), .CK(n_0_1), .Q(B[2]), .QN());
   DFF_X1 \B_reg[1]  (.D(n_0_195), .CK(n_0_1), .Q(B[1]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_0_288), .CK(n_0_1), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_0_287), .CK(n_0_1), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_0_286), .CK(n_0_1), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_0_285), .CK(n_0_1), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_0_284), .CK(n_0_1), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_0_283), .CK(n_0_1), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_0_282), .CK(n_0_1), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_0_281), .CK(n_0_1), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_0_280), .CK(n_0_1), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_0_279), .CK(n_0_1), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_0_278), .CK(n_0_1), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_0_277), .CK(n_0_1), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_0_276), .CK(n_0_1), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_0_275), .CK(n_0_1), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_0_274), .CK(n_0_1), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_0_273), .CK(n_0_1), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_0_272), .CK(n_0_1), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_0_271), .CK(n_0_1), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_0_270), .CK(n_0_1), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_0_269), .CK(n_0_1), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_0_268), .CK(n_0_1), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_0_267), .CK(n_0_1), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_0_266), .CK(n_0_1), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_0_265), .CK(n_0_1), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_0_264), .CK(n_0_1), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_0_263), .CK(n_0_1), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_0_262), .CK(n_0_1), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_0_261), .CK(n_0_1), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_0_260), .CK(n_0_1), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_0_259), .CK(n_0_1), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0_258), .CK(n_0_1), .Q(Q[0]), .QN());
   DFFR_X1 \Accumulator_reg[63]  (.D(n_0_194), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[63]), .QN());
   DFFR_X1 \Accumulator_reg[62]  (.D(n_0_193), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[62]), .QN());
   DFFR_X1 \Accumulator_reg[61]  (.D(n_0_192), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[61]), .QN());
   DFFR_X1 \Accumulator_reg[60]  (.D(n_0_191), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[60]), .QN());
   DFFR_X1 \Accumulator_reg[59]  (.D(n_0_190), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[59]), .QN());
   DFFR_X1 \Accumulator_reg[58]  (.D(n_0_189), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[58]), .QN());
   DFFR_X1 \Accumulator_reg[57]  (.D(n_0_188), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[57]), .QN());
   DFFR_X1 \Accumulator_reg[56]  (.D(n_0_187), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[56]), .QN());
   DFFR_X1 \Accumulator_reg[55]  (.D(n_0_186), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[55]), .QN());
   DFFR_X1 \Accumulator_reg[54]  (.D(n_0_185), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[54]), .QN());
   DFFR_X1 \Accumulator_reg[53]  (.D(n_0_184), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[53]), .QN());
   DFFR_X1 \Accumulator_reg[52]  (.D(n_0_183), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[52]), .QN());
   DFFR_X1 \Accumulator_reg[51]  (.D(n_0_182), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[51]), .QN());
   DFFR_X1 \Accumulator_reg[50]  (.D(n_0_181), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[50]), .QN());
   DFFR_X1 \Accumulator_reg[49]  (.D(n_0_180), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[49]), .QN());
   DFFR_X1 \Accumulator_reg[48]  (.D(n_0_179), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[48]), .QN());
   DFFR_X1 \Accumulator_reg[47]  (.D(n_0_178), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[47]), .QN());
   DFFR_X1 \Accumulator_reg[46]  (.D(n_0_177), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[46]), .QN());
   DFFR_X1 \Accumulator_reg[45]  (.D(n_0_176), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[45]), .QN());
   DFFR_X1 \Accumulator_reg[44]  (.D(n_0_175), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[44]), .QN());
   DFFR_X1 \Accumulator_reg[43]  (.D(n_0_174), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[43]), .QN());
   DFFR_X1 \Accumulator_reg[42]  (.D(n_0_173), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[42]), .QN());
   DFFR_X1 \Accumulator_reg[41]  (.D(n_0_172), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[41]), .QN());
   DFFR_X1 \Accumulator_reg[40]  (.D(n_0_171), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[40]), .QN());
   DFFR_X1 \Accumulator_reg[39]  (.D(n_0_170), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[39]), .QN());
   DFFR_X1 \Accumulator_reg[38]  (.D(n_0_169), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[38]), .QN());
   DFFR_X1 \Accumulator_reg[37]  (.D(n_0_168), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[37]), .QN());
   DFFR_X1 \Accumulator_reg[36]  (.D(n_0_167), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[36]), .QN());
   DFFR_X1 \Accumulator_reg[35]  (.D(n_0_166), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[35]), .QN());
   DFFR_X1 \Accumulator_reg[34]  (.D(n_0_165), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[34]), .QN());
   DFFR_X1 \Accumulator_reg[33]  (.D(n_0_164), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[33]), .QN());
   DFFR_X1 \Accumulator_reg[32]  (.D(n_0_163), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[32]), .QN());
   DFFR_X1 \Accumulator_reg[31]  (.D(n_0_162), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[31]), .QN());
   DFFR_X1 \Accumulator_reg[30]  (.D(n_0_161), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[30]), .QN());
   DFFR_X1 \Accumulator_reg[29]  (.D(n_0_160), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[29]), .QN());
   DFFR_X1 \Accumulator_reg[28]  (.D(n_0_159), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[28]), .QN());
   DFFR_X1 \Accumulator_reg[27]  (.D(n_0_158), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[27]), .QN());
   DFFR_X1 \Accumulator_reg[26]  (.D(n_0_157), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[26]), .QN());
   DFFR_X1 \Accumulator_reg[25]  (.D(n_0_156), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[25]), .QN());
   DFFR_X1 \Accumulator_reg[24]  (.D(n_0_155), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[24]), .QN());
   DFFR_X1 \Accumulator_reg[23]  (.D(n_0_154), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[23]), .QN());
   DFFR_X1 \Accumulator_reg[22]  (.D(n_0_153), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[22]), .QN());
   DFFR_X1 \Accumulator_reg[21]  (.D(n_0_152), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[21]), .QN());
   DFFR_X1 \Accumulator_reg[20]  (.D(n_0_151), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[20]), .QN());
   DFFR_X1 \Accumulator_reg[19]  (.D(n_0_150), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[19]), .QN());
   DFFR_X1 \Accumulator_reg[18]  (.D(n_0_149), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[18]), .QN());
   DFFR_X1 \Accumulator_reg[17]  (.D(n_0_148), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[17]), .QN());
   DFFR_X1 \Accumulator_reg[16]  (.D(n_0_147), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[16]), .QN());
   DFFR_X1 \Accumulator_reg[15]  (.D(n_0_146), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[15]), .QN());
   DFFR_X1 \Accumulator_reg[14]  (.D(n_0_145), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[14]), .QN());
   DFFR_X1 \Accumulator_reg[13]  (.D(n_0_144), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[13]), .QN());
   DFFR_X1 \Accumulator_reg[12]  (.D(n_0_143), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[12]), .QN());
   DFFR_X1 \Accumulator_reg[11]  (.D(n_0_142), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[11]), .QN());
   DFFR_X1 \Accumulator_reg[10]  (.D(n_0_141), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[10]), .QN());
   DFFR_X1 \Accumulator_reg[9]  (.D(n_0_140), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[9]), .QN());
   DFFR_X1 \Accumulator_reg[8]  (.D(n_0_139), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[8]), .QN());
   DFFR_X1 \Accumulator_reg[7]  (.D(n_0_138), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[7]), .QN());
   DFFR_X1 \Accumulator_reg[6]  (.D(n_0_137), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[6]), .QN());
   DFFR_X1 \Accumulator_reg[5]  (.D(n_0_136), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[5]), .QN());
   DFFR_X1 \Accumulator_reg[4]  (.D(n_0_135), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[4]), .QN());
   DFFR_X1 \Accumulator_reg[3]  (.D(n_0_134), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[3]), .QN());
   DFFR_X1 \Accumulator_reg[2]  (.D(n_0_133), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[2]), .QN());
   DFFR_X1 \Accumulator_reg[1]  (.D(n_0_132), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[1]), .QN());
   DFFR_X1 \Accumulator_reg[0]  (.D(n_0_131), .RN(n_0_289), .CK(clk), .Q(
      Accumulator[0]), .QN());
   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_0_289), .SE(1'b0), .GCK(n_0_1));
   HA_X1 i_0_0_0 (.A(counter[1]), .B(counter[0]), .CO(n_0_0_0), .S(n_0_0_6));
   HA_X1 i_0_0_1 (.A(counter[2]), .B(n_0_0_0), .CO(n_0_0_1), .S(n_0_0_7));
   HA_X1 i_0_0_2 (.A(counter[3]), .B(n_0_0_1), .CO(n_0_0_2), .S(n_0_0_8));
   HA_X1 i_0_0_3 (.A(counter[4]), .B(n_0_0_2), .CO(n_0_0_3), .S(n_0_0_9));
   HA_X1 i_0_0_4 (.A(counter[5]), .B(n_0_0_3), .CO(n_0_0_4), .S(n_0_0_10));
   HA_X1 i_0_0_5 (.A(counter[6]), .B(n_0_0_4), .CO(n_0_0_5), .S(n_0_0_11));
   MUX2_X1 i_0_0_6 (.A(b[1]), .B(Q[1]), .S(n_0_0_87), .Z(n_0_258));
   MUX2_X1 i_0_0_7 (.A(b[2]), .B(Q[2]), .S(n_0_0_87), .Z(n_0_259));
   MUX2_X1 i_0_0_8 (.A(b[3]), .B(Q[3]), .S(n_0_0_87), .Z(n_0_260));
   MUX2_X1 i_0_0_9 (.A(b[4]), .B(Q[4]), .S(n_0_0_87), .Z(n_0_261));
   MUX2_X1 i_0_0_10 (.A(b[5]), .B(Q[5]), .S(n_0_0_87), .Z(n_0_262));
   MUX2_X1 i_0_0_11 (.A(b[6]), .B(Q[6]), .S(n_0_0_87), .Z(n_0_263));
   MUX2_X1 i_0_0_12 (.A(b[7]), .B(Q[7]), .S(n_0_0_87), .Z(n_0_264));
   MUX2_X1 i_0_0_13 (.A(b[8]), .B(Q[8]), .S(n_0_0_87), .Z(n_0_265));
   MUX2_X1 i_0_0_14 (.A(b[9]), .B(Q[9]), .S(n_0_0_87), .Z(n_0_266));
   MUX2_X1 i_0_0_15 (.A(b[10]), .B(Q[10]), .S(n_0_0_87), .Z(n_0_267));
   MUX2_X1 i_0_0_16 (.A(b[11]), .B(Q[11]), .S(n_0_0_87), .Z(n_0_268));
   MUX2_X1 i_0_0_17 (.A(b[12]), .B(Q[12]), .S(n_0_0_87), .Z(n_0_269));
   MUX2_X1 i_0_0_18 (.A(b[13]), .B(Q[13]), .S(n_0_0_87), .Z(n_0_270));
   MUX2_X1 i_0_0_19 (.A(b[14]), .B(Q[14]), .S(n_0_0_87), .Z(n_0_271));
   MUX2_X1 i_0_0_20 (.A(b[15]), .B(Q[15]), .S(n_0_0_87), .Z(n_0_272));
   MUX2_X1 i_0_0_21 (.A(b[16]), .B(Q[16]), .S(n_0_0_87), .Z(n_0_273));
   MUX2_X1 i_0_0_22 (.A(b[17]), .B(Q[17]), .S(n_0_0_87), .Z(n_0_274));
   MUX2_X1 i_0_0_23 (.A(b[18]), .B(Q[18]), .S(n_0_0_87), .Z(n_0_275));
   MUX2_X1 i_0_0_24 (.A(b[19]), .B(Q[19]), .S(n_0_0_87), .Z(n_0_276));
   MUX2_X1 i_0_0_25 (.A(b[20]), .B(Q[20]), .S(n_0_0_87), .Z(n_0_277));
   MUX2_X1 i_0_0_26 (.A(b[21]), .B(Q[21]), .S(n_0_0_87), .Z(n_0_278));
   MUX2_X1 i_0_0_27 (.A(b[22]), .B(Q[22]), .S(n_0_0_87), .Z(n_0_279));
   MUX2_X1 i_0_0_28 (.A(b[23]), .B(Q[23]), .S(n_0_0_87), .Z(n_0_280));
   MUX2_X1 i_0_0_29 (.A(b[24]), .B(Q[24]), .S(n_0_0_87), .Z(n_0_281));
   MUX2_X1 i_0_0_30 (.A(b[25]), .B(Q[25]), .S(n_0_0_87), .Z(n_0_282));
   MUX2_X1 i_0_0_31 (.A(b[26]), .B(Q[26]), .S(n_0_0_87), .Z(n_0_283));
   MUX2_X1 i_0_0_32 (.A(b[27]), .B(Q[27]), .S(n_0_0_87), .Z(n_0_284));
   MUX2_X1 i_0_0_33 (.A(b[28]), .B(Q[28]), .S(n_0_0_87), .Z(n_0_285));
   MUX2_X1 i_0_0_34 (.A(b[29]), .B(Q[29]), .S(n_0_0_87), .Z(n_0_286));
   MUX2_X1 i_0_0_35 (.A(b[30]), .B(Q[30]), .S(n_0_0_87), .Z(n_0_287));
   MUX2_X1 i_0_0_36 (.A(b[31]), .B(Q[30]), .S(n_0_0_87), .Z(n_0_288));
   MUX2_X1 i_0_0_37 (.A(a[1]), .B(B[1]), .S(n_0_0_87), .Z(n_0_196));
   MUX2_X1 i_0_0_38 (.A(a[2]), .B(B[2]), .S(n_0_0_87), .Z(n_0_197));
   MUX2_X1 i_0_0_39 (.A(a[3]), .B(B[3]), .S(n_0_0_87), .Z(n_0_198));
   MUX2_X1 i_0_0_40 (.A(a[4]), .B(B[4]), .S(n_0_0_87), .Z(n_0_199));
   MUX2_X1 i_0_0_41 (.A(a[5]), .B(B[5]), .S(n_0_0_87), .Z(n_0_200));
   MUX2_X1 i_0_0_42 (.A(a[6]), .B(B[6]), .S(n_0_0_87), .Z(n_0_201));
   MUX2_X1 i_0_0_43 (.A(a[7]), .B(B[7]), .S(n_0_0_87), .Z(n_0_202));
   MUX2_X1 i_0_0_44 (.A(a[8]), .B(B[8]), .S(n_0_0_87), .Z(n_0_203));
   MUX2_X1 i_0_0_45 (.A(a[9]), .B(B[9]), .S(n_0_0_87), .Z(n_0_204));
   MUX2_X1 i_0_0_46 (.A(a[10]), .B(B[10]), .S(n_0_0_87), .Z(n_0_205));
   MUX2_X1 i_0_0_47 (.A(a[11]), .B(B[11]), .S(n_0_0_87), .Z(n_0_206));
   MUX2_X1 i_0_0_48 (.A(a[12]), .B(B[12]), .S(n_0_0_87), .Z(n_0_207));
   MUX2_X1 i_0_0_49 (.A(a[13]), .B(B[13]), .S(n_0_0_87), .Z(n_0_208));
   MUX2_X1 i_0_0_50 (.A(a[14]), .B(B[14]), .S(n_0_0_87), .Z(n_0_209));
   MUX2_X1 i_0_0_51 (.A(a[15]), .B(B[15]), .S(n_0_0_87), .Z(n_0_210));
   MUX2_X1 i_0_0_52 (.A(a[16]), .B(B[16]), .S(n_0_0_87), .Z(n_0_211));
   MUX2_X1 i_0_0_53 (.A(a[17]), .B(B[17]), .S(n_0_0_87), .Z(n_0_212));
   MUX2_X1 i_0_0_54 (.A(a[18]), .B(B[18]), .S(n_0_0_87), .Z(n_0_213));
   MUX2_X1 i_0_0_55 (.A(a[19]), .B(B[19]), .S(n_0_0_87), .Z(n_0_214));
   MUX2_X1 i_0_0_56 (.A(a[20]), .B(B[20]), .S(n_0_0_87), .Z(n_0_215));
   MUX2_X1 i_0_0_57 (.A(a[21]), .B(B[21]), .S(n_0_0_87), .Z(n_0_216));
   MUX2_X1 i_0_0_58 (.A(a[22]), .B(B[22]), .S(n_0_0_87), .Z(n_0_217));
   MUX2_X1 i_0_0_59 (.A(a[23]), .B(B[23]), .S(n_0_0_87), .Z(n_0_218));
   MUX2_X1 i_0_0_60 (.A(a[24]), .B(B[24]), .S(n_0_0_87), .Z(n_0_219));
   MUX2_X1 i_0_0_61 (.A(a[25]), .B(B[25]), .S(n_0_0_87), .Z(n_0_220));
   MUX2_X1 i_0_0_62 (.A(a[26]), .B(B[26]), .S(n_0_0_87), .Z(n_0_221));
   MUX2_X1 i_0_0_63 (.A(a[27]), .B(B[27]), .S(n_0_0_87), .Z(n_0_222));
   MUX2_X1 i_0_0_64 (.A(a[28]), .B(B[28]), .S(n_0_0_87), .Z(n_0_223));
   MUX2_X1 i_0_0_65 (.A(a[29]), .B(B[29]), .S(n_0_0_87), .Z(n_0_224));
   MUX2_X1 i_0_0_66 (.A(a[30]), .B(B[30]), .S(n_0_0_87), .Z(n_0_225));
   OAI21_X1 i_0_0_67 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_54), .ZN(n_0_226));
   OAI21_X1 i_0_0_68 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_55), .ZN(n_0_227));
   OAI21_X1 i_0_0_69 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_56), .ZN(n_0_228));
   OAI21_X1 i_0_0_70 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_57), .ZN(n_0_229));
   OAI21_X1 i_0_0_71 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_58), .ZN(n_0_230));
   OAI21_X1 i_0_0_72 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_59), .ZN(n_0_231));
   OAI21_X1 i_0_0_73 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_60), .ZN(n_0_232));
   OAI21_X1 i_0_0_74 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_61), .ZN(n_0_233));
   OAI21_X1 i_0_0_75 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_62), .ZN(n_0_234));
   OAI21_X1 i_0_0_76 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_63), .ZN(n_0_235));
   OAI21_X1 i_0_0_77 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_64), .ZN(n_0_236));
   OAI21_X1 i_0_0_78 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_65), .ZN(n_0_237));
   OAI21_X1 i_0_0_79 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_66), .ZN(n_0_238));
   OAI21_X1 i_0_0_80 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_67), .ZN(n_0_239));
   OAI21_X1 i_0_0_81 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_68), .ZN(n_0_240));
   OAI21_X1 i_0_0_82 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_69), .ZN(n_0_241));
   OAI21_X1 i_0_0_83 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_70), .ZN(n_0_242));
   OAI21_X1 i_0_0_84 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_71), .ZN(n_0_243));
   OAI21_X1 i_0_0_85 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_72), .ZN(n_0_244));
   OAI21_X1 i_0_0_86 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_73), .ZN(n_0_245));
   OAI21_X1 i_0_0_87 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_74), .ZN(n_0_246));
   OAI21_X1 i_0_0_88 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_75), .ZN(n_0_247));
   OAI21_X1 i_0_0_89 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_76), .ZN(n_0_248));
   OAI21_X1 i_0_0_90 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_77), .ZN(n_0_249));
   OAI21_X1 i_0_0_91 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_78), .ZN(n_0_250));
   OAI21_X1 i_0_0_92 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_79), .ZN(n_0_251));
   OAI21_X1 i_0_0_93 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_80), .ZN(n_0_252));
   OAI21_X1 i_0_0_94 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_81), .ZN(n_0_253));
   OAI21_X1 i_0_0_95 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_82), .ZN(n_0_254));
   OAI21_X1 i_0_0_96 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_83), .ZN(n_0_255));
   OAI21_X1 i_0_0_97 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_84), .ZN(n_0_256));
   OAI21_X1 i_0_0_98 (.A(n_0_0_44), .B1(n_0_0_47), .B2(n_0_0_85), .ZN(n_0_257));
   AND2_X1 i_0_0_99 (.A1(n_0_0_87), .A2(Accumulator[0]), .ZN(n_0_67));
   AND2_X1 i_0_0_100 (.A1(n_0_0_87), .A2(Accumulator[1]), .ZN(n_0_68));
   AND2_X1 i_0_0_101 (.A1(n_0_0_87), .A2(Accumulator[2]), .ZN(n_0_69));
   AND2_X1 i_0_0_102 (.A1(n_0_0_87), .A2(Accumulator[3]), .ZN(n_0_70));
   AND2_X1 i_0_0_103 (.A1(n_0_0_87), .A2(Accumulator[4]), .ZN(n_0_71));
   AND2_X1 i_0_0_104 (.A1(n_0_0_87), .A2(Accumulator[5]), .ZN(n_0_72));
   AND2_X1 i_0_0_105 (.A1(n_0_0_87), .A2(Accumulator[6]), .ZN(n_0_73));
   AND2_X1 i_0_0_106 (.A1(n_0_0_87), .A2(Accumulator[7]), .ZN(n_0_74));
   AND2_X1 i_0_0_107 (.A1(n_0_0_87), .A2(Accumulator[8]), .ZN(n_0_75));
   AND2_X1 i_0_0_108 (.A1(n_0_0_87), .A2(Accumulator[9]), .ZN(n_0_76));
   AND2_X1 i_0_0_109 (.A1(n_0_0_87), .A2(Accumulator[10]), .ZN(n_0_77));
   AND2_X1 i_0_0_110 (.A1(n_0_0_87), .A2(Accumulator[11]), .ZN(n_0_78));
   AND2_X1 i_0_0_111 (.A1(n_0_0_87), .A2(Accumulator[12]), .ZN(n_0_79));
   AND2_X1 i_0_0_112 (.A1(n_0_0_87), .A2(Accumulator[13]), .ZN(n_0_80));
   AND2_X1 i_0_0_113 (.A1(n_0_0_87), .A2(Accumulator[14]), .ZN(n_0_81));
   AND2_X1 i_0_0_114 (.A1(n_0_0_87), .A2(Accumulator[15]), .ZN(n_0_82));
   AND2_X1 i_0_0_115 (.A1(n_0_0_87), .A2(Accumulator[16]), .ZN(n_0_83));
   AND2_X1 i_0_0_116 (.A1(n_0_0_87), .A2(Accumulator[17]), .ZN(n_0_84));
   AND2_X1 i_0_0_117 (.A1(n_0_0_87), .A2(Accumulator[18]), .ZN(n_0_85));
   AND2_X1 i_0_0_118 (.A1(n_0_0_87), .A2(Accumulator[19]), .ZN(n_0_86));
   AND2_X1 i_0_0_119 (.A1(n_0_0_87), .A2(Accumulator[20]), .ZN(n_0_87));
   AND2_X1 i_0_0_120 (.A1(n_0_0_87), .A2(Accumulator[21]), .ZN(n_0_88));
   AND2_X1 i_0_0_121 (.A1(n_0_0_87), .A2(Accumulator[22]), .ZN(n_0_89));
   AND2_X1 i_0_0_122 (.A1(n_0_0_87), .A2(Accumulator[23]), .ZN(n_0_90));
   AND2_X1 i_0_0_123 (.A1(n_0_0_87), .A2(Accumulator[24]), .ZN(n_0_91));
   AND2_X1 i_0_0_124 (.A1(n_0_0_87), .A2(Accumulator[25]), .ZN(n_0_92));
   AND2_X1 i_0_0_125 (.A1(n_0_0_87), .A2(Accumulator[26]), .ZN(n_0_93));
   AND2_X1 i_0_0_126 (.A1(n_0_0_87), .A2(Accumulator[27]), .ZN(n_0_94));
   AND2_X1 i_0_0_127 (.A1(n_0_0_87), .A2(Accumulator[28]), .ZN(n_0_95));
   AND2_X1 i_0_0_128 (.A1(n_0_0_87), .A2(Accumulator[29]), .ZN(n_0_96));
   AND2_X1 i_0_0_129 (.A1(n_0_0_87), .A2(Accumulator[30]), .ZN(n_0_97));
   AND2_X1 i_0_0_130 (.A1(n_0_0_87), .A2(Accumulator[31]), .ZN(n_0_98));
   AND2_X1 i_0_0_131 (.A1(n_0_0_87), .A2(Accumulator[32]), .ZN(n_0_99));
   AND2_X1 i_0_0_132 (.A1(n_0_0_87), .A2(Accumulator[33]), .ZN(n_0_100));
   AND2_X1 i_0_0_133 (.A1(n_0_0_87), .A2(Accumulator[34]), .ZN(n_0_101));
   AND2_X1 i_0_0_134 (.A1(n_0_0_87), .A2(Accumulator[35]), .ZN(n_0_102));
   AND2_X1 i_0_0_135 (.A1(n_0_0_87), .A2(Accumulator[36]), .ZN(n_0_103));
   AND2_X1 i_0_0_136 (.A1(n_0_0_87), .A2(Accumulator[37]), .ZN(n_0_104));
   AND2_X1 i_0_0_137 (.A1(n_0_0_87), .A2(Accumulator[38]), .ZN(n_0_105));
   AND2_X1 i_0_0_138 (.A1(n_0_0_87), .A2(Accumulator[39]), .ZN(n_0_106));
   AND2_X1 i_0_0_139 (.A1(n_0_0_87), .A2(Accumulator[40]), .ZN(n_0_107));
   AND2_X1 i_0_0_140 (.A1(n_0_0_87), .A2(Accumulator[41]), .ZN(n_0_108));
   AND2_X1 i_0_0_141 (.A1(n_0_0_87), .A2(Accumulator[42]), .ZN(n_0_109));
   AND2_X1 i_0_0_142 (.A1(n_0_0_87), .A2(Accumulator[43]), .ZN(n_0_110));
   AND2_X1 i_0_0_143 (.A1(n_0_0_87), .A2(Accumulator[44]), .ZN(n_0_111));
   AND2_X1 i_0_0_144 (.A1(n_0_0_87), .A2(Accumulator[45]), .ZN(n_0_112));
   AND2_X1 i_0_0_145 (.A1(n_0_0_87), .A2(Accumulator[46]), .ZN(n_0_113));
   AND2_X1 i_0_0_146 (.A1(n_0_0_87), .A2(Accumulator[47]), .ZN(n_0_114));
   AND2_X1 i_0_0_147 (.A1(n_0_0_87), .A2(Accumulator[48]), .ZN(n_0_115));
   AND2_X1 i_0_0_148 (.A1(n_0_0_87), .A2(Accumulator[49]), .ZN(n_0_116));
   AND2_X1 i_0_0_149 (.A1(n_0_0_87), .A2(Accumulator[50]), .ZN(n_0_117));
   AND2_X1 i_0_0_150 (.A1(n_0_0_87), .A2(Accumulator[51]), .ZN(n_0_118));
   AND2_X1 i_0_0_151 (.A1(n_0_0_87), .A2(Accumulator[52]), .ZN(n_0_119));
   AND2_X1 i_0_0_152 (.A1(n_0_0_87), .A2(Accumulator[53]), .ZN(n_0_120));
   AND2_X1 i_0_0_153 (.A1(n_0_0_87), .A2(Accumulator[54]), .ZN(n_0_121));
   AND2_X1 i_0_0_154 (.A1(n_0_0_87), .A2(Accumulator[55]), .ZN(n_0_122));
   AND2_X1 i_0_0_155 (.A1(n_0_0_87), .A2(Accumulator[56]), .ZN(n_0_123));
   AND2_X1 i_0_0_156 (.A1(n_0_0_87), .A2(Accumulator[57]), .ZN(n_0_124));
   AND2_X1 i_0_0_157 (.A1(n_0_0_87), .A2(Accumulator[58]), .ZN(n_0_125));
   AND2_X1 i_0_0_158 (.A1(n_0_0_87), .A2(Accumulator[59]), .ZN(n_0_126));
   AND2_X1 i_0_0_159 (.A1(n_0_0_87), .A2(Accumulator[60]), .ZN(n_0_127));
   AND2_X1 i_0_0_160 (.A1(n_0_0_87), .A2(Accumulator[61]), .ZN(n_0_128));
   AND2_X1 i_0_0_161 (.A1(n_0_0_87), .A2(Accumulator[62]), .ZN(n_0_129));
   AND2_X1 i_0_0_162 (.A1(n_0_0_87), .A2(Accumulator[63]), .ZN(n_0_130));
   AND2_X1 i_0_0_163 (.A1(b[0]), .A2(n_0_195), .ZN(n_0_3));
   AND2_X1 i_0_0_164 (.A1(a[0]), .A2(n_0_0_47), .ZN(n_0_195));
   INV_X1 i_0_0_165 (.A(n_0_0_12), .ZN(n_0_4));
   AOI22_X1 i_0_0_166 (.A1(B[1]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[1]), 
      .ZN(n_0_0_12));
   INV_X1 i_0_0_167 (.A(n_0_0_13), .ZN(n_0_5));
   AOI22_X1 i_0_0_168 (.A1(B[2]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[2]), 
      .ZN(n_0_0_13));
   INV_X1 i_0_0_169 (.A(n_0_0_14), .ZN(n_0_6));
   AOI22_X1 i_0_0_170 (.A1(B[3]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[3]), 
      .ZN(n_0_0_14));
   INV_X1 i_0_0_171 (.A(n_0_0_15), .ZN(n_0_7));
   AOI22_X1 i_0_0_172 (.A1(B[4]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[4]), 
      .ZN(n_0_0_15));
   INV_X1 i_0_0_173 (.A(n_0_0_16), .ZN(n_0_8));
   AOI22_X1 i_0_0_174 (.A1(B[5]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[5]), 
      .ZN(n_0_0_16));
   INV_X1 i_0_0_175 (.A(n_0_0_17), .ZN(n_0_9));
   AOI22_X1 i_0_0_176 (.A1(B[6]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[6]), 
      .ZN(n_0_0_17));
   INV_X1 i_0_0_177 (.A(n_0_0_18), .ZN(n_0_10));
   AOI22_X1 i_0_0_178 (.A1(B[7]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[7]), 
      .ZN(n_0_0_18));
   INV_X1 i_0_0_179 (.A(n_0_0_19), .ZN(n_0_11));
   AOI22_X1 i_0_0_180 (.A1(B[8]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[8]), 
      .ZN(n_0_0_19));
   INV_X1 i_0_0_181 (.A(n_0_0_20), .ZN(n_0_12));
   AOI22_X1 i_0_0_182 (.A1(B[9]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[9]), 
      .ZN(n_0_0_20));
   INV_X1 i_0_0_183 (.A(n_0_0_21), .ZN(n_0_13));
   AOI22_X1 i_0_0_184 (.A1(B[10]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[10]), 
      .ZN(n_0_0_21));
   INV_X1 i_0_0_185 (.A(n_0_0_22), .ZN(n_0_14));
   AOI22_X1 i_0_0_186 (.A1(B[11]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[11]), 
      .ZN(n_0_0_22));
   INV_X1 i_0_0_187 (.A(n_0_0_23), .ZN(n_0_15));
   AOI22_X1 i_0_0_188 (.A1(B[12]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[12]), 
      .ZN(n_0_0_23));
   INV_X1 i_0_0_189 (.A(n_0_0_24), .ZN(n_0_16));
   AOI22_X1 i_0_0_190 (.A1(B[13]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[13]), 
      .ZN(n_0_0_24));
   INV_X1 i_0_0_191 (.A(n_0_0_25), .ZN(n_0_17));
   AOI22_X1 i_0_0_192 (.A1(B[14]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[14]), 
      .ZN(n_0_0_25));
   INV_X1 i_0_0_193 (.A(n_0_0_26), .ZN(n_0_18));
   AOI22_X1 i_0_0_194 (.A1(B[15]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[15]), 
      .ZN(n_0_0_26));
   INV_X1 i_0_0_195 (.A(n_0_0_27), .ZN(n_0_19));
   AOI22_X1 i_0_0_196 (.A1(B[16]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[16]), 
      .ZN(n_0_0_27));
   INV_X1 i_0_0_197 (.A(n_0_0_28), .ZN(n_0_20));
   AOI22_X1 i_0_0_198 (.A1(B[17]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[17]), 
      .ZN(n_0_0_28));
   INV_X1 i_0_0_199 (.A(n_0_0_29), .ZN(n_0_21));
   AOI22_X1 i_0_0_200 (.A1(B[18]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[18]), 
      .ZN(n_0_0_29));
   INV_X1 i_0_0_201 (.A(n_0_0_30), .ZN(n_0_22));
   AOI22_X1 i_0_0_202 (.A1(B[19]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[19]), 
      .ZN(n_0_0_30));
   INV_X1 i_0_0_203 (.A(n_0_0_31), .ZN(n_0_23));
   AOI22_X1 i_0_0_204 (.A1(B[20]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[20]), 
      .ZN(n_0_0_31));
   INV_X1 i_0_0_205 (.A(n_0_0_32), .ZN(n_0_24));
   AOI22_X1 i_0_0_206 (.A1(B[21]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[21]), 
      .ZN(n_0_0_32));
   INV_X1 i_0_0_207 (.A(n_0_0_33), .ZN(n_0_25));
   AOI22_X1 i_0_0_208 (.A1(B[22]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[22]), 
      .ZN(n_0_0_33));
   INV_X1 i_0_0_209 (.A(n_0_0_34), .ZN(n_0_26));
   AOI22_X1 i_0_0_210 (.A1(B[23]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[23]), 
      .ZN(n_0_0_34));
   INV_X1 i_0_0_211 (.A(n_0_0_35), .ZN(n_0_27));
   AOI22_X1 i_0_0_212 (.A1(B[24]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[24]), 
      .ZN(n_0_0_35));
   INV_X1 i_0_0_213 (.A(n_0_0_36), .ZN(n_0_28));
   AOI22_X1 i_0_0_214 (.A1(B[25]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[25]), 
      .ZN(n_0_0_36));
   INV_X1 i_0_0_215 (.A(n_0_0_37), .ZN(n_0_29));
   AOI22_X1 i_0_0_216 (.A1(B[26]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[26]), 
      .ZN(n_0_0_37));
   INV_X1 i_0_0_217 (.A(n_0_0_38), .ZN(n_0_30));
   AOI22_X1 i_0_0_218 (.A1(B[27]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[27]), 
      .ZN(n_0_0_38));
   INV_X1 i_0_0_219 (.A(n_0_0_39), .ZN(n_0_31));
   AOI22_X1 i_0_0_220 (.A1(B[28]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[28]), 
      .ZN(n_0_0_39));
   INV_X1 i_0_0_221 (.A(n_0_0_40), .ZN(n_0_32));
   AOI22_X1 i_0_0_222 (.A1(B[29]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[29]), 
      .ZN(n_0_0_40));
   INV_X1 i_0_0_223 (.A(n_0_0_41), .ZN(n_0_33));
   AOI22_X1 i_0_0_224 (.A1(B[30]), .A2(n_0_0_46), .B1(n_0_0_42), .B2(a[30]), 
      .ZN(n_0_0_41));
   OAI21_X1 i_0_0_225 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_54), .ZN(n_0_34));
   OAI21_X1 i_0_0_226 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_55), .ZN(n_0_35));
   OAI21_X1 i_0_0_227 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_56), .ZN(n_0_36));
   OAI21_X1 i_0_0_228 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_57), .ZN(n_0_37));
   OAI21_X1 i_0_0_229 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_58), .ZN(n_0_38));
   OAI21_X1 i_0_0_230 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_59), .ZN(n_0_39));
   OAI21_X1 i_0_0_231 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_60), .ZN(n_0_40));
   OAI21_X1 i_0_0_232 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_61), .ZN(n_0_41));
   OAI21_X1 i_0_0_233 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_62), .ZN(n_0_42));
   OAI21_X1 i_0_0_234 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_63), .ZN(n_0_43));
   OAI21_X1 i_0_0_235 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_64), .ZN(n_0_44));
   OAI21_X1 i_0_0_236 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_65), .ZN(n_0_45));
   OAI21_X1 i_0_0_237 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_66), .ZN(n_0_46));
   OAI21_X1 i_0_0_238 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_67), .ZN(n_0_47));
   OAI21_X1 i_0_0_239 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_68), .ZN(n_0_48));
   OAI21_X1 i_0_0_240 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_69), .ZN(n_0_49));
   OAI21_X1 i_0_0_241 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_70), .ZN(n_0_50));
   OAI21_X1 i_0_0_242 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_71), .ZN(n_0_51));
   OAI21_X1 i_0_0_243 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_72), .ZN(n_0_52));
   OAI21_X1 i_0_0_244 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_73), .ZN(n_0_53));
   OAI21_X1 i_0_0_245 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_74), .ZN(n_0_54));
   OAI21_X1 i_0_0_246 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_75), .ZN(n_0_55));
   OAI21_X1 i_0_0_247 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_76), .ZN(n_0_56));
   OAI21_X1 i_0_0_248 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_77), .ZN(n_0_57));
   OAI21_X1 i_0_0_249 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_78), .ZN(n_0_58));
   OAI21_X1 i_0_0_250 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_79), .ZN(n_0_59));
   OAI21_X1 i_0_0_251 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_80), .ZN(n_0_60));
   OAI21_X1 i_0_0_252 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_81), .ZN(n_0_61));
   OAI21_X1 i_0_0_253 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_82), .ZN(n_0_62));
   OAI21_X1 i_0_0_254 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_83), .ZN(n_0_63));
   OAI21_X1 i_0_0_255 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_84), .ZN(n_0_64));
   OAI21_X1 i_0_0_256 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_85), .ZN(n_0_65));
   OAI21_X1 i_0_0_257 (.A(n_0_0_43), .B1(n_0_0_45), .B2(n_0_0_86), .ZN(n_0_66));
   AND2_X1 i_0_0_258 (.A1(b[0]), .A2(n_0_0_47), .ZN(n_0_0_42));
   NAND3_X1 i_0_0_259 (.A1(a[31]), .A2(b[0]), .A3(n_0_0_47), .ZN(n_0_0_43));
   NAND2_X1 i_0_0_260 (.A1(a[31]), .A2(n_0_0_47), .ZN(n_0_0_44));
   INV_X1 i_0_0_261 (.A(n_0_0_46), .ZN(n_0_0_45));
   AND2_X1 i_0_0_262 (.A1(n_0_0_87), .A2(Q[0]), .ZN(n_0_0_46));
   AND3_X1 i_0_0_263 (.A1(n_0_0_51), .A2(n_0_0_49), .A3(n_0_0_48), .ZN(n_0_0_47));
   NOR2_X1 i_0_0_264 (.A1(counter[5]), .A2(counter[4]), .ZN(n_0_0_48));
   NOR4_X1 i_0_0_265 (.A1(counter[3]), .A2(counter[2]), .A3(counter[1]), 
      .A4(counter[0]), .ZN(n_0_0_49));
   AND2_X1 i_0_0_266 (.A1(n_0_0_50), .A2(n_0_0_6), .ZN(n_0_291));
   AND2_X1 i_0_0_267 (.A1(n_0_0_50), .A2(n_0_0_7), .ZN(n_0_292));
   AND2_X1 i_0_0_268 (.A1(n_0_0_50), .A2(n_0_0_8), .ZN(n_0_293));
   AND2_X1 i_0_0_269 (.A1(n_0_0_50), .A2(n_0_0_9), .ZN(n_0_294));
   AND2_X1 i_0_0_270 (.A1(n_0_0_50), .A2(n_0_0_10), .ZN(n_0_295));
   AND2_X1 i_0_0_271 (.A1(n_0_0_50), .A2(n_0_0_11), .ZN(n_0_296));
   NOR2_X1 i_0_0_272 (.A1(n_0_2), .A2(n_0_0_53), .ZN(n_0_297));
   INV_X1 i_0_0_273 (.A(n_0_0_50), .ZN(n_0_2));
   NAND4_X1 i_0_0_274 (.A1(counter[5]), .A2(counter[4]), .A3(n_0_0_52), .A4(
      n_0_0_51), .ZN(n_0_0_50));
   NOR2_X1 i_0_0_275 (.A1(counter[7]), .A2(counter[6]), .ZN(n_0_0_51));
   AND4_X1 i_0_0_276 (.A1(counter[3]), .A2(counter[2]), .A3(counter[1]), 
      .A4(counter[0]), .ZN(n_0_0_52));
   XNOR2_X1 i_0_0_277 (.A(counter[7]), .B(n_0_0_5), .ZN(n_0_0_53));
   INV_X1 i_0_0_278 (.A(B[31]), .ZN(n_0_0_54));
   INV_X1 i_0_0_279 (.A(B[32]), .ZN(n_0_0_55));
   INV_X1 i_0_0_280 (.A(B[33]), .ZN(n_0_0_56));
   INV_X1 i_0_0_281 (.A(B[34]), .ZN(n_0_0_57));
   INV_X1 i_0_0_282 (.A(B[35]), .ZN(n_0_0_58));
   INV_X1 i_0_0_283 (.A(B[36]), .ZN(n_0_0_59));
   INV_X1 i_0_0_284 (.A(B[37]), .ZN(n_0_0_60));
   INV_X1 i_0_0_285 (.A(B[38]), .ZN(n_0_0_61));
   INV_X1 i_0_0_286 (.A(B[39]), .ZN(n_0_0_62));
   INV_X1 i_0_0_287 (.A(B[40]), .ZN(n_0_0_63));
   INV_X1 i_0_0_288 (.A(B[41]), .ZN(n_0_0_64));
   INV_X1 i_0_0_289 (.A(B[42]), .ZN(n_0_0_65));
   INV_X1 i_0_0_290 (.A(B[43]), .ZN(n_0_0_66));
   INV_X1 i_0_0_291 (.A(B[44]), .ZN(n_0_0_67));
   INV_X1 i_0_0_292 (.A(B[45]), .ZN(n_0_0_68));
   INV_X1 i_0_0_293 (.A(B[46]), .ZN(n_0_0_69));
   INV_X1 i_0_0_294 (.A(B[47]), .ZN(n_0_0_70));
   INV_X1 i_0_0_295 (.A(B[48]), .ZN(n_0_0_71));
   INV_X1 i_0_0_296 (.A(B[49]), .ZN(n_0_0_72));
   INV_X1 i_0_0_297 (.A(B[50]), .ZN(n_0_0_73));
   INV_X1 i_0_0_298 (.A(B[51]), .ZN(n_0_0_74));
   INV_X1 i_0_0_299 (.A(B[52]), .ZN(n_0_0_75));
   INV_X1 i_0_0_300 (.A(B[53]), .ZN(n_0_0_76));
   INV_X1 i_0_0_301 (.A(B[54]), .ZN(n_0_0_77));
   INV_X1 i_0_0_302 (.A(B[55]), .ZN(n_0_0_78));
   INV_X1 i_0_0_303 (.A(B[56]), .ZN(n_0_0_79));
   INV_X1 i_0_0_304 (.A(B[57]), .ZN(n_0_0_80));
   INV_X1 i_0_0_305 (.A(B[58]), .ZN(n_0_0_81));
   INV_X1 i_0_0_306 (.A(B[59]), .ZN(n_0_0_82));
   INV_X1 i_0_0_307 (.A(B[60]), .ZN(n_0_0_83));
   INV_X1 i_0_0_308 (.A(B[61]), .ZN(n_0_0_84));
   INV_X1 i_0_0_309 (.A(B[62]), .ZN(n_0_0_85));
   INV_X1 i_0_0_310 (.A(B[63]), .ZN(n_0_0_86));
   INV_X1 i_0_0_311 (.A(rst), .ZN(n_0_289));
   INV_X1 i_0_0_312 (.A(counter[0]), .ZN(n_0_290));
   INV_X1 i_0_0_313 (.A(n_0_0_47), .ZN(n_0_0_87));
endmodule
