* SPICE NETLIST
***************************************

.SUBCKT MGC_via2_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT via2_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT WELLTAP
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_3
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X2
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_4
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT INV_X1 A VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4
** N=4 EP=4 IP=7 FDC=2
X1 3 1 2 4 INV_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT NOR2_X1 A2 VDD A1 ZN VSS
** N=6 EP=5 IP=0 FDC=4
M0 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 6 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 ZN A1 6 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X4
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AOI22_X1 B2 B1 VDD A1 ZN A2 VSS
** N=10 EP=7 IP=0 FDC=8
M0 9 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN B1 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 10 A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 VSS A2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 VDD B2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 8 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 8 A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN 6
** N=8 EP=6 IP=0 FDC=6
M0 8 A1 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A1 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI21_X1 B2 B1 ZN A VSS VDD
** N=8 EP=6 IP=0 FDC=6
M0 8 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN B1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 7 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2_X1 VSS A ZN B VDD
** N=9 EP=5 IP=0 FDC=10
M0 9 A 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=155 $Y=90 $D=1
M1 VSS B 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=345 $Y=90 $D=1
M2 7 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=540 $Y=90 $D=1
M3 ZN A 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 7 B ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 6 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=155 $Y=995 $D=0
M6 VDD B 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=345 $Y=995 $D=0
M7 ZN 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=540 $Y=680 $D=0
M8 8 A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M9 VDD B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS
** N=9 EP=5 IP=0 FDC=10
M0 6 A VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 9 A Z VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 8 A 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 7 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 7 B Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X8
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_16
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT OR3_X1 A1 A2 A3 VSS VDD ZN
** N=9 EP=6 IP=0 FDC=8
M0 VSS A1 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 7 A2 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 VSS A3 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=525 $Y=90 $D=1
M3 ZN 7 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 8 A1 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M5 9 A2 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M6 VDD A3 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=525 $Y=995 $D=0
M7 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT OAI21_X1 B2 B1 ZN A VSS VDD
** N=8 EP=6 IP=0 FDC=6
M0 ZN B2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 7 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS A 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 8 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M4 ZN B1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M5 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=6
X1 3 4 1 2 5 1 AND2_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6
** N=6 EP=6 IP=9 FDC=6
X1 3 4 1 2 5 6 AND2_X1 $T=950 0 1 180 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_29
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT DFF_X1 D CK VSS VDD Q 6
** N=21 EP=6 IP=0 FDC=28
M0 VSS 10 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=160 $Y=180 $D=1
M1 18 9 VSS 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=350 $Y=300 $D=1
M2 8 7 18 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.6e-14 AS=1.26e-14 PD=8.4e-07 PS=4.6e-07 $X=540 $Y=300 $D=1
M3 19 10 8 6 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=2.6e-14 PD=8.3e-07 PS=8.4e-07 $X=735 $Y=180 $D=1
M4 VSS D 19 6 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.395e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=925 $Y=180 $D=1
M5 9 8 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=3.395e-14 PD=6.3e-07 PS=8.3e-07 $X=1115 $Y=180 $D=1
M6 VSS CK 10 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1530 $Y=255 $D=1
M7 20 8 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1720 $Y=255 $D=1
M8 11 7 20 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1910 $Y=255 $D=1
M9 21 10 11 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.1e-14 PD=4.7e-07 PS=7e-07 $X=2100 $Y=300 $D=1
M10 VSS 13 21 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.305e-14 PD=7e-07 PS=4.7e-07 $X=2295 $Y=300 $D=1
M11 13 11 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.1e-14 PD=6.3e-07 PS=7e-07 $X=2485 $Y=255 $D=1
M12 VSS 11 QN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=2825 $Y=90 $D=1
M13 Q 13 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=3015 $Y=90 $D=1
M14 VDD 10 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=160 $Y=785 $D=0
M15 14 9 VDD VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=350 $Y=1010 $D=0
M16 8 10 14 VDD PMOS_VTL L=5e-08 W=9e-08 AD=3.615e-14 AS=1.26e-14 PD=1.13e-06 PS=4.6e-07 $X=540 $Y=1010 $D=0
M17 15 7 8 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=3.615e-14 PD=1.12e-06 PS=1.13e-06 $X=735 $Y=765 $D=0
M18 VDD D 15 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.145e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=925 $Y=765 $D=0
M19 9 8 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=5.145e-14 PD=9.9e-07 PS=1.12e-06 $X=1115 $Y=870 $D=0
M20 VDD CK 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1530 $Y=870 $D=0
M21 16 8 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1720 $Y=870 $D=0
M22 11 10 16 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1910 $Y=870 $D=0
M23 17 7 11 VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.835e-14 PD=4.7e-07 PS=9.1e-07 $X=2100 $Y=1095 $D=0
M24 VDD 13 17 VDD PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.305e-14 PD=9.1e-07 PS=4.7e-07 $X=2295 $Y=1095 $D=0
M25 13 11 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=2.835e-14 PD=8.4e-07 PS=9.1e-07 $X=2485 $Y=870 $D=0
M26 VDD 11 QN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=2825 $Y=680 $D=0
M27 Q 13 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3015 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_34 1 2 3 4 5 6
** N=6 EP=6 IP=9 FDC=28
X1 3 4 1 2 5 6 DFF_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT NAND2_X1 A2 VSS A1 ZN VDD
** N=6 EP=5 IP=0 FDC=4
M0 6 A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN A1 6 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_35
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X16
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_37
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT via1_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_38
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4
** N=4 EP=4 IP=7 FDC=2
X0 1 2 3 4 INV_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT OR2_X1 A1 A2 VSS VDD ZN
** N=7 EP=5 IP=0 FDC=6
M0 6 A1 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A1 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_40
** N=2 EP=0 IP=5 FDC=0
.ENDS
***************************************
.SUBCKT ICV_41
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_42
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_43
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_44
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_45
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_46
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_47
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AOI222_X1 C2 C1 VDD B1 B2 A2 VSS A1 ZN
** N=14 EP=9 IP=0 FDC=12
M0 12 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN C1 12 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=1.2035e-13 AS=5.81e-14 PD=1.41e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 13 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=1.2035e-13 PD=1.11e-06 PS=1.41e-06 $X=675 $Y=90 $D=1
M3 VSS B2 13 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=865 $Y=90 $D=1
M4 14 A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1055 $Y=90 $D=1
M5 ZN A1 14 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1245 $Y=90 $D=1
M6 10 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M7 VDD C1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M8 10 B1 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=675 $Y=680 $D=0
M9 11 B2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=865 $Y=680 $D=0
M10 ZN A2 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1055 $Y=680 $D=0
M11 11 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1245 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_48
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_49
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_50
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI221_X1 B2 B1 VSS A C2 VDD C1 ZN
** N=12 EP=8 IP=0 FDC=10
M0 VSS B2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 9 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 10 A 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN C2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 10 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 11 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 ZN B1 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 12 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 ZN C1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_51
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT OAI22_X1 B2 B1 VSS ZN A1 A2 VDD
** N=10 EP=7 IP=0 FDC=8
M0 VSS B2 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 8 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 8 A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 9 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 ZN B1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 10 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 VDD A2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_52
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_53 1 2 3 4
** N=4 EP=4 IP=7 FDC=2
X0 1 2 3 4 INV_X1 $T=380 0 0 0 $X=265 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_54
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_55 1 2 3 4 5 6 7 8 9 10 11 12
** N=12 EP=12 IP=14 FDC=16
X0 1 2 3 4 5 6 7 AOI22_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 8 9 3 10 11 12 7 AOI22_X1 $T=950 0 0 0 $X=835 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_56
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_57 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=4
X1 3 1 4 5 2 NAND2_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT FILLCELL_X32
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_58 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=8
X1 3 4 2 5 6 7 1 AOI22_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_59
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_60
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_61
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_62
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_63
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT OAI211_X1 C2 C1 A VDD B ZN VSS
** N=10 EP=7 IP=0 FDC=8
M0 ZN C2 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 8 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 10 A 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS B 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 9 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN C1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 ZN B VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI221_X1 B2 B1 VDD A C2 VSS C1 ZN
** N=12 EP=8 IP=0 FDC=10
M0 11 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN B1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 12 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN C1 12 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VDD B2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 9 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 10 A 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 ZN C2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 10 C1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_64 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=11 FDC=10
X0 1 2 3 4 5 6 OAI21_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 7 5 8 9 6 NAND2_X1 $T=1330 0 1 180 $X=645 $Y=-115
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_65
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_66
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_67
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_68
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT NAND4_X1 A4 VSS A3 A2 A1 ZN VDD
** N=10 EP=7 IP=0 FDC=8
M0 8 A4 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 9 A3 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 10 A2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN A4 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 VDD A3 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_69
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_70
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT NOR3_X1 A3 VDD A2 A1 VSS ZN
** N=8 EP=6 IP=0 FDC=6
M0 ZN A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 8 A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_71
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_72 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=56
X0 1 2 3 4 5 3 DFF_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 6 7 3 4 8 3 DFF_X1 $T=3230 0 0 0 $X=3115 $Y=-115
.ENDS
***************************************
.SUBCKT NOR4_X1 A4 VDD A3 A2 A1 ZN VSS
** N=10 EP=7 IP=0 FDC=8
M0 ZN A4 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A3 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 8 A4 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 9 A3 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 10 A2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 ZN A1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI211_X1 C2 C1 B VSS A ZN VDD
** N=10 EP=7 IP=0 FDC=8
M0 10 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN C1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS B ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 ZN C2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 8 C1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 9 B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3_X1 A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
M0 7 A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 8 A2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 VDD A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_73 1 2 3 4
** N=4 EP=4 IP=7 FDC=2
X0 1 2 3 4 INV_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_AUTO_NDR_MGC_CLK_NDR_1.0w2.0s_via2_single_MA_north
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND3_X1 A1 A2 A3 VSS VDD ZN
** N=9 EP=6 IP=0 FDC=8
M0 8 A1 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 9 A2 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 VSS A3 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=525 $Y=90 $D=1
M3 ZN 7 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 VDD A1 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M5 7 A2 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M6 VDD A3 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=525 $Y=995 $D=0
M7 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR2_X2 A1 ZN A2 VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 6 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN A1 6 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 7 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR3_X2 A1 ZN A2 A3 VSS VDD
** N=10 EP=6 IP=0 FDC=12
M0 ZN A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=945 $Y=90 $D=1
M5 VSS A3 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1135 $Y=90 $D=1
M6 7 A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M7 8 A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M8 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M9 9 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
M10 10 A2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=945 $Y=680 $D=0
M11 VDD A3 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1135 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUF_X1 A VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS A 5 VSS NMOS_VTL L=5e-08 W=9.5e-08 AD=2.03e-14 AS=9.975e-15 PD=6.7e-07 PS=4e-07 $X=165 $Y=160 $D=1
M1 Z 5 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.03e-14 PD=6e-07 PS=6.7e-07 $X=355 $Y=160 $D=1
M2 VDD A 5 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=165 $Y=995 $D=0
M3 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=355 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI21_X2 A VSS B1 ZN B2 VDD
** N=9 EP=6 IP=0 FDC=12
M0 VSS A 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 7 A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN B2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN B1 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 7 B2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1095 $Y=90 $D=1
M6 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M7 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M8 8 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M9 ZN B1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M10 9 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
M11 VDD B2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1095 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT HA_X1 S B A VSS VDD CO
** N=12 EP=6 IP=0 FDC=16
M0 11 B VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 S A 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 8 S VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.48e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 8 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.48e-14 PD=7e-07 PS=1.12e-06 $X=760 $Y=90 $D=1
M4 VSS A 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=950 $Y=90 $D=1
M5 12 A 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1320 $Y=90 $D=1
M6 VSS B 12 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=1510 $Y=90 $D=1
M7 CO 9 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1700 $Y=90 $D=1
M8 S B 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 7 A S VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 VDD 8 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.7725e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 10 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.7725e-14 PD=9.1e-07 PS=1.55e-06 $X=760 $Y=870 $D=0
M12 8 A 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=950 $Y=870 $D=0
M13 9 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1320 $Y=870 $D=0
M14 VDD B 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=1510 $Y=870 $D=0
M15 CO 9 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1700 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI222_X2 C1 VDD C2 B1 B2 A1 A2 ZN VSS
** N=17 EP=9 IP=0 FDC=24
M0 13 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN C1 13 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 14 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS C2 14 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 15 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 ZN B1 15 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1095 $Y=90 $D=1
M6 16 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1285 $Y=90 $D=1
M7 VSS B2 16 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1475 $Y=90 $D=1
M8 ZN A1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=1850 $Y=90 $D=1
M9 17 A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2040 $Y=90 $D=1
M10 VSS A2 17 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2230 $Y=90 $D=1
M11 11 A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=2420 $Y=90 $D=1
M12 VDD C2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M13 10 C1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M14 VDD C1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M15 10 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M16 12 B2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
M17 10 B1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1095 $Y=680 $D=0
M18 12 B1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1285 $Y=680 $D=0
M19 10 B2 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1475 $Y=680 $D=0
M20 ZN A1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=1850 $Y=680 $D=0
M21 12 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2040 $Y=680 $D=0
M22 ZN A2 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2230 $Y=680 $D=0
M23 12 A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=2420 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FA_X1 CO CI B A VDD VSS
** N=19 EP=6 IP=0 FDC=28
M0 VSS 7 CO VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 17 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=360 $Y=215 $D=1
M2 7 A 17 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=550 $Y=215 $D=1
M3 8 CI 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07 $X=740 $Y=215 $D=1
M4 VSS A 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=935 $Y=215 $D=1
M5 8 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1125 $Y=215 $D=1
M6 10 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1465 $Y=90 $D=1
M7 VSS CI 10 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1655 $Y=90 $D=1
M8 10 A VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1845 $Y=90 $D=1
M9 12 7 10 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07 $X=2035 $Y=90 $D=1
M10 18 CI 12 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07 $X=2235 $Y=90 $D=1
M11 19 B 18 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2425 $Y=90 $D=1
M12 VSS A 19 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=2615 $Y=90 $D=1
M13 S 12 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M14 VDD 7 CO VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M15 14 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=360 $Y=870 $D=0
M16 7 A 14 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=550 $Y=870 $D=0
M17 9 CI 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06 PS=9.1e-07 $X=740 $Y=870 $D=0
M18 VDD A 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06 $X=935 $Y=945 $D=0
M19 9 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1125 $Y=945 $D=0
M20 11 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1465 $Y=995 $D=0
M21 VDD CI 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1655 $Y=995 $D=0
M22 11 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1845 $Y=995 $D=0
M23 12 7 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07 $X=2035 $Y=995 $D=0
M24 15 CI 12 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07 $X=2235 $Y=995 $D=0
M25 16 B 15 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2425 $Y=995 $D=0
M26 VDD A 16 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2615 $Y=995 $D=0
M27 S 12 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI33_X1 B3 B2 B1 VSS A1 A2 A3 ZN VDD
** N=14 EP=9 IP=0 FDC=12
M0 10 B3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS B2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 10 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 ZN A1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 10 A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 ZN A3 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1110 $Y=90 $D=1
M6 11 B3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M7 12 B2 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M8 ZN B1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M9 13 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M10 14 A2 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
M11 VDD A3 14 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1110 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT CLKGATETST_X1 SE E CK VDD VSS GCK 7
** N=19 EP=7 IP=0 FDC=24
M0 8 SE VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=205 $D=1
M1 VSS E 8 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.94e-14 PD=8.3e-07 PS=7e-07 $X=335 $Y=205 $D=1
M2 17 8 VSS 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=8.3e-07 $X=525 $Y=140 $D=1
M3 9 12 17 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=2.915e-14 AS=3.85e-14 PD=9.1e-07 PS=8.3e-07 $X=715 $Y=140 $D=1
M4 18 10 9 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.915e-14 PD=4.6e-07 PS=9.1e-07 $X=945 $Y=300 $D=1
M5 VSS 11 18 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.26e-14 PD=7e-07 PS=4.6e-07 $X=1135 $Y=300 $D=1
M6 10 12 VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.1e-14 PD=6.3e-07 PS=7e-07 $X=1325 $Y=180 $D=1
M7 VSS 9 11 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1665 $Y=315 $D=1
M8 12 CK VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1855 $Y=315 $D=1
M9 19 CK 13 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=2240 $Y=295 $D=1
M10 VSS 9 19 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.835e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2430 $Y=295 $D=1
M11 GCK 13 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.835e-14 PD=6e-07 PS=7e-07 $X=2620 $Y=310 $D=1
M12 14 SE 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=890 $D=0
M13 VDD E 14 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=4.41e-14 PD=1.12e-06 PS=9.1e-07 $X=335 $Y=890 $D=0
M14 15 8 VDD VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=525 $Y=890 $D=0
M15 9 10 15 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=3.93e-14 AS=5.88e-14 PD=1.2e-06 PS=1.12e-06 $X=715 $Y=890 $D=0
M16 16 12 9 VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.93e-14 PD=4.6e-07 PS=1.2e-06 $X=945 $Y=990 $D=0
M17 VDD 11 16 VDD PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.26e-14 PD=9.1e-07 PS=4.6e-07 $X=1135 $Y=990 $D=0
M18 10 12 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=2.835e-14 PD=8.4e-07 PS=9.1e-07 $X=1325 $Y=990 $D=0
M19 VDD 9 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1665 $Y=870 $D=0
M20 12 CK VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1855 $Y=870 $D=0
M21 13 CK VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=2240 $Y=870 $D=0
M22 VDD 9 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2430 $Y=870 $D=0
M23 GCK 13 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2620 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT fp_adder_buff
** N=1265 EP=0 IP=22316 FDC=9712
M0 271 504 506 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=3045 $Y=45515 $D=1
M1 23 506 271 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=3235 $Y=45515 $D=1
M2 271 506 23 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=3425 $Y=45515 $D=1
M3 23 506 271 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=3615 $Y=45515 $D=1
M4 1256 169 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=19980 $Y=34095 $D=1
M5 151 562 1256 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=20170 $Y=34095 $D=1
M6 1257 562 151 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=20360 $Y=34095 $D=1
M7 271 169 1257 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=20550 $Y=34095 $D=1
M8 609 271 271 271 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=30240 $Y=15090 $D=1
M9 271 610 609 271 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=30430 $Y=15090 $D=1
M10 271 628 618 271 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.205e-14 PD=8.3e-07 PS=6.3e-07 $X=30770 $Y=15090 $D=1
M11 1258 609 271 271 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=8.3e-07 $X=30960 $Y=15090 $D=1
M12 271 339 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=31020 $Y=43090 $D=1
M13 643 628 1258 271 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.0125e-14 AS=3.85e-14 PD=8.7e-07 PS=8.3e-07 $X=31150 $Y=15090 $D=1
M14 271 339 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=31210 $Y=43090 $D=1
M15 1259 618 643 271 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.0125e-14 PD=4.6e-07 PS=8.7e-07 $X=31360 $Y=15160 $D=1
M16 271 339 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=31400 $Y=43090 $D=1
M17 271 624 1259 271 NMOS_VTL L=5e-08 W=9e-08 AD=3.58e-14 AS=1.26e-14 PD=1.12e-06 PS=4.6e-07 $X=31550 $Y=15160 $D=1
M18 271 339 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=31590 $Y=43090 $D=1
M19 624 643 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.58e-14 PD=1.11e-06 PS=1.12e-06 $X=31745 $Y=15090 $D=1
M20 271 643 624 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=31935 $Y=15090 $D=1
M21 271 273 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=31965 $Y=43090 $D=1
M22 271 273 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=32155 $Y=43090 $D=1
M23 271 23 628 271 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.69e-14 AS=3.36e-14 PD=1.14e-06 PS=7.4e-07 $X=32330 $Y=15090 $D=1
M24 271 273 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=32345 $Y=43090 $D=1
M25 1260 23 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.69e-14 PD=1.11e-06 PS=1.14e-06 $X=32535 $Y=15090 $D=1
M26 271 273 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=32535 $Y=43090 $D=1
M27 646 643 1260 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=32725 $Y=15090 $D=1
M28 271 288 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=32725 $Y=43090 $D=1
M29 1261 643 646 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=32915 $Y=15090 $D=1
M30 271 288 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=32915 $Y=43090 $D=1
M31 271 23 1261 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33105 $Y=15090 $D=1
M32 271 288 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33105 $Y=43090 $D=1
M33 1262 23 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33295 $Y=15090 $D=1
M34 271 288 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=33295 $Y=43090 $D=1
M35 646 643 1262 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33485 $Y=15090 $D=1
M36 1263 643 646 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33675 $Y=15090 $D=1
M37 271 23 1263 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.27e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33865 $Y=15090 $D=1
M38 38 646 271 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.27e-14 PD=6.7e-07 PS=1.11e-06 $X=34055 $Y=15090 $D=1
M39 271 646 38 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=34245 $Y=15090 $D=1
M40 38 646 271 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=34435 $Y=15090 $D=1
M41 271 646 38 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=34625 $Y=15090 $D=1
M42 38 646 271 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=34815 $Y=15090 $D=1
M43 271 646 38 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=35005 $Y=15090 $D=1
M44 38 646 271 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=35195 $Y=15090 $D=1
M45 271 646 38 271 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=35385 $Y=15090 $D=1
M46 271 693 695 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=42375 $Y=17890 $D=1
M47 695 693 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=42565 $Y=17890 $D=1
M48 271 693 695 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=42755 $Y=17890 $D=1
M49 695 693 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=42945 $Y=17890 $D=1
M50 196 704 695 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43135 $Y=17890 $D=1
M51 695 700 196 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43325 $Y=17890 $D=1
M52 196 700 695 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43515 $Y=17890 $D=1
M53 695 704 196 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43705 $Y=17890 $D=1
M54 196 704 695 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=43895 $Y=17890 $D=1
M55 695 700 196 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=44085 $Y=17890 $D=1
M56 196 700 695 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=44275 $Y=17890 $D=1
M57 695 704 196 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=44465 $Y=17890 $D=1
M58 394 421 719 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=45080 $Y=20095 $D=1
M59 719 450 394 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=45270 $Y=20095 $D=1
M60 723 426 719 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=45460 $Y=20095 $D=1
M61 719 706 723 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=45650 $Y=20095 $D=1
M62 723 721 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=46015 $Y=20095 $D=1
M63 271 458 723 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=46205 $Y=20095 $D=1
M64 726 727 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=46565 $Y=31890 $D=1
M65 271 727 726 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=46755 $Y=31890 $D=1
M66 1264 445 271 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=46945 $Y=31890 $D=1
M67 727 729 1264 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=47135 $Y=31890 $D=1
M68 726 729 393 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=47520 $Y=31890 $D=1
M69 393 729 726 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=47710 $Y=31890 $D=1
M70 726 445 393 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=47900 $Y=31890 $D=1
M71 393 445 726 271 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=48090 $Y=31890 $D=1
M72 502 504 506 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=3045 $Y=44490 $D=0
M73 23 506 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3235 $Y=44490 $D=0
M74 502 506 23 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3425 $Y=44490 $D=0
M75 23 506 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3615 $Y=44490 $D=0
M76 151 169 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=19980 $Y=33290 $D=0
M77 502 562 151 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=20170 $Y=33290 $D=0
M78 151 562 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=20360 $Y=33290 $D=0
M79 502 169 151 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=20550 $Y=33290 $D=0
M80 1245 271 609 502 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=30240 $Y=15995 $D=0
M81 502 610 1245 502 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=30430 $Y=15995 $D=0
M82 502 628 618 502 PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=3.3075e-14 PD=1.12e-06 PS=8.4e-07 $X=30770 $Y=15995 $D=0
M83 1246 609 502 502 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=30960 $Y=15890 $D=0
M84 630 339 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=31020 $Y=43680 $D=0
M85 643 618 1246 502 PMOS_VTL L=5e-08 W=4.2e-07 AD=4.245e-14 AS=5.88e-14 PD=1.16e-06 PS=1.12e-06 $X=31150 $Y=15890 $D=0
M86 502 339 630 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=31210 $Y=43680 $D=0
M87 1247 628 643 502 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=4.245e-14 PD=4.6e-07 PS=1.16e-06 $X=31360 $Y=16080 $D=0
M88 630 339 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=31400 $Y=43680 $D=0
M89 502 624 1247 502 PMOS_VTL L=5e-08 W=9e-08 AD=5.085e-14 AS=1.26e-14 PD=1.55e-06 PS=4.6e-07 $X=31550 $Y=16080 $D=0
M90 502 339 630 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=31590 $Y=43680 $D=0
M91 624 643 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=5.085e-14 PD=1.54e-06 PS=1.55e-06 $X=31745 $Y=15680 $D=0
M92 502 643 624 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=31935 $Y=15680 $D=0
M93 630 273 642 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=31965 $Y=43680 $D=0
M94 642 273 630 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=32155 $Y=43680 $D=0
M95 502 23 628 502 PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=5.04e-14 PD=1.57e-06 PS=9.5e-07 $X=32330 $Y=15790 $D=0
M96 630 273 642 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=32345 $Y=43680 $D=0
M97 646 23 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06 PS=1.57e-06 $X=32535 $Y=15680 $D=0
M98 642 273 630 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=32535 $Y=43680 $D=0
M99 502 643 646 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=32725 $Y=15680 $D=0
M100 271 288 642 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=32725 $Y=43680 $D=0
M101 646 643 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=32915 $Y=15680 $D=0
M102 642 288 271 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=32915 $Y=43680 $D=0
M103 502 23 646 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33105 $Y=15680 $D=0
M104 271 288 642 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33105 $Y=43680 $D=0
M105 646 23 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33295 $Y=15680 $D=0
M106 642 288 271 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=33295 $Y=43680 $D=0
M107 502 643 646 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33485 $Y=15680 $D=0
M108 646 643 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33675 $Y=15680 $D=0
M109 502 23 646 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33865 $Y=15680 $D=0
M110 38 646 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=34055 $Y=15680 $D=0
M111 502 646 38 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=34245 $Y=15680 $D=0
M112 38 646 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=34435 $Y=15680 $D=0
M113 502 646 38 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=34625 $Y=15680 $D=0
M114 38 646 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=34815 $Y=15680 $D=0
M115 502 646 38 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=35005 $Y=15680 $D=0
M116 38 646 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=35195 $Y=15680 $D=0
M117 502 646 38 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=35385 $Y=15680 $D=0
M118 196 693 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=42375 $Y=18480 $D=0
M119 502 693 196 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=42565 $Y=18480 $D=0
M120 196 693 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=42755 $Y=18480 $D=0
M121 502 693 196 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=42945 $Y=18480 $D=0
M122 1248 704 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43135 $Y=18480 $D=0
M123 196 700 1248 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43325 $Y=18480 $D=0
M124 1249 700 196 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43515 $Y=18480 $D=0
M125 502 704 1249 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43705 $Y=18480 $D=0
M126 1250 704 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=43895 $Y=18480 $D=0
M127 196 700 1250 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=44085 $Y=18480 $D=0
M128 1251 700 196 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=44275 $Y=18480 $D=0
M129 502 704 1251 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=44465 $Y=18480 $D=0
M130 1252 421 394 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=45080 $Y=19290 $D=0
M131 502 450 1252 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=45270 $Y=19290 $D=0
M132 1253 426 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=45460 $Y=19290 $D=0
M133 394 706 1253 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=1.9845e-13 AS=8.82e-14 PD=1.89e-06 PS=1.54e-06 $X=45650 $Y=19290 $D=0
M134 1254 721 394 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.9845e-13 PD=1.54e-06 PS=1.89e-06 $X=46015 $Y=19290 $D=0
M135 502 458 1254 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=46205 $Y=19290 $D=0
M136 393 727 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=46565 $Y=32480 $D=0
M137 502 727 393 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=46755 $Y=32480 $D=0
M138 727 445 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=46945 $Y=32480 $D=0
M139 502 729 727 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=47135 $Y=32480 $D=0
M140 393 729 728 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=47520 $Y=32480 $D=0
M141 1255 729 393 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=47710 $Y=32480 $D=0
M142 502 445 1255 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=47900 $Y=32480 $D=0
M143 728 445 502 502 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=48090 $Y=32480 $D=0
X10707 22 271 502 500 INV_X1 $T=1760 15000 0 180 $X=1265 $Y=13485
X10708 22 271 502 588 INV_X1 $T=2900 15000 1 0 $X=2785 $Y=13485
X10709 22 271 502 510 INV_X1 $T=5750 48600 0 0 $X=5635 $Y=48485
X10710 1154 271 502 43 INV_X1 $T=7840 51400 1 180 $X=7345 $Y=51285
X10711 958 271 502 528 INV_X1 $T=8220 26200 1 0 $X=8105 $Y=24685
X10712 765 271 502 512 INV_X1 $T=8790 23400 1 180 $X=8295 $Y=23285
X10713 966 271 502 50 INV_X1 $T=9170 54200 0 180 $X=8675 $Y=52685
X10714 959 271 502 774 INV_X1 $T=9740 31800 1 0 $X=9625 $Y=30285
X10715 772 271 502 84 INV_X1 $T=10310 29000 1 180 $X=9815 $Y=28885
X10716 529 271 502 516 INV_X1 $T=10500 17800 0 180 $X=10005 $Y=16285
X10717 967 271 502 525 INV_X1 $T=10120 43000 1 0 $X=10005 $Y=41485
X10718 524 271 502 970 INV_X1 $T=10880 48600 0 180 $X=10385 $Y=47085
X10719 63 271 502 57 INV_X1 $T=10690 48600 0 0 $X=10575 $Y=48485
X10720 526 271 502 67 INV_X1 $T=11260 20600 0 180 $X=10765 $Y=19085
X10721 981 271 502 40 INV_X1 $T=11070 43000 0 0 $X=10955 $Y=42885
X10722 513 271 502 82 INV_X1 $T=11830 40200 0 0 $X=11715 $Y=40085
X10723 779 271 502 534 INV_X1 $T=12400 9400 1 0 $X=12285 $Y=7885
X10724 1104 271 502 533 INV_X1 $T=12590 40200 1 0 $X=12475 $Y=38685
X10725 72 271 502 76 INV_X1 $T=12780 20600 0 0 $X=12665 $Y=20485
X10726 70 271 502 58 INV_X1 $T=13350 48600 1 180 $X=12855 $Y=48485
X10727 976 271 502 86 INV_X1 $T=14110 43000 0 180 $X=13615 $Y=41485
X10728 803 271 502 787 INV_X1 $T=14490 37400 0 180 $X=13995 $Y=35885
X10729 1106 271 502 105 INV_X1 $T=14870 15000 1 0 $X=14755 $Y=13485
X10730 85 271 502 108 INV_X1 $T=15250 45800 1 0 $X=15135 $Y=44285
X10731 982 271 502 80 INV_X1 $T=15630 54200 0 180 $X=15135 $Y=52685
X10732 795 271 502 650 INV_X1 $T=15440 26200 0 0 $X=15325 $Y=26085
X10733 86 271 502 134 INV_X1 $T=16010 51400 1 0 $X=15895 $Y=49885
X10734 117 271 502 121 INV_X1 $T=17150 26200 0 180 $X=16655 $Y=24685
X10735 783 271 502 986 INV_X1 $T=16770 37400 0 0 $X=16655 $Y=37285
X10736 109 271 502 560 INV_X1 $T=17150 20600 0 0 $X=17035 $Y=20485
X10737 553 271 502 987 INV_X1 $T=17340 31800 1 0 $X=17225 $Y=30285
X10738 802 271 502 145 INV_X1 $T=17530 31800 0 0 $X=17415 $Y=31685
X10739 801 271 502 125 INV_X1 $T=18100 29000 0 180 $X=17605 $Y=27485
X10740 693 271 502 91 INV_X1 $T=18100 40200 0 180 $X=17605 $Y=38685
X10741 191 271 502 137 INV_X1 $T=18290 12200 1 0 $X=18175 $Y=10685
X10742 151 271 502 130 INV_X1 $T=18670 34600 1 0 $X=18555 $Y=33085
X10743 793 271 502 989 INV_X1 $T=18670 45800 1 0 $X=18555 $Y=44285
X10744 561 271 502 812 INV_X1 $T=19430 17800 1 0 $X=19315 $Y=16285
X10745 564 271 502 141 INV_X1 $T=19810 43000 1 180 $X=19315 $Y=42885
X10746 185 271 502 99 INV_X1 $T=19620 9400 1 0 $X=19505 $Y=7885
X10747 991 271 502 163 INV_X1 $T=19810 51400 1 0 $X=19695 $Y=49885
X10748 157 271 502 123 INV_X1 $T=20000 6600 0 0 $X=19885 $Y=6485
X10749 166 271 502 198 INV_X1 $T=20000 9400 1 0 $X=19885 $Y=7885
X10750 225 271 502 187 INV_X1 $T=20000 26200 1 0 $X=19885 $Y=24685
X10751 816 271 502 992 INV_X1 $T=20570 37400 1 180 $X=20075 $Y=37285
X10752 778 271 502 144 INV_X1 $T=20190 43000 1 0 $X=20075 $Y=41485
X10753 201 271 502 60 INV_X1 $T=20380 6600 0 0 $X=20265 $Y=6485
X10754 119 271 502 566 INV_X1 $T=20760 29000 0 180 $X=20265 $Y=27485
X10755 1112 271 502 186 INV_X1 $T=20570 20600 0 0 $X=20455 $Y=20485
X10756 993 271 502 817 INV_X1 $T=20570 43000 1 0 $X=20455 $Y=41485
X10757 764 271 502 568 INV_X1 $T=20760 6600 0 0 $X=20645 $Y=6485
X10758 995 271 502 61 INV_X1 $T=21140 9400 1 0 $X=21025 $Y=7885
X10759 74 271 502 132 INV_X1 $T=21900 9400 0 180 $X=21405 $Y=7885
X10760 569 271 502 1179 INV_X1 $T=21520 17800 0 0 $X=21405 $Y=17685
X10761 188 271 502 149 INV_X1 $T=21900 34600 1 180 $X=21405 $Y=34485
X10762 116 271 502 178 INV_X1 $T=21520 51400 1 0 $X=21405 $Y=49885
X10763 98 271 502 1158 INV_X1 $T=22090 48600 1 0 $X=21975 $Y=47085
X10764 196 271 502 156 INV_X1 $T=22660 40200 1 180 $X=22165 $Y=40085
X10765 108 271 502 823 INV_X1 $T=22280 45800 0 0 $X=22165 $Y=45685
X10766 154 271 502 182 INV_X1 $T=23040 31800 0 180 $X=22545 $Y=30285
X10767 215 271 502 177 INV_X1 $T=23420 31800 0 180 $X=22925 $Y=30285
X10768 288 271 502 798 INV_X1 $T=23230 43000 1 0 $X=23115 $Y=41485
X10769 273 271 502 575 INV_X1 $T=23800 40200 1 180 $X=23305 $Y=40085
X10770 141 271 502 228 INV_X1 $T=23420 48600 1 0 $X=23305 $Y=47085
X10771 144 271 502 226 INV_X1 $T=23420 48600 0 0 $X=23305 $Y=48485
X10772 285 271 502 1004 INV_X1 $T=24180 6600 0 180 $X=23685 $Y=5085
X10773 1005 271 502 90 INV_X1 $T=24370 45800 0 180 $X=23875 $Y=44285
X10774 205 271 502 1007 INV_X1 $T=25320 6600 1 0 $X=25205 $Y=5085
X10775 831 271 502 828 INV_X1 $T=26270 37400 1 180 $X=25775 $Y=37285
X10776 577 271 502 237 INV_X1 $T=26270 15000 0 0 $X=26155 $Y=14885
X10777 1011 271 502 219 INV_X1 $T=26840 31800 0 180 $X=26345 $Y=30285
X10778 179 271 502 593 INV_X1 $T=26650 17800 1 0 $X=26535 $Y=16285
X10779 589 271 502 1122 INV_X1 $T=26840 6600 1 0 $X=26725 $Y=5085
X10780 128 271 502 595 INV_X1 $T=26840 12200 0 0 $X=26725 $Y=12085
X10781 594 271 502 171 INV_X1 $T=27220 31800 0 180 $X=26725 $Y=30285
X10782 207 271 502 235 INV_X1 $T=27030 9400 0 0 $X=26915 $Y=9285
X10783 224 271 502 244 INV_X1 $T=27220 17800 0 0 $X=27105 $Y=17685
X10784 1010 271 502 1009 INV_X1 $T=27600 37400 0 180 $X=27105 $Y=35885
X10785 240 271 502 249 INV_X1 $T=27410 9400 0 0 $X=27295 $Y=9285
X10786 366 271 502 236 INV_X1 $T=27980 15000 0 180 $X=27485 $Y=13485
X10787 112 271 502 233 INV_X1 $T=27980 20600 1 180 $X=27485 $Y=20485
X10788 339 271 502 305 INV_X1 $T=27600 43000 0 0 $X=27485 $Y=42885
X10789 840 271 502 200 INV_X1 $T=28170 3800 1 180 $X=27675 $Y=3685
X10790 260 271 502 328 INV_X1 $T=27790 23400 1 0 $X=27675 $Y=21885
X10791 292 271 502 315 INV_X1 $T=27980 48600 1 0 $X=27865 $Y=47085
X10792 247 271 502 1125 INV_X1 $T=28550 20600 0 180 $X=28055 $Y=19085
X10793 243 271 502 270 INV_X1 $T=28550 9400 1 0 $X=28435 $Y=7885
X10794 250 271 502 599 INV_X1 $T=29120 43000 1 180 $X=28625 $Y=42885
X10795 265 271 502 254 INV_X1 $T=29310 29000 1 0 $X=29195 $Y=27485
X10796 423 271 502 298 INV_X1 $T=29500 6600 1 0 $X=29385 $Y=5085
X10797 242 271 502 836 INV_X1 $T=29500 9400 1 0 $X=29385 $Y=7885
X10798 252 271 502 234 INV_X1 $T=29880 26200 1 180 $X=29385 $Y=26085
X10799 335 271 502 602 INV_X1 $T=30070 12200 0 180 $X=29575 $Y=10685
X10800 371 271 502 385 INV_X1 $T=30070 12200 1 180 $X=29575 $Y=12085
X10801 344 271 502 852 INV_X1 $T=29880 17800 0 0 $X=29765 $Y=17685
X10802 832 271 502 387 INV_X1 $T=30450 6600 1 180 $X=29955 $Y=6485
X10803 598 271 502 638 INV_X1 $T=30070 12200 0 0 $X=29955 $Y=12085
X10804 308 271 502 267 INV_X1 $T=30450 20600 1 180 $X=29955 $Y=20485
X10805 204 271 502 606 INV_X1 $T=30260 15000 1 0 $X=30145 $Y=13485
X10806 274 271 502 277 INV_X1 $T=30830 12200 1 180 $X=30335 $Y=12085
X10807 278 271 502 319 INV_X1 $T=30640 15000 1 0 $X=30525 $Y=13485
X10808 377 271 502 1008 INV_X1 $T=30640 17800 1 0 $X=30525 $Y=16285
X10809 69 271 502 290 INV_X1 $T=31020 17800 1 0 $X=30905 $Y=16285
X10810 623 271 502 261 INV_X1 $T=31780 26200 0 180 $X=31285 $Y=24685
X10811 453 271 502 853 INV_X1 $T=31590 12200 1 0 $X=31475 $Y=10685
X10812 854 271 502 614 INV_X1 $T=31970 26200 1 180 $X=31475 $Y=26085
X10813 1126 271 502 851 INV_X1 $T=32540 34600 1 180 $X=32045 $Y=34485
X10814 603 271 502 855 INV_X1 $T=33110 37400 0 180 $X=32615 $Y=35885
X10815 300 271 502 325 INV_X1 $T=34250 17800 1 180 $X=33755 $Y=17685
X10816 604 271 502 357 INV_X1 $T=34630 20600 1 180 $X=34135 $Y=20485
X10817 203 271 502 309 INV_X1 $T=34820 26200 1 180 $X=34325 $Y=26085
X10818 654 271 502 316 INV_X1 $T=35200 26200 0 180 $X=34705 $Y=24685
X10819 1240 271 502 667 INV_X1 $T=35770 17800 1 0 $X=35655 $Y=16285
X10820 209 271 502 146 INV_X1 $T=35960 23400 1 0 $X=35845 $Y=21885
X10821 1220 271 502 349 INV_X1 $T=36340 23400 0 0 $X=36225 $Y=23285
X10822 867 271 502 1165 INV_X1 $T=37290 26200 1 180 $X=36795 $Y=26085
X10823 665 271 502 1027 INV_X1 $T=37480 37400 0 180 $X=36985 $Y=35885
X10824 346 271 502 867 INV_X1 $T=37670 26200 1 180 $X=37175 $Y=26085
X10825 671 271 502 669 INV_X1 $T=38050 23400 1 180 $X=37555 $Y=23285
X10826 1035 271 502 880 INV_X1 $T=38240 23400 1 0 $X=38125 $Y=21885
X10827 375 271 502 1034 INV_X1 $T=38620 51400 0 180 $X=38125 $Y=49885
X10828 670 271 502 367 INV_X1 $T=38430 37400 1 0 $X=38315 $Y=35885
X10829 1037 271 502 879 INV_X1 $T=39570 34600 0 180 $X=39075 $Y=33085
X10830 396 271 502 386 INV_X1 $T=39380 20600 1 0 $X=39265 $Y=19085
X10831 679 271 502 837 INV_X1 $T=39570 12200 1 0 $X=39455 $Y=10685
X10832 682 271 502 692 INV_X1 $T=40330 20600 1 0 $X=40215 $Y=19085
X10833 684 271 502 1043 INV_X1 $T=40520 15000 1 0 $X=40405 $Y=13485
X10834 857 271 502 687 INV_X1 $T=40900 9400 1 0 $X=40785 $Y=7885
X10835 269 271 502 221 INV_X1 $T=42610 17800 0 180 $X=42115 $Y=16285
X10836 404 271 502 903 INV_X1 $T=42230 20600 1 0 $X=42115 $Y=19085
X10837 317 271 502 895 INV_X1 $T=42610 34600 1 180 $X=42115 $Y=34485
X10838 1048 271 502 401 INV_X1 $T=42990 20600 0 180 $X=42495 $Y=19085
X10839 680 271 502 412 INV_X1 $T=43370 34600 0 0 $X=43255 $Y=34485
X10840 418 271 502 410 INV_X1 $T=43940 15000 1 0 $X=43825 $Y=13485
X10841 903 271 502 703 INV_X1 $T=43940 20600 0 0 $X=43825 $Y=20485
X10842 378 271 502 419 INV_X1 $T=44700 37400 1 0 $X=44585 $Y=35885
X10843 407 271 502 432 INV_X1 $T=45650 26200 0 180 $X=45155 $Y=24685
X10844 706 271 502 403 INV_X1 $T=45650 20600 0 0 $X=45535 $Y=20485
X10845 389 271 502 427 INV_X1 $T=46220 37400 0 180 $X=45725 $Y=35885
X10846 477 271 502 462 INV_X1 $T=46030 15000 0 0 $X=45915 $Y=14885
X10847 721 271 502 416 INV_X1 $T=46030 20600 0 0 $X=45915 $Y=20485
X10848 910 271 502 911 INV_X1 $T=46030 31800 0 0 $X=45915 $Y=31685
X10849 263 271 502 456 INV_X1 $T=46600 51400 0 180 $X=46105 $Y=49885
X10850 216 271 502 426 INV_X1 $T=46790 20600 1 180 $X=46295 $Y=20485
X10851 718 271 502 291 INV_X1 $T=46790 48600 1 180 $X=46295 $Y=48485
X10852 442 271 502 461 INV_X1 $T=47550 15000 1 0 $X=47435 $Y=13485
X10853 1146 271 502 915 INV_X1 $T=48310 17800 1 180 $X=47815 $Y=17685
X10854 450 271 502 452 INV_X1 $T=47930 23400 1 0 $X=47815 $Y=21885
X10855 365 271 502 455 INV_X1 $T=47930 34600 1 0 $X=47815 $Y=33085
X10856 314 271 502 913 INV_X1 $T=49260 34600 1 180 $X=48765 $Y=34485
X10857 320 271 502 1073 INV_X1 $T=49830 20600 0 0 $X=49715 $Y=20485
X10858 583 271 502 927 INV_X1 $T=50400 20600 1 0 $X=50285 $Y=19085
X10859 746 271 502 1067 INV_X1 $T=51540 29000 1 180 $X=51045 $Y=28885
X10860 1071 271 502 931 INV_X1 $T=51540 31800 1 0 $X=51425 $Y=30285
X10861 482 271 502 929 INV_X1 $T=51920 12200 0 0 $X=51805 $Y=12085
X10862 493 271 502 494 INV_X1 $T=53630 20600 1 0 $X=53515 $Y=19085
X10863 496 271 502 451 INV_X1 $T=53820 17800 1 0 $X=53705 $Y=16285
X10864 271 502 962 29 ICV_5 $T=7080 48600 1 0 $X=6965 $Y=47085
X10865 271 502 770 771 ICV_5 $T=9740 23400 0 0 $X=9625 $Y=23285
X10866 271 502 768 775 ICV_5 $T=9740 40200 1 0 $X=9625 $Y=38685
X10867 271 502 975 790 ICV_5 $T=12970 34600 1 0 $X=12855 $Y=33085
X10868 271 502 780 107 ICV_5 $T=13730 9400 1 0 $X=13615 $Y=7885
X10869 271 502 794 111 ICV_5 $T=15060 34600 0 0 $X=14945 $Y=34485
X10870 271 502 71 116 ICV_5 $T=16960 40200 0 0 $X=16845 $Y=40085
X10871 271 502 202 143 ICV_5 $T=22660 17800 1 0 $X=22545 $Y=16285
X10872 271 502 124 208 ICV_5 $T=24180 26200 0 0 $X=24065 $Y=26085
X10873 271 502 465 458 ICV_5 $T=47170 20600 0 0 $X=47055 $Y=20485
X10874 271 502 1060 918 ICV_5 $T=47550 51400 1 0 $X=47435 $Y=49885
X10875 271 502 924 483 ICV_5 $T=50020 12200 1 0 $X=49905 $Y=10685
X10876 271 502 454 1153 ICV_5 $T=51920 20600 0 0 $X=51805 $Y=20485
X10877 271 502 947 1077 ICV_5 $T=55910 29000 0 0 $X=55795 $Y=28885
X10878 507 502 501 759 271 NOR2_X1 $T=2330 48600 1 0 $X=2215 $Y=47085
X10879 507 502 760 961 271 NOR2_X1 $T=4800 45800 1 180 $X=4115 $Y=45685
X10880 768 502 960 967 271 NOR2_X1 $T=8410 40200 0 0 $X=8295 $Y=40085
X10881 973 502 517 524 271 NOR2_X1 $T=9550 45800 0 0 $X=9435 $Y=45685
X10882 773 502 527 969 271 NOR2_X1 $T=10310 26200 0 0 $X=10195 $Y=26085
X10883 774 502 62 527 271 NOR2_X1 $T=10310 29000 0 0 $X=10195 $Y=28885
X10884 55 502 67 511 271 NOR2_X1 $T=10500 17800 1 0 $X=10385 $Y=16285
X10885 775 502 960 550 271 NOR2_X1 $T=10500 37400 0 0 $X=10385 $Y=37285
X10886 529 502 76 118 271 NOR2_X1 $T=12210 20600 1 0 $X=12095 $Y=19085
X10887 533 502 87 783 271 NOR2_X1 $T=12590 37400 1 0 $X=12475 $Y=35885
X10888 79 502 84 64 271 NOR2_X1 $T=12970 26200 0 0 $X=12855 $Y=26085
X10889 113 502 72 75 271 NOR2_X1 $T=13160 20600 0 0 $X=13045 $Y=20485
X10890 529 502 72 142 271 NOR2_X1 $T=13730 17800 1 0 $X=13615 $Y=16285
X10891 544 502 529 978 271 NOR2_X1 $T=14680 20600 0 180 $X=13995 $Y=19085
X10892 76 502 106 115 271 NOR2_X1 $T=15250 23400 0 0 $X=15135 $Y=23285
X10893 120 502 693 981 271 NOR2_X1 $T=15820 40200 1 180 $X=15135 $Y=40085
X10894 790 502 101 984 271 NOR2_X1 $T=16010 31800 1 180 $X=15325 $Y=31685
X10895 550 502 980 139 271 NOR2_X1 $T=16580 37400 1 0 $X=16465 $Y=35885
X10896 1158 502 546 83 271 NOR2_X1 $T=18100 48600 0 180 $X=17415 $Y=47085
X10897 139 502 554 562 271 NOR2_X1 $T=18670 34600 0 180 $X=17985 $Y=33085
X10898 812 502 121 994 271 NOR2_X1 $T=20570 17800 1 0 $X=20455 $Y=16285
X10899 196 502 174 1000 271 NOR2_X1 $T=22850 34600 1 180 $X=22165 $Y=34485
X10900 196 502 578 1185 271 NOR2_X1 $T=23610 34600 0 0 $X=23495 $Y=34485
X10901 196 502 1218 1233 271 NOR2_X1 $T=27030 31800 1 180 $X=26345 $Y=31685
X10902 1015 502 1014 194 271 NOR2_X1 $T=28360 40200 0 180 $X=27675 $Y=38685
X10903 196 502 1161 1191 271 NOR2_X1 $T=28360 31800 0 0 $X=28245 $Y=31685
X10904 273 502 798 323 271 NOR2_X1 $T=28360 43000 1 0 $X=28245 $Y=41485
X10905 598 502 607 278 271 NOR2_X1 $T=29690 15000 1 0 $X=29575 $Y=13485
X10906 638 502 607 293 271 NOR2_X1 $T=30070 12200 1 0 $X=29955 $Y=10685
X10907 273 502 288 318 271 NOR2_X1 $T=30260 43000 1 0 $X=30145 $Y=41485
X10908 196 502 1162 621 271 NOR2_X1 $T=31970 31800 1 180 $X=31285 $Y=31685
X10909 575 502 288 370 271 NOR2_X1 $T=32160 43000 0 180 $X=31475 $Y=41485
X10910 196 502 613 856 271 NOR2_X1 $T=32540 31800 0 180 $X=31855 $Y=30285
X10911 196 502 651 652 271 NOR2_X1 $T=34440 31800 1 0 $X=34325 $Y=30285
X10912 662 502 69 330 271 NOR2_X1 $T=34820 12200 1 0 $X=34705 $Y=10685
X10913 662 502 290 355 271 NOR2_X1 $T=36910 9400 0 0 $X=36795 $Y=9285
X10914 196 502 668 1032 271 NOR2_X1 $T=37100 29000 0 0 $X=36985 $Y=28885
X10915 196 502 675 878 271 NOR2_X1 $T=37860 20600 0 0 $X=37745 $Y=20485
X10916 196 502 1167 883 271 NOR2_X1 $T=39190 29000 0 0 $X=39075 $Y=28885
X10917 386 502 681 886 271 NOR2_X1 $T=40710 23400 1 180 $X=40025 $Y=23285
X10918 680 502 697 373 271 NOR2_X1 $T=40900 40200 0 180 $X=40215 $Y=38685
X10919 196 502 392 1200 271 NOR2_X1 $T=40520 26200 0 0 $X=40405 $Y=26085
X10920 391 502 378 884 271 NOR2_X1 $T=42040 37400 1 0 $X=41925 $Y=35885
X10921 196 502 696 1235 271 NOR2_X1 $T=42990 26200 1 0 $X=42875 $Y=24685
X10922 365 502 326 1049 271 NOR2_X1 $T=42990 37400 0 0 $X=42875 $Y=37285
X10923 1051 502 702 424 271 NOR2_X1 $T=44510 29000 1 0 $X=44395 $Y=27485
X10924 196 502 905 1206 271 NOR2_X1 $T=45460 26200 1 180 $X=44775 $Y=26085
X10925 493 502 720 440 271 NOR2_X1 $T=46790 17800 1 180 $X=46105 $Y=17685
X10926 196 502 1143 1222 271 NOR2_X1 $T=46790 26200 1 180 $X=46105 $Y=26085
X10927 724 502 421 917 271 NOR2_X1 $T=47740 29000 0 0 $X=47625 $Y=28885
X10928 196 502 919 731 271 NOR2_X1 $T=49070 26200 1 180 $X=48385 $Y=26085
X10929 196 502 1068 734 271 NOR2_X1 $T=50780 23400 0 180 $X=50095 $Y=21885
X10930 196 502 1065 930 271 NOR2_X1 $T=51350 15000 0 180 $X=50665 $Y=13485
X10931 196 502 934 1145 271 NOR2_X1 $T=50970 20600 0 0 $X=50855 $Y=20485
X10932 196 502 932 1210 271 NOR2_X1 $T=51540 17800 1 0 $X=51425 $Y=16285
X10933 927 502 943 710 271 NOR2_X1 $T=51920 20600 1 0 $X=51805 $Y=19085
X10934 196 502 937 1078 271 NOR2_X1 $T=54580 15000 0 180 $X=53895 $Y=13485
X10935 196 502 752 942 271 NOR2_X1 $T=55720 15000 1 180 $X=55035 $Y=14885
X10936 196 502 1080 946 271 NOR2_X1 $T=56480 20600 0 180 $X=55795 $Y=19085
X11324 511 119 502 577 777 516 271 AOI22_X1 $T=8980 15000 0 0 $X=8865 $Y=14885
X11325 84 79 502 62 773 774 271 AOI22_X1 $T=9550 29000 1 0 $X=9435 $Y=27485
X11326 520 525 502 767 42 59 271 AOI22_X1 $T=9930 51400 1 0 $X=9815 $Y=49885
X11327 516 106 502 92 78 522 271 AOI22_X1 $T=10310 15000 1 0 $X=10195 $Y=13485
X11328 151 958 502 765 778 130 271 AOI22_X1 $T=10880 29000 0 0 $X=10765 $Y=28885
X11329 511 762 502 202 65 516 271 AOI22_X1 $T=11070 17800 1 0 $X=10955 $Y=16285
X11330 151 87 502 1104 49 130 271 AOI22_X1 $T=12020 40200 0 180 $X=10955 $Y=38685
X11331 109 764 502 76 779 531 271 AOI22_X1 $T=11260 9400 0 0 $X=11145 $Y=9285
X11332 118 81 502 76 780 515 271 AOI22_X1 $T=12400 9400 0 180 $X=11335 $Y=7885
X11333 151 772 502 79 85 130 271 AOI22_X1 $T=11640 31800 1 0 $X=11525 $Y=30285
X11334 1102 83 502 781 782 91 271 AOI22_X1 $T=12780 48600 0 180 $X=11715 $Y=47085
X11335 522 198 502 67 73 68 271 AOI22_X1 $T=12210 15000 0 0 $X=12095 $Y=14885
X11336 532 96 502 89 1110 789 271 AOI22_X1 $T=12400 29000 1 0 $X=12285 $Y=27485
X11337 1217 1103 502 798 972 86 271 AOI22_X1 $T=12590 43000 0 0 $X=12475 $Y=42885
X11338 535 76 502 72 977 78 271 AOI22_X1 $T=12780 17800 1 0 $X=12665 $Y=16285
X11339 151 101 502 975 976 130 271 AOI22_X1 $T=12780 37400 0 0 $X=12665 $Y=37285
X11340 783 787 502 87 1157 533 271 AOI22_X1 $T=13160 37400 1 0 $X=13045 $Y=35885
X11341 118 92 502 76 1106 73 271 AOI22_X1 $T=14870 15000 0 180 $X=13805 $Y=13485
X11342 75 577 502 112 1109 118 271 AOI22_X1 $T=16580 17800 1 180 $X=15515 $Y=17685
X11343 976 288 502 798 1103 86 271 AOI22_X1 $T=15630 43000 1 0 $X=15515 $Y=41485
X11344 75 224 502 762 1113 118 271 AOI22_X1 $T=16580 17800 0 0 $X=16465 $Y=17685
X11345 131 1115 502 273 1217 71 271 AOI22_X1 $T=18290 43000 0 180 $X=17225 $Y=41485
X11346 116 575 502 273 1115 71 271 AOI22_X1 $T=18480 40200 1 180 $X=17415 $Y=40085
X11347 75 225 502 204 1118 109 271 AOI22_X1 $T=18100 20600 0 0 $X=17985 $Y=20485
X11348 75 119 502 112 811 109 271 AOI22_X1 $T=18290 23400 1 0 $X=18175 $Y=21885
X11349 91 130 502 992 821 156 271 AOI22_X1 $T=18480 37400 0 0 $X=18365 $Y=37285
X11350 545 121 502 117 206 809 271 AOI22_X1 $T=19810 15000 1 180 $X=18745 $Y=14885
X11351 557 117 502 121 569 974 271 AOI22_X1 $T=19810 20600 0 180 $X=18745 $Y=19085
X11352 561 121 502 117 1159 158 271 AOI22_X1 $T=19430 15000 1 0 $X=19315 $Y=13485
X11353 1178 805 502 225 154 151 271 AOI22_X1 $T=19430 29000 0 0 $X=19315 $Y=28885
X11354 805 117 502 119 188 151 271 AOI22_X1 $T=21330 29000 1 180 $X=20265 $Y=28885
X11355 571 121 502 117 582 140 271 AOI22_X1 $T=21900 9400 1 180 $X=20835 $Y=9285
X11356 152 117 502 121 271 1118 271 AOI22_X1 $T=20950 20600 0 0 $X=20835 $Y=20485
X11357 1118 117 502 121 573 811 271 AOI22_X1 $T=21900 23400 0 180 $X=20835 $Y=21885
X11358 567 989 502 292 818 564 271 AOI22_X1 $T=20950 45800 1 0 $X=20835 $Y=44285
X11359 152 121 502 117 1182 572 271 AOI22_X1 $T=21330 20600 1 0 $X=21215 $Y=19085
X11360 1184 805 502 762 215 151 271 AOI22_X1 $T=22280 29000 1 180 $X=21215 $Y=28885
X11361 144 305 502 339 993 778 271 AOI22_X1 $T=22280 43000 1 0 $X=22165 $Y=41485
X11362 220 828 502 580 183 824 271 AOI22_X1 $T=24750 37400 1 180 $X=23685 $Y=37285
X11363 74 270 502 576 239 585 271 AOI22_X1 $T=24560 9400 1 0 $X=24445 $Y=7885
X11364 230 1009 502 219 831 830 271 AOI22_X1 $T=26460 37400 0 180 $X=25395 $Y=35885
X11365 478 825 502 283 590 479 271 AOI22_X1 $T=25510 43000 1 0 $X=25395 $Y=41485
X11366 1188 253 502 368 594 146 271 AOI22_X1 $T=27030 26200 0 180 $X=25965 $Y=24685
X11367 1121 253 502 303 1011 146 271 AOI22_X1 $T=27030 29000 0 180 $X=25965 $Y=27485
X11368 595 371 502 1124 1123 597 271 AOI22_X1 $T=27220 12200 0 0 $X=27105 $Y=12085
X11369 1013 839 502 171 1010 838 271 AOI22_X1 $T=28170 34600 1 180 $X=27105 $Y=34485
X11370 92 277 502 385 597 128 271 AOI22_X1 $T=29120 12200 1 180 $X=28055 $Y=12085
X11371 221 368 502 252 600 269 271 AOI22_X1 $T=28170 23400 1 0 $X=28055 $Y=21885
X11372 204 852 502 1219 1016 266 271 AOI22_X1 $T=28360 17800 0 0 $X=28245 $Y=17685
X11373 718 847 502 283 1017 478 271 AOI22_X1 $T=29310 48600 0 180 $X=28245 $Y=47085
X11374 593 356 502 344 266 606 271 AOI22_X1 $T=29120 15000 0 0 $X=29005 $Y=14885
X11375 294 851 502 614 262 848 271 AOI22_X1 $T=30830 34600 1 180 $X=29765 $Y=34485
X11376 258 854 502 614 1020 282 271 AOI22_X1 $T=30640 26200 0 0 $X=30525 $Y=26085
X11377 362 308 502 335 634 278 271 AOI22_X1 $T=30830 12200 0 0 $X=30715 $Y=12085
X11378 362 366 502 303 850 293 271 AOI22_X1 $T=31970 6600 0 180 $X=30905 $Y=5085
X11379 362 252 502 620 331 278 271 AOI22_X1 $T=31020 15000 1 0 $X=30905 $Y=13485
X11380 479 295 502 603 284 478 271 AOI22_X1 $T=32540 48600 1 180 $X=31475 $Y=48485
X11381 293 368 502 371 633 362 271 AOI22_X1 $T=31970 6600 1 0 $X=31855 $Y=5085
X11382 278 853 502 607 334 1022 271 AOI22_X1 $T=31970 12200 1 0 $X=31855 $Y=10685
X11383 1128 1127 502 644 1126 625 271 AOI22_X1 $T=33490 34600 0 180 $X=32425 $Y=33085
X11384 629 389 502 250 302 271 271 AOI22_X1 $T=32540 40200 1 0 $X=32425 $Y=38685
X11385 479 639 502 295 324 478 271 AOI22_X1 $T=33490 48600 1 180 $X=32425 $Y=48485
X11386 660 292 502 315 636 635 271 AOI22_X1 $T=33680 48600 0 180 $X=32615 $Y=47085
X11387 634 290 502 69 684 331 271 AOI22_X1 $T=33680 15000 1 0 $X=33565 $Y=13485
X11388 69 303 502 247 1240 290 271 AOI22_X1 $T=33680 17800 1 0 $X=33565 $Y=16285
X11389 478 639 502 653 862 479 271 AOI22_X1 $T=34250 51400 1 0 $X=34135 $Y=49885
X11390 1132 339 502 305 329 647 271 AOI22_X1 $T=35390 45800 1 180 $X=34325 $Y=45685
X11391 329 315 502 292 327 1024 271 AOI22_X1 $T=34630 48600 1 0 $X=34515 $Y=47085
X11392 330 679 502 69 1164 661 271 AOI22_X1 $T=34820 6600 1 0 $X=34705 $Y=5085
X11393 629 430 502 888 641 322 271 AOI22_X1 $T=36150 40200 1 180 $X=35085 $Y=40085
X11394 370 430 502 888 657 318 271 AOI22_X1 $T=35200 43000 0 0 $X=35085 $Y=42885
X11395 863 1221 502 316 645 864 271 AOI22_X1 $T=36530 31800 1 180 $X=35465 $Y=31685
X11396 1040 292 502 315 342 660 271 AOI22_X1 $T=35580 48600 1 0 $X=35465 $Y=47085
X11397 370 389 502 670 1132 318 271 AOI22_X1 $T=36720 43000 0 180 $X=35655 $Y=41485
X11398 372 669 502 349 1029 346 271 AOI22_X1 $T=37290 26200 0 180 $X=36225 $Y=24685
X11399 676 671 502 1220 873 867 271 AOI22_X1 $T=37670 23400 1 180 $X=36605 $Y=23285
X11400 663 326 502 697 865 364 271 AOI22_X1 $T=37290 45800 1 0 $X=37175 $Y=44285
X11401 881 879 502 669 358 876 271 AOI22_X1 $T=38620 31800 1 180 $X=37555 $Y=31685
X11402 318 317 502 314 871 370 271 AOI22_X1 $T=37860 43000 0 0 $X=37745 $Y=42885
X11403 685 292 502 315 375 1024 271 AOI22_X1 $T=38050 48600 1 0 $X=37935 $Y=47085
X11404 479 347 502 665 374 478 271 AOI22_X1 $T=38050 48600 0 0 $X=37935 $Y=48485
X11405 352 269 502 221 1039 686 271 AOI22_X1 $T=38810 17800 1 0 $X=38695 $Y=16285
X11406 370 391 502 347 869 318 271 AOI22_X1 $T=39760 43000 1 180 $X=38695 $Y=42885
X11407 890 292 502 315 1041 1040 271 AOI22_X1 $T=39000 48600 1 0 $X=38885 $Y=47085
X11408 882 655 502 221 382 379 271 AOI22_X1 $T=40520 15000 0 180 $X=39455 $Y=13485
X11409 382 357 502 304 885 1039 271 AOI22_X1 $T=40710 17800 0 180 $X=39645 $Y=16285
X11410 395 1134 502 692 1037 673 271 AOI22_X1 $T=39760 31800 1 0 $X=39645 $Y=30285
X11411 364 378 502 380 678 663 271 AOI22_X1 $T=39760 43000 0 0 $X=39645 $Y=42885
X11412 656 221 502 269 388 891 271 AOI22_X1 $T=39950 9400 1 0 $X=39835 $Y=7885
X11413 1050 269 502 221 690 332 271 AOI22_X1 $T=40900 9400 1 180 $X=39835 $Y=9285
X11414 1047 456 502 347 1136 478 271 AOI22_X1 $T=41660 48600 1 180 $X=40595 $Y=48485
X11415 896 269 502 221 411 891 271 AOI22_X1 $T=41850 6600 1 180 $X=40785 $Y=6485
X11416 690 304 502 357 1042 388 271 AOI22_X1 $T=41850 9400 1 180 $X=40785 $Y=9285
X11417 686 269 502 221 409 691 271 AOI22_X1 $T=40900 15000 1 0 $X=40785 $Y=13485
X11418 889 1138 502 1135 1045 892 271 AOI22_X1 $T=41850 29000 1 180 $X=40785 $Y=28885
X11419 663 393 502 359 1038 364 271 AOI22_X1 $T=40900 45800 1 0 $X=40785 $Y=44285
X11420 1043 221 502 269 701 379 271 AOI22_X1 $T=42230 15000 1 0 $X=42115 $Y=13485
X11421 404 401 502 1048 406 903 271 AOI22_X1 $T=42230 20600 0 0 $X=42115 $Y=20485
X11422 691 269 502 221 438 898 271 AOI22_X1 $T=42420 12200 0 0 $X=42305 $Y=12085
X11423 1139 456 502 670 1052 479 271 AOI22_X1 $T=42800 51400 1 0 $X=42685 $Y=49885
X11424 1139 718 502 317 1055 479 271 AOI22_X1 $T=43180 48600 1 0 $X=43065 $Y=47085
X11425 364 326 502 430 428 271 271 AOI22_X1 $T=43750 40200 1 0 $X=43635 $Y=38685
X11426 478 317 502 359 1057 479 271 AOI22_X1 $T=44700 45800 1 180 $X=43635 $Y=45685
X11427 714 718 502 456 420 901 271 AOI22_X1 $T=44130 48600 1 0 $X=44015 $Y=47085
X11428 364 393 502 391 422 271 271 AOI22_X1 $T=45270 43000 0 180 $X=44205 $Y=41485
X11429 364 380 502 314 1054 271 271 AOI22_X1 $T=45460 37400 1 180 $X=44395 $Y=37285
X11430 701 304 502 357 1141 438 271 AOI22_X1 $T=44700 12200 0 0 $X=44585 $Y=12085
X11431 478 359 502 718 1058 901 271 AOI22_X1 $T=44700 45800 0 0 $X=44585 $Y=45685
X11432 364 365 502 389 722 271 271 AOI22_X1 $T=45460 40200 0 0 $X=45345 $Y=40085
X11433 479 391 502 456 1063 716 271 AOI22_X1 $T=46410 37400 0 0 $X=46295 $Y=37285
X11434 725 326 502 380 468 732 271 AOI22_X1 $T=47930 48600 0 180 $X=46865 $Y=47085
X11435 716 718 502 430 1225 479 271 AOI22_X1 $T=48500 37400 0 180 $X=47435 $Y=35885
X11436 909 456 502 718 933 713 271 AOI22_X1 $T=47740 43000 1 0 $X=47625 $Y=41485
X11437 909 718 502 378 737 478 271 AOI22_X1 $T=48120 40200 1 0 $X=48005 $Y=38685
X11438 478 697 502 456 738 713 271 AOI22_X1 $T=49070 43000 1 180 $X=48005 $Y=42885
X11439 478 314 502 393 470 479 271 AOI22_X1 $T=50020 43000 0 0 $X=49905 $Y=42885
X11440 927 1146 502 1073 1147 477 271 AOI22_X1 $T=50210 17800 0 0 $X=50095 $Y=17685
X11441 741 926 502 416 1071 735 271 AOI22_X1 $T=50210 31800 1 0 $X=50095 $Y=30285
X11442 479 389 502 456 1070 743 271 AOI22_X1 $T=51350 40200 0 180 $X=50285 $Y=38685
X11443 745 931 502 439 1148 928 271 AOI22_X1 $T=51540 26200 1 180 $X=50475 $Y=26085
X11444 479 378 502 680 744 478 271 AOI22_X1 $T=51540 43000 0 180 $X=50475 $Y=41485
X11445 750 935 502 1073 484 748 271 AOI22_X1 $T=52680 23400 1 180 $X=51615 $Y=23285
X11446 1150 1077 502 720 746 751 271 AOI22_X1 $T=53630 31800 1 0 $X=53515 $Y=30285
X11447 1081 940 502 1153 947 1083 271 AOI22_X1 $T=55530 26200 1 0 $X=55415 $Y=24685
X12224 500 1 271 502 948 271 AND2_X1 $T=1000 3800 0 0 $X=885 $Y=3685
X12225 500 2 271 502 949 271 AND2_X1 $T=1000 9400 1 0 $X=885 $Y=7885
X12226 500 3 271 502 1087 271 AND2_X1 $T=1000 12200 0 0 $X=885 $Y=12085
X12227 500 4 271 502 1088 271 AND2_X1 $T=1000 17800 0 0 $X=885 $Y=17685
X12228 500 9 271 502 48 271 AND2_X1 $T=1760 31800 1 180 $X=885 $Y=31685
X12229 500 10 271 502 1086 271 AND2_X1 $T=1760 37400 0 180 $X=885 $Y=35885
X12230 500 5 271 502 950 271 AND2_X1 $T=1190 9400 0 0 $X=1075 $Y=9285
X12231 500 11 271 502 1090 271 AND2_X1 $T=1760 23400 1 0 $X=1645 $Y=21885
X12232 588 12 271 502 952 271 AND2_X1 $T=1760 40200 0 0 $X=1645 $Y=40085
X12233 588 13 271 502 45 271 AND2_X1 $T=2710 26200 1 180 $X=1835 $Y=26085
X12234 500 14 271 502 758 271 AND2_X1 $T=2140 37400 1 0 $X=2025 $Y=35885
X12235 500 27 271 502 1226 271 AND2_X1 $T=3090 3800 0 180 $X=2215 $Y=2285
X12236 500 16 271 502 953 271 AND2_X1 $T=2330 6600 0 0 $X=2215 $Y=6485
X12237 500 17 271 502 1091 271 AND2_X1 $T=2330 15000 0 0 $X=2215 $Y=14885
X12238 588 18 271 502 954 271 AND2_X1 $T=2330 23400 0 0 $X=2215 $Y=23285
X12239 500 19 271 502 1228 271 AND2_X1 $T=2330 29000 1 0 $X=2215 $Y=27485
X12240 500 25 271 502 955 271 AND2_X1 $T=2330 34600 1 0 $X=2215 $Y=33085
X12241 500 26 271 502 505 271 AND2_X1 $T=2330 34600 0 0 $X=2215 $Y=34485
X12242 588 20 271 502 1092 271 AND2_X1 $T=2330 37400 0 0 $X=2215 $Y=37285
X12243 588 21 271 502 956 271 AND2_X1 $T=2330 43000 1 0 $X=2215 $Y=41485
X12244 588 28 271 502 1093 271 AND2_X1 $T=2520 40200 0 0 $X=2405 $Y=40085
X12245 500 31 271 502 1094 271 AND2_X1 $T=3090 15000 0 0 $X=2975 $Y=14885
X12246 588 32 271 502 1229 271 AND2_X1 $T=3090 34600 1 0 $X=2975 $Y=33085
X12247 500 33 271 502 1096 271 AND2_X1 $T=3470 20600 1 0 $X=3355 $Y=19085
X12248 500 34 271 502 957 271 AND2_X1 $T=3660 12200 0 0 $X=3545 $Y=12085
X12249 588 36 271 502 1095 271 AND2_X1 $T=4420 29000 1 180 $X=3545 $Y=28885
X12250 500 35 271 502 1097 271 AND2_X1 $T=3850 9400 0 0 $X=3735 $Y=9285
X12251 588 37 271 502 761 271 AND2_X1 $T=4230 20600 1 0 $X=4115 $Y=19085
X12252 500 39 271 502 1171 271 AND2_X1 $T=4420 29000 0 0 $X=4305 $Y=28885
X12253 588 41 271 502 509 271 AND2_X1 $T=5370 37400 0 0 $X=5255 $Y=37285
X12254 510 42 271 502 763 271 AND2_X1 $T=6320 54200 0 180 $X=5445 $Y=52685
X12255 510 43 271 502 1098 271 AND2_X1 $T=6320 54200 1 0 $X=6205 $Y=52685
X12256 500 44 271 502 1099 271 AND2_X1 $T=6510 3800 0 0 $X=6395 $Y=3685
X12257 500 1214 271 502 1100 1265 AND2_X1 $T=6890 1000 0 0 $X=6775 $Y=885
X12258 510 50 271 502 1101 271 AND2_X1 $T=8030 54200 1 0 $X=7915 $Y=52685
X12259 500 54 271 502 968 1265 AND2_X1 $T=9930 1000 0 0 $X=9815 $Y=885
X12260 529 68 271 502 535 271 AND2_X1 $T=12020 17800 0 0 $X=11905 $Y=17685
X12261 500 77 271 502 785 271 AND2_X1 $T=13920 3800 0 180 $X=13045 $Y=2285
X12262 500 88 271 502 1105 271 AND2_X1 $T=14680 3800 0 180 $X=13805 $Y=2285
X12263 500 102 271 502 792 1265 AND2_X1 $T=15630 1000 1 180 $X=14755 $Y=885
X12264 500 110 271 502 551 271 AND2_X1 $T=15820 3800 1 0 $X=15705 $Y=2285
X12265 500 122 271 502 1114 1265 AND2_X1 $T=16960 1000 0 0 $X=16845 $Y=885
X12266 109 125 271 502 805 271 AND2_X1 $T=17530 29000 0 0 $X=17415 $Y=28885
X12267 588 150 271 502 810 271 AND2_X1 $T=20000 3800 0 180 $X=19125 $Y=2285
X12268 813 156 271 502 1116 271 AND2_X1 $T=20190 37400 1 180 $X=19315 $Y=37285
X12269 813 162 271 502 816 271 AND2_X1 $T=20190 37400 1 0 $X=20075 $Y=35885
X12270 510 163 271 502 148 271 AND2_X1 $T=20380 54200 1 0 $X=20265 $Y=52685
X12271 588 167 271 502 997 1265 AND2_X1 $T=20950 1000 0 0 $X=20835 $Y=885
X12272 155 193 271 502 578 271 AND2_X1 $T=23040 34600 1 0 $X=22925 $Y=33085
X12273 588 1215 271 502 1187 1265 AND2_X1 $T=25890 1000 0 0 $X=25775 $Y=885
X12274 510 229 271 502 835 271 AND2_X1 $T=26080 54200 1 0 $X=25965 $Y=52685
X12275 510 251 271 502 272 271 AND2_X1 $T=28360 51400 0 0 $X=28245 $Y=51285
X12276 195 255 271 502 1161 271 AND2_X1 $T=28550 31800 1 0 $X=28435 $Y=30285
X12277 510 264 271 502 1192 271 AND2_X1 $T=29120 51400 0 0 $X=29005 $Y=51285
X12278 588 275 271 502 1193 1265 AND2_X1 $T=30450 1000 0 0 $X=30335 $Y=885
X12279 510 299 271 502 1195 271 AND2_X1 $T=32350 51400 0 0 $X=32235 $Y=51285
X12280 510 306 271 502 1130 271 AND2_X1 $T=33110 51400 0 0 $X=32995 $Y=51285
X12281 588 311 271 502 1129 1265 AND2_X1 $T=34250 1000 1 180 $X=33375 $Y=885
X12282 510 343 271 502 1131 271 AND2_X1 $T=36530 54200 0 180 $X=35655 $Y=52685
X12283 588 348 271 502 872 1265 AND2_X1 $T=36530 1000 0 0 $X=36415 $Y=885
X12284 510 360 271 502 1198 271 AND2_X1 $T=37100 51400 0 0 $X=36985 $Y=51285
X12285 510 381 271 502 1133 271 AND2_X1 $T=40140 51400 1 180 $X=39265 $Y=51285
X12286 588 390 271 502 376 1265 AND2_X1 $T=40520 1000 0 0 $X=40405 $Y=885
X12287 510 399 271 502 1201 271 AND2_X1 $T=41090 51400 0 0 $X=40975 $Y=51285
X12288 588 402 271 502 1234 271 AND2_X1 $T=42990 3800 0 180 $X=42115 $Y=2285
X12289 588 408 271 502 1204 271 AND2_X1 $T=42990 3800 0 0 $X=42875 $Y=3685
X12290 510 431 271 502 1223 271 AND2_X1 $T=45460 51400 1 0 $X=45345 $Y=49885
X12291 1061 1207 271 502 1143 271 AND2_X1 $T=46410 26200 0 180 $X=45535 $Y=24685
X12292 315 271 271 502 725 271 AND2_X1 $T=45650 45800 0 0 $X=45535 $Y=45685
X12293 510 437 271 502 417 271 AND2_X1 $T=46030 51400 0 0 $X=45915 $Y=51285
X12294 588 441 271 502 709 1265 AND2_X1 $T=46980 1000 1 180 $X=46105 $Y=885
X12295 588 444 271 502 1208 1265 AND2_X1 $T=46980 1000 0 0 $X=46865 $Y=885
X12296 292 271 271 502 732 271 AND2_X1 $T=46980 43000 1 0 $X=46865 $Y=41485
X12297 510 459 271 502 472 271 AND2_X1 $T=49450 54200 0 180 $X=48575 $Y=52685
X12298 588 460 271 502 740 1265 AND2_X1 $T=49070 1000 0 0 $X=48955 $Y=885
X12299 510 469 271 502 1236 271 AND2_X1 $T=50970 37400 0 180 $X=50095 $Y=35885
X12300 510 471 271 502 1209 271 AND2_X1 $T=50590 51400 0 0 $X=50475 $Y=51285
X12301 1069 473 271 502 932 271 AND2_X1 $T=50780 17800 1 0 $X=50665 $Y=16285
X12302 510 475 271 502 747 271 AND2_X1 $T=50780 54200 1 0 $X=50665 $Y=52685
X12303 510 476 271 502 749 271 AND2_X1 $T=50970 48600 1 0 $X=50855 $Y=47085
X12304 510 480 271 502 1075 271 AND2_X1 $T=52110 37400 1 0 $X=51995 $Y=35885
X12305 510 481 271 502 936 271 AND2_X1 $T=52110 48600 0 0 $X=51995 $Y=48485
X12306 588 487 271 502 1149 271 AND2_X1 $T=54390 9400 0 180 $X=53515 $Y=7885
X12307 510 490 271 502 1211 271 AND2_X1 $T=54390 45800 1 180 $X=53515 $Y=45685
X12308 588 491 271 502 1212 1265 AND2_X1 $T=54770 1000 1 180 $X=53895 $Y=885
X12309 588 492 271 502 1151 271 AND2_X1 $T=54770 3800 1 180 $X=53895 $Y=3685
X12310 588 498 271 502 1239 271 AND2_X1 $T=56100 9400 0 180 $X=55225 $Y=7885
X12311 588 499 271 502 1152 271 AND2_X1 $T=56100 9400 1 180 $X=55225 $Y=9285
X12312 588 495 271 502 1079 271 AND2_X1 $T=55340 15000 1 0 $X=55225 $Y=13485
X12313 943 497 271 502 1080 271 AND2_X1 $T=55340 17800 0 0 $X=55225 $Y=17685
X12314 973 83 963 53 271 502 AOI21_X1 $T=10120 45800 0 0 $X=10005 $Y=45685
X12315 768 960 803 967 271 502 AOI21_X1 $T=10310 40200 1 0 $X=10195 $Y=38685
X12316 774 62 795 527 271 502 AOI21_X1 $T=10500 29000 1 0 $X=10385 $Y=27485
X12317 795 64 523 527 271 502 AOI21_X1 $T=10880 26200 0 0 $X=10765 $Y=26085
X12318 91 63 59 525 271 502 AOI21_X1 $T=11640 51400 0 180 $X=10765 $Y=49885
X12319 79 84 124 64 271 502 AOI21_X1 $T=13540 26200 0 0 $X=13425 $Y=26085
X12320 533 87 980 803 271 502 AOI21_X1 $T=13730 37400 0 0 $X=13615 $Y=37285
X12321 1110 95 553 984 271 502 AOI21_X1 $T=14300 31800 1 0 $X=14185 $Y=30285
X12322 974 117 1112 797 271 502 AOI21_X1 $T=17150 20600 1 180 $X=16275 $Y=20485
X12323 1107 126 558 554 271 502 AOI21_X1 $T=17340 34600 1 0 $X=17225 $Y=33085
X12324 117 138 1178 1117 271 502 AOI21_X1 $T=18100 29000 1 0 $X=17985 $Y=27485
X12325 574 146 1155 130 271 502 AOI21_X1 $T=19810 34600 0 180 $X=18935 $Y=33085
X12326 121 119 1117 208 271 502 AOI21_X1 $T=20000 26200 1 180 $X=19125 $Y=26085
X12327 572 121 217 994 271 502 AOI21_X1 $T=21900 17800 0 180 $X=21025 $Y=16285
X12328 196 188 824 1000 271 502 AOI21_X1 $T=23610 34600 1 180 $X=22735 $Y=34485
X12329 210 194 98 196 271 502 AOI21_X1 $T=23800 43000 1 180 $X=22925 $Y=42885
X12330 827 566 1184 221 271 502 AOI21_X1 $T=23800 29000 1 0 $X=23685 $Y=27485
X12331 586 209 580 1186 271 502 AOI21_X1 $T=24180 29000 0 0 $X=24065 $Y=28885
X12332 208 209 1186 252 271 502 AOI21_X1 $T=24560 29000 1 0 $X=24445 $Y=27485
X12333 196 215 830 1185 271 502 AOI21_X1 $T=25320 34600 0 180 $X=24445 $Y=33085
X12334 196 154 838 1233 271 502 AOI21_X1 $T=25320 34600 1 0 $X=25205 $Y=33085
X12335 202 236 232 1123 271 502 AOI21_X1 $T=26840 15000 1 0 $X=26725 $Y=13485
X12336 244 247 1216 1016 271 502 AOI21_X1 $T=27600 17800 0 0 $X=27485 $Y=17685
X12337 596 599 1005 283 271 502 AOI21_X1 $T=27980 43000 0 0 $X=27865 $Y=42885
X12338 847 456 1012 1021 271 502 AOI21_X1 $T=29690 45800 1 180 $X=28815 $Y=45685
X12339 196 265 845 1191 271 502 AOI21_X1 $T=30070 31800 0 180 $X=29195 $Y=30285
X12340 608 280 211 616 271 502 AOI21_X1 $T=30450 40200 1 0 $X=30335 $Y=38685
X12341 196 282 848 621 271 502 AOI21_X1 $T=30830 31800 1 0 $X=30715 $Y=30285
X12342 271 283 617 1023 271 502 AOI21_X1 $T=30830 45800 1 0 $X=30715 $Y=44285
X12343 361 281 874 615 271 502 AOI21_X1 $T=31780 17800 1 180 $X=30905 $Y=17685
X12344 361 605 286 611 271 502 AOI21_X1 $T=32160 20600 1 180 $X=31285 $Y=20485
X12345 196 301 625 856 271 502 AOI21_X1 $T=33300 31800 0 180 $X=32425 $Y=30285
X12346 290 303 631 221 271 502 AOI21_X1 $T=32920 17800 1 0 $X=32805 $Y=16285
X12347 866 321 1196 639 271 502 AOI21_X1 $T=33870 37400 1 0 $X=33755 $Y=35885
X12348 196 203 864 652 271 502 AOI21_X1 $T=34250 29000 0 0 $X=34135 $Y=28885
X12349 341 344 336 269 271 502 AOI21_X1 $T=35960 12200 0 0 $X=35845 $Y=12085
X12350 196 346 1026 1032 271 502 AOI21_X1 $T=37100 29000 1 180 $X=36225 $Y=28885
X12351 196 1035 892 878 271 502 AOI21_X1 $T=37480 23400 1 0 $X=37365 $Y=21885
X12352 894 367 1031 888 271 502 AOI21_X1 $T=38050 34600 0 0 $X=37935 $Y=34485
X12353 196 372 876 883 271 502 AOI21_X1 $T=38430 29000 0 0 $X=38315 $Y=28885
X12354 361 308 882 221 271 502 AOI21_X1 $T=38810 15000 1 0 $X=38695 $Y=13485
X12355 196 396 673 1200 271 502 AOI21_X1 $T=39760 26200 0 0 $X=39645 $Y=26085
X12356 196 404 1169 1235 271 502 AOI21_X1 $T=42230 26200 1 0 $X=42115 $Y=24685
X12357 705 412 1168 697 271 502 AOI21_X1 $T=44510 34600 1 180 $X=43635 $Y=34485
X12358 196 407 1051 1206 271 502 AOI21_X1 $T=44130 26200 0 0 $X=44015 $Y=26085
X12359 914 427 907 430 271 502 AOI21_X1 $T=45080 37400 1 0 $X=44965 $Y=35885
X12360 196 216 433 1222 271 502 AOI21_X1 $T=45460 26200 0 0 $X=45345 $Y=26085
X12361 403 433 910 717 271 502 AOI21_X1 $T=46410 31800 0 180 $X=45535 $Y=30285
X12362 725 718 1060 479 271 502 AOI21_X1 $T=47550 48600 1 180 $X=46675 $Y=48485
X12363 445 447 926 917 271 502 AOI21_X1 $T=47170 31800 1 0 $X=47055 $Y=30285
X12364 196 450 724 731 271 502 AOI21_X1 $T=48500 26200 1 180 $X=47625 $Y=26085
X12365 380 455 733 326 271 502 AOI21_X1 $T=48880 34600 1 180 $X=48005 $Y=34485
X12366 196 465 735 734 271 502 AOI21_X1 $T=50400 23400 1 180 $X=49525 $Y=23285
X12367 196 583 739 1145 271 502 AOI21_X1 $T=50970 20600 1 180 $X=50095 $Y=20485
X12368 196 477 748 1210 271 502 AOI21_X1 $T=51160 17800 0 0 $X=51045 $Y=17685
X12369 196 442 928 930 271 502 AOI21_X1 $T=52300 15000 1 180 $X=51425 $Y=14885
X12370 196 482 938 1078 271 502 AOI21_X1 $T=54010 15000 0 180 $X=53135 $Y=13485
X12371 196 493 751 946 271 502 AOI21_X1 $T=55150 20600 1 180 $X=54275 $Y=20485
X12372 196 496 1083 942 271 502 AOI21_X1 $T=56100 17800 0 180 $X=55225 $Y=16285
X12800 271 82 693 94 502 XNOR2_X1 $T=14110 40200 0 0 $X=13995 $Y=40085
X12801 271 1115 555 131 502 XNOR2_X1 $T=17530 43000 0 0 $X=17415 $Y=42885
X12802 271 831 283 220 502 XNOR2_X1 $T=25890 37400 1 180 $X=24635 $Y=37285
X12803 271 1010 250 230 502 XNOR2_X1 $T=26270 37400 0 0 $X=26155 $Y=37285
X12804 271 1126 639 294 502 XNOR2_X1 $T=31590 37400 1 0 $X=31475 $Y=35885
X12805 271 645 653 1128 502 XNOR2_X1 $T=33110 34600 0 0 $X=32995 $Y=34485
X12806 271 867 668 353 502 XNOR2_X1 $T=36530 29000 1 0 $X=36415 $Y=27485
X12807 271 676 1167 886 502 XNOR2_X1 $T=38620 26200 0 0 $X=38505 $Y=26085
X12808 271 1037 888 881 502 XNOR2_X1 $T=40710 34600 0 180 $X=39455 $Y=33085
X12809 271 1045 670 395 502 XNOR2_X1 $T=40710 34600 1 0 $X=40595 $Y=33085
X12810 271 906 365 698 502 XNOR2_X1 $T=44510 34600 0 180 $X=43255 $Y=33085
X12811 271 903 696 710 502 XNOR2_X1 $T=43750 20600 1 0 $X=43635 $Y=19085
X12812 271 717 326 429 502 XNOR2_X1 $T=45270 34600 0 0 $X=45155 $Y=34485
X12813 271 403 429 433 502 XNOR2_X1 $T=46790 34600 0 180 $X=45535 $Y=33085
X12814 271 746 697 736 502 XNOR2_X1 $T=48310 34600 1 0 $X=48195 $Y=33085
X12815 271 1148 430 750 502 XNOR2_X1 $T=51350 29000 1 0 $X=51235 $Y=27485
X12816 271 1071 389 745 502 XNOR2_X1 $T=51540 31800 0 0 $X=51425 $Y=31685
X12817 271 947 680 1150 502 XNOR2_X1 $T=56100 31800 1 180 $X=54845 $Y=31685
X12818 502 771 72 523 271 XOR2_X1 $T=9740 23400 1 0 $X=9625 $Y=21885
X12819 502 1103 971 1217 271 XOR2_X1 $T=12590 43000 1 180 $X=11335 $Y=42885
X12820 502 96 526 532 271 XOR2_X1 $T=13350 23400 0 180 $X=12095 $Y=21885
X12821 502 89 96 789 271 XOR2_X1 $T=14490 29000 0 180 $X=13235 $Y=27485
X12822 502 64 1156 795 271 XOR2_X1 $T=14300 26200 0 0 $X=14185 $Y=26085
X12823 502 1110 55 800 271 XOR2_X1 $T=15440 29000 1 0 $X=15325 $Y=27485
X12824 502 103 598 800 271 XOR2_X1 $T=17720 29000 0 180 $X=16465 $Y=27485
X12825 502 793 806 567 271 XOR2_X1 $T=17530 45800 1 0 $X=17415 $Y=44285
X12826 502 1116 161 990 271 XOR2_X1 $T=19050 40200 1 0 $X=18935 $Y=38685
X12827 502 149 174 155 271 XOR2_X1 $T=20760 34600 1 0 $X=20645 $Y=33085
X12828 502 993 1180 818 271 XOR2_X1 $T=20760 45800 0 0 $X=20645 $Y=45685
X12829 502 580 1003 188 271 XOR2_X1 $T=22280 29000 0 0 $X=22165 $Y=28885
X12830 502 580 220 824 271 XOR2_X1 $T=22280 37400 1 0 $X=22165 $Y=35885
X12831 502 183 825 998 271 XOR2_X1 $T=23230 40200 1 0 $X=23115 $Y=38685
X12832 502 219 230 830 271 XOR2_X1 $T=24180 34600 0 0 $X=24065 $Y=34485
X12833 502 182 1218 195 271 XOR2_X1 $T=25320 31800 0 0 $X=25205 $Y=31685
X12834 502 171 1013 838 271 XOR2_X1 $T=26080 34600 1 0 $X=25965 $Y=33085
X12835 502 839 603 1013 271 XOR2_X1 $T=27600 37400 1 0 $X=27485 $Y=35885
X12836 502 262 295 846 271 XOR2_X1 $T=28740 37400 1 0 $X=28625 $Y=35885
X12837 502 258 1162 268 271 XOR2_X1 $T=30070 29000 0 0 $X=29955 $Y=28885
X12838 502 614 294 848 271 XOR2_X1 $T=31590 34600 0 180 $X=30335 $Y=33085
X12839 502 287 613 626 271 XOR2_X1 $T=32730 29000 0 180 $X=31475 $Y=27485
X12840 502 644 1128 625 271 XOR2_X1 $T=33110 31800 1 180 $X=31855 $Y=31685
X12841 502 309 651 345 271 XOR2_X1 $T=33870 29000 1 0 $X=33755 $Y=27485
X12842 502 316 863 864 271 XOR2_X1 $T=34440 31800 0 0 $X=34325 $Y=31685
X12843 502 1221 665 863 271 XOR2_X1 $T=36150 34600 0 180 $X=34895 $Y=33085
X12844 502 358 347 870 271 XOR2_X1 $T=37290 34600 0 180 $X=36035 $Y=33085
X12845 502 669 881 876 271 XOR2_X1 $T=39760 31800 0 180 $X=38505 $Y=30285
X12846 502 880 675 1140 271 XOR2_X1 $T=40330 20600 1 180 $X=39075 $Y=20485
X12847 502 1135 889 892 271 XOR2_X1 $T=39760 29000 0 0 $X=39645 $Y=28885
X12848 502 1135 1044 880 271 XOR2_X1 $T=39950 23400 1 0 $X=39835 $Y=21885
X12849 502 692 395 673 271 XOR2_X1 $T=40520 31800 0 0 $X=40405 $Y=31685
X12850 502 386 392 681 271 XOR2_X1 $T=41850 23400 1 180 $X=40595 $Y=23285
X12851 502 1138 317 889 271 XOR2_X1 $T=41660 31800 0 0 $X=41545 $Y=31685
X12852 502 923 359 1046 271 XOR2_X1 $T=42230 31800 1 0 $X=42115 $Y=30285
X12853 502 410 380 436 271 XOR2_X1 $T=43940 31800 1 180 $X=42685 $Y=31685
X12854 502 702 698 1051 271 XOR2_X1 $T=44510 29000 0 180 $X=43255 $Y=27485
X12855 502 432 905 436 271 XOR2_X1 $T=44130 26200 1 0 $X=44015 $Y=24685
X12856 502 421 729 724 271 XOR2_X1 $T=46790 29000 0 180 $X=45535 $Y=27485
X12857 502 452 919 1061 271 XOR2_X1 $T=47550 26200 1 0 $X=47435 $Y=24685
X12858 502 458 1068 920 271 XOR2_X1 $T=47740 20600 0 0 $X=47625 $Y=20485
X12859 502 461 1065 463 271 XOR2_X1 $T=47930 15000 1 0 $X=47815 $Y=13485
X12860 502 416 741 735 271 XOR2_X1 $T=48880 31800 0 0 $X=48765 $Y=31685
X12861 502 926 314 741 271 XOR2_X1 $T=50590 34600 0 180 $X=49335 $Y=33085
X12862 502 439 745 928 271 XOR2_X1 $T=50020 26200 1 0 $X=49905 $Y=24685
X12863 502 915 736 739 271 XOR2_X1 $T=51350 29000 0 180 $X=50095 $Y=27485
X12864 502 927 934 943 271 XOR2_X1 $T=50780 20600 1 0 $X=50665 $Y=19085
X12865 502 1073 750 748 271 XOR2_X1 $T=50780 23400 1 0 $X=50665 $Y=21885
X12866 502 929 937 1069 271 XOR2_X1 $T=52110 15000 1 0 $X=51995 $Y=13485
X12867 502 484 391 941 271 XOR2_X1 $T=54010 26200 1 180 $X=52755 $Y=26085
X12868 502 720 1150 751 271 XOR2_X1 $T=54770 29000 1 180 $X=53515 $Y=28885
X12869 502 451 752 488 271 XOR2_X1 $T=54200 17800 1 0 $X=54085 $Y=16285
X12870 502 1153 1081 1083 271 XOR2_X1 $T=54960 23400 1 0 $X=54845 $Y=21885
X12871 502 940 378 1081 271 XOR2_X1 $T=56100 29000 0 180 $X=54845 $Y=27485
X13340 155 149 151 271 502 813 OR3_X1 $T=19240 37400 1 0 $X=19125 $Y=35885
X13341 195 182 177 271 502 155 OR3_X1 $T=23230 31800 1 180 $X=22165 $Y=31685
X13342 268 258 254 271 502 195 OR3_X1 $T=29310 29000 1 180 $X=28245 $Y=28885
X13343 426 432 436 271 502 1061 OR3_X1 $T=45840 23400 1 0 $X=45725 $Y=21885
X13344 463 461 462 271 502 1069 OR3_X1 $T=49070 15000 1 0 $X=48955 $Y=13485
X13345 488 451 494 271 502 943 OR3_X1 $T=54390 17800 0 0 $X=54275 $Y=17685
X13534 113 60 531 514 271 502 OAI21_X1 $T=10500 12200 1 0 $X=10385 $Y=10685
X13535 113 61 515 777 271 502 OAI21_X1 $T=10500 12200 0 0 $X=10385 $Y=12085
X13536 512 958 788 536 271 502 OAI21_X1 $T=11070 26200 1 0 $X=10955 $Y=24685
X13537 969 770 69 536 271 502 OAI21_X1 $T=12020 23400 0 0 $X=11905 $Y=23285
X13538 535 76 974 1242 271 502 OAI21_X1 $T=12780 20600 1 0 $X=12665 $Y=19085
X13539 539 70 66 782 271 502 OAI21_X1 $T=13540 48600 0 180 $X=12665 $Y=47085
X13540 1155 82 56 784 271 502 OAI21_X1 $T=13350 40200 0 0 $X=13235 $Y=40085
X13541 789 89 103 93 271 502 OAI21_X1 $T=13920 29000 0 0 $X=13805 $Y=28885
X13542 788 96 607 93 271 502 OAI21_X1 $T=15250 23400 1 180 $X=14375 $Y=23285
X13543 113 99 104 65 271 502 OAI21_X1 $T=14680 12200 0 0 $X=14565 $Y=12085
X13544 790 101 800 95 271 502 OAI21_X1 $T=14680 31800 0 0 $X=14565 $Y=31685
X13545 984 103 160 95 271 502 OAI21_X1 $T=15820 31800 0 180 $X=14945 $Y=30285
X13546 560 123 100 799 271 502 OAI21_X1 $T=17910 9400 0 180 $X=17035 $Y=7885
X13547 560 132 129 988 271 502 OAI21_X1 $T=17910 9400 1 0 $X=17795 $Y=7885
X13548 194 134 808 804 271 502 OAI21_X1 $T=18860 51400 1 180 $X=17985 $Y=51285
X13549 560 143 557 1113 271 502 OAI21_X1 $T=19430 17800 0 180 $X=18555 $Y=16285
X13550 987 145 209 562 271 502 OAI21_X1 $T=18860 31800 1 0 $X=18745 $Y=30285
X13551 149 155 162 151 271 502 OAI21_X1 $T=19430 34600 0 0 $X=19315 $Y=34485
X13552 545 121 192 565 271 502 OAI21_X1 $T=19810 17800 1 0 $X=19695 $Y=16285
X13553 558 160 223 169 271 502 OAI21_X1 $T=19810 31800 0 0 $X=19695 $Y=31685
X13554 821 146 998 999 271 502 OAI21_X1 $T=21710 40200 1 0 $X=21595 $Y=38685
X13555 210 178 1002 1001 271 502 OAI21_X1 $T=22280 51400 1 0 $X=22165 $Y=49885
X13556 998 183 990 999 271 502 OAI21_X1 $T=22470 40200 1 0 $X=22355 $Y=38685
X13557 182 195 193 177 271 502 OAI21_X1 $T=23990 31800 1 180 $X=23115 $Y=31685
X13558 845 261 846 841 271 502 OAI21_X1 $T=29690 31800 1 180 $X=28815 $Y=31685
X13559 846 262 839 841 271 502 OAI21_X1 $T=29880 34600 1 180 $X=29005 $Y=34485
X13560 258 268 255 254 271 502 OAI21_X1 $T=29310 29000 0 0 $X=29195 $Y=28885
X13561 260 270 351 1018 271 502 OAI21_X1 $T=30640 9400 0 180 $X=29765 $Y=7885
X13562 319 276 661 850 271 502 OAI21_X1 $T=31210 6600 1 180 $X=30335 $Y=6485
X13563 619 234 313 612 271 502 OAI21_X1 $T=31400 23400 1 180 $X=30525 $Y=23285
X13564 1196 295 596 855 271 502 OAI21_X1 $T=32540 37400 1 180 $X=31665 $Y=37285
X13565 319 298 312 633 271 502 OAI21_X1 $T=32160 6600 0 0 $X=32045 $Y=6485
X13566 632 305 1023 641 271 502 OAI21_X1 $T=32730 45800 1 0 $X=32615 $Y=44285
X13567 648 305 859 649 271 502 OAI21_X1 $T=34250 45800 0 180 $X=33375 $Y=44285
X13568 657 339 1040 865 271 502 OAI21_X1 $T=35390 45800 0 0 $X=35275 $Y=45685
X13569 869 305 659 664 271 502 OAI21_X1 $T=36910 43000 1 180 $X=36035 $Y=42885
X13570 1031 347 866 1027 271 502 OAI21_X1 $T=37100 37400 0 180 $X=36225 $Y=35885
X13571 655 269 369 874 271 502 OAI21_X1 $T=36720 17800 0 0 $X=36605 $Y=17685
X13572 870 358 1221 875 271 502 OAI21_X1 $T=36910 31800 0 0 $X=36795 $Y=31685
X13573 877 363 608 674 271 502 OAI21_X1 $T=37670 37400 0 0 $X=37555 $Y=37285
X13574 1132 339 685 677 271 502 OAI21_X1 $T=38240 45800 1 0 $X=38125 $Y=44285
X13575 871 339 890 678 271 502 OAI21_X1 $T=38430 45800 0 0 $X=38315 $Y=45685
X13576 869 339 1024 1038 271 502 OAI21_X1 $T=39000 45800 1 0 $X=38885 $Y=44285
X13577 209 387 702 1042 271 502 OAI21_X1 $T=39950 12200 1 0 $X=39835 $Y=10685
X13578 209 385 1135 885 271 502 OAI21_X1 $T=40710 17800 1 180 $X=39835 $Y=17685
X13579 1168 359 894 895 271 502 OAI21_X1 $T=41090 34600 0 0 $X=40975 $Y=34485
X13580 397 900 398 884 271 502 OAI21_X1 $T=41280 37400 1 0 $X=41165 $Y=35885
X13581 400 315 1047 271 271 502 OAI21_X1 $T=42040 45800 1 180 $X=41165 $Y=45685
X13582 1169 401 1046 897 271 502 OAI21_X1 $T=42040 26200 0 0 $X=41925 $Y=26085
X13583 405 315 1139 893 271 502 OAI21_X1 $T=42800 45800 1 180 $X=41925 $Y=45685
X13584 1046 923 1138 897 271 502 OAI21_X1 $T=42230 29000 1 0 $X=42115 $Y=27485
X13585 465 416 904 708 271 502 OAI21_X1 $T=43940 23400 0 0 $X=43825 $Y=23285
X13586 209 200 421 902 271 502 OAI21_X1 $T=44890 12200 0 180 $X=44015 $Y=10685
X13587 907 391 705 419 271 502 OAI21_X1 $T=45270 34600 1 180 $X=44395 $Y=34485
X13588 906 424 717 908 271 502 OAI21_X1 $T=44890 29000 0 0 $X=44775 $Y=28885
X13589 209 837 720 1141 271 502 OAI21_X1 $T=45650 12200 0 0 $X=45535 $Y=12085
X13590 436 432 1207 426 271 502 OAI21_X1 $T=46410 23400 1 180 $X=45535 $Y=23285
X13591 403 433 445 911 271 502 OAI21_X1 $T=47170 31800 0 180 $X=46295 $Y=30285
X13592 733 393 914 913 271 502 OAI21_X1 $T=48120 34600 1 180 $X=47245 $Y=34485
X13593 1054 292 743 1062 271 502 OAI21_X1 $T=47360 40200 1 0 $X=47245 $Y=38685
X13594 461 463 473 462 271 502 OAI21_X1 $T=49070 15000 0 0 $X=48955 $Y=14885
X13595 1066 263 471 922 271 502 OAI21_X1 $T=49450 51400 1 0 $X=49335 $Y=49885
X13596 474 263 489 1074 271 502 OAI21_X1 $T=51540 45800 1 0 $X=51425 $Y=44285
X13597 941 484 940 939 271 502 OAI21_X1 $T=53440 26200 1 0 $X=53325 $Y=24685
X13598 451 488 497 494 271 502 OAI21_X1 $T=53630 17800 0 0 $X=53515 $Y=17685
X13599 938 483 941 939 271 502 OAI21_X1 $T=54390 20600 1 180 $X=53515 $Y=20485
X13649 271 502 500 6 503 ICV_27 $T=1000 20600 1 0 $X=885 $Y=19085
X13650 271 502 500 7 1089 ICV_27 $T=1000 26200 1 0 $X=885 $Y=24685
X13651 271 502 500 8 951 ICV_27 $T=1000 29000 0 0 $X=885 $Y=28885
X13652 271 502 510 46 1173 ICV_27 $T=6510 51400 0 0 $X=6395 $Y=51285
X13653 271 502 500 52 521 ICV_27 $T=9550 3800 1 0 $X=9435 $Y=2285
X13654 271 502 510 56 1175 ICV_27 $T=10120 43000 0 0 $X=10005 $Y=42885
X13655 271 502 209 223 253 ICV_27 $T=26080 29000 0 0 $X=25965 $Y=28885
X13656 271 502 208 253 304 ICV_27 $T=28360 26200 0 0 $X=28245 $Y=26085
X13657 271 502 588 464 1144 ICV_27 $T=49260 3800 1 0 $X=49145 $Y=2285
X13658 271 502 510 485 1213 ICV_27 $T=53440 37400 0 0 $X=53325 $Y=37285
X13659 271 502 510 486 1238 ICV_27 $T=53440 45800 1 0 $X=53325 $Y=44285
X13660 271 502 510 66 518 271 ICV_28 $T=10880 54200 1 0 $X=10765 $Y=52685
X13661 271 502 510 80 786 271 ICV_28 $T=12970 54200 1 0 $X=12855 $Y=52685
X13662 271 502 546 98 962 271 ICV_28 $T=14300 48600 1 0 $X=14185 $Y=47085
X13663 271 502 510 135 1176 271 ICV_28 $T=17720 54200 0 0 $X=17605 $Y=54085
X13664 271 502 588 199 1119 1265 ICV_28 $T=23610 1000 0 0 $X=23495 $Y=885
X13665 271 502 588 257 1189 1265 ICV_28 $T=28360 1000 0 0 $X=28245 $Y=885
X13666 271 502 588 383 1199 1265 ICV_28 $T=39570 1000 0 0 $X=39455 $Y=885
X13667 271 502 510 413 1205 271 ICV_28 $T=43370 51400 0 0 $X=43255 $Y=51285
X13668 271 502 510 489 1237 271 ICV_28 $T=53440 43000 1 0 $X=53325 $Y=41485
X13745 1226 15 271 502 207 1265 DFF_X1 $T=1000 1000 0 0 $X=885 $Y=885
X13746 1172 23 271 502 760 271 DFF_X1 $T=1000 45800 0 0 $X=885 $Y=45685
X13747 1227 23 271 502 501 271 DFF_X1 $T=4230 51400 0 180 $X=885 $Y=49885
X13748 948 15 271 502 92 271 DFF_X1 $T=1760 3800 0 0 $X=1645 $Y=3685
X13749 1087 15 271 502 112 271 DFF_X1 $T=2330 12200 1 0 $X=2215 $Y=10685
X13750 1088 15 271 502 119 271 DFF_X1 $T=2330 17800 1 0 $X=2215 $Y=16285
X13751 1089 15 271 502 958 271 DFF_X1 $T=2330 26200 1 0 $X=2215 $Y=24685
X13752 951 15 271 502 959 271 DFF_X1 $T=2330 31800 1 0 $X=2215 $Y=30285
X13753 1173 24 271 502 1231 271 DFF_X1 $T=2330 54200 1 0 $X=2215 $Y=52685
X13754 1098 24 271 502 508 271 DFF_X1 $T=2330 57000 1 0 $X=2215 $Y=55485
X13755 1228 15 271 502 89 271 DFF_X1 $T=2710 26200 0 0 $X=2595 $Y=26085
X13756 1100 15 271 502 74 271 DFF_X1 $T=3090 3800 1 0 $X=2975 $Y=2285
X13757 953 15 271 502 764 271 DFF_X1 $T=3090 6600 0 0 $X=2975 $Y=6485
X13758 954 38 271 502 765 271 DFF_X1 $T=3090 23400 0 0 $X=2975 $Y=23285
X13759 1095 38 271 502 62 271 DFF_X1 $T=3090 29000 1 0 $X=2975 $Y=27485
X13760 1093 38 271 502 513 271 DFF_X1 $T=3090 43000 1 0 $X=2975 $Y=41485
X13761 952 38 271 502 768 271 DFF_X1 $T=3280 40200 0 0 $X=3165 $Y=40085
X13762 1094 15 271 502 106 271 DFF_X1 $T=3850 15000 0 0 $X=3735 $Y=14885
X13763 957 15 271 502 224 271 DFF_X1 $T=4420 12200 0 0 $X=4305 $Y=12085
X13764 950 15 271 502 204 271 DFF_X1 $T=4610 9400 0 0 $X=4495 $Y=9285
X13765 761 38 271 502 252 271 DFF_X1 $T=4990 20600 1 0 $X=4875 $Y=19085
X13766 1171 15 271 502 772 271 DFF_X1 $T=5560 31800 1 0 $X=5445 $Y=30285
X13767 1096 15 271 502 577 271 DFF_X1 $T=5750 17800 0 0 $X=5635 $Y=17685
X13768 505 15 271 502 87 271 DFF_X1 $T=5750 37400 1 0 $X=5635 $Y=35885
X13769 1175 24 271 502 769 271 DFF_X1 $T=5750 45800 1 0 $X=5635 $Y=44285
X13770 45 38 271 502 79 271 DFF_X1 $T=5940 26200 0 0 $X=5825 $Y=26085
X13771 1099 15 271 502 81 271 DFF_X1 $T=8980 3800 0 0 $X=8865 $Y=3685
X13772 1092 38 271 502 541 271 DFF_X1 $T=8980 37400 1 0 $X=8865 $Y=35885
X13773 956 38 271 502 1104 271 DFF_X1 $T=10500 43000 1 0 $X=10385 $Y=41485
X13774 1105 15 271 502 185 271 DFF_X1 $T=15440 3800 1 180 $X=12095 $Y=3685
X13775 1176 24 271 502 983 271 DFF_X1 $T=18670 57000 0 180 $X=15325 $Y=55485
X13776 551 15 271 502 201 271 DFF_X1 $T=16770 6600 0 0 $X=16655 $Y=6485
X13777 792 15 271 502 995 1265 DFF_X1 $T=17720 1000 0 0 $X=17605 $Y=885
X13778 148 24 271 502 1181 271 DFF_X1 $T=18670 57000 1 0 $X=18555 $Y=55485
X13779 1119 38 271 502 368 271 DFF_X1 $T=25510 3800 1 180 $X=22165 $Y=3685
X13780 272 24 271 502 1194 271 DFF_X1 $T=29310 54200 1 0 $X=29195 $Y=52685
X13781 1189 38 271 502 620 271 DFF_X1 $T=30450 3800 0 0 $X=30335 $Y=3685
X13782 1193 38 271 502 247 271 DFF_X1 $T=32160 3800 1 0 $X=32045 $Y=2285
X13783 1195 24 271 502 1197 271 DFF_X1 $T=32540 54200 1 0 $X=32425 $Y=52685
X13784 1129 38 271 502 371 271 DFF_X1 $T=33680 3800 0 0 $X=33565 $Y=3685
X13785 872 38 271 502 356 271 DFF_X1 $T=38620 3800 0 180 $X=35275 $Y=2285
X13786 1199 38 271 502 683 271 DFF_X1 $T=38620 3800 1 0 $X=38505 $Y=2285
X13787 376 38 271 502 366 271 DFF_X1 $T=38620 6600 1 0 $X=38505 $Y=5085
X13788 1198 24 271 502 1202 271 DFF_X1 $T=38620 54200 1 0 $X=38505 $Y=52685
X13789 1131 24 271 502 1203 271 DFF_X1 $T=38620 57000 1 0 $X=38505 $Y=55485
X13790 1234 38 271 502 679 1265 DFF_X1 $T=41280 1000 0 0 $X=41165 $Y=885
X13791 1204 38 271 502 274 271 DFF_X1 $T=42230 6600 1 0 $X=42115 $Y=5085
X13792 1205 24 271 502 1056 271 DFF_X1 $T=42230 57000 1 0 $X=42115 $Y=55485
X13793 417 24 271 502 1059 271 DFF_X1 $T=43560 54200 0 0 $X=43445 $Y=54085
X13794 709 38 271 502 243 271 DFF_X1 $T=43750 3800 0 0 $X=43635 $Y=3685
X13795 1208 38 271 502 335 271 DFF_X1 $T=49640 6600 0 0 $X=49525 $Y=6485
X13796 472 24 271 502 1076 271 DFF_X1 $T=50020 57000 1 0 $X=49905 $Y=55485
X13797 1149 38 271 502 344 271 DFF_X1 $T=53630 9400 0 180 $X=50285 $Y=7885
X13798 740 38 271 502 285 1265 DFF_X1 $T=50780 1000 0 0 $X=50665 $Y=885
X13799 1144 38 271 502 423 271 DFF_X1 $T=50780 3800 0 0 $X=50665 $Y=3685
X13800 1152 38 271 502 377 271 DFF_X1 $T=55340 9400 1 180 $X=51995 $Y=9285
X13801 1212 38 271 502 242 271 DFF_X1 $T=52870 3800 1 0 $X=52755 $Y=2285
X13802 1239 38 271 502 190 271 DFF_X1 $T=56100 6600 1 180 $X=52755 $Y=6485
X13803 1075 24 271 502 944 271 DFF_X1 $T=52870 37400 1 0 $X=52755 $Y=35885
X13804 1237 24 271 502 753 271 DFF_X1 $T=52870 40200 0 0 $X=52755 $Y=40085
X13805 1211 24 271 502 945 271 DFF_X1 $T=52870 48600 0 0 $X=52755 $Y=48485
X13806 936 24 271 502 1082 271 DFF_X1 $T=52870 51400 0 0 $X=52755 $Y=51285
X13807 1151 38 271 502 453 271 DFF_X1 $T=53250 6600 1 0 $X=53135 $Y=5085
X13808 1079 38 271 502 308 271 DFF_X1 $T=53250 12200 1 0 $X=53135 $Y=10685
X13809 1238 24 271 502 755 271 DFF_X1 $T=53250 43000 0 0 $X=53135 $Y=42885
X13810 749 24 271 502 756 271 DFF_X1 $T=53250 48600 1 0 $X=53135 $Y=47085
X13811 1209 24 271 502 757 271 DFF_X1 $T=53250 54200 1 0 $X=53135 $Y=52685
X13812 747 24 271 502 1085 271 DFF_X1 $T=53250 57000 1 0 $X=53135 $Y=55485
X13848 271 502 1091 15 225 271 ICV_34 $T=3280 15000 1 0 $X=3165 $Y=13485
X13849 271 502 1229 38 965 271 ICV_34 $T=5750 31800 0 0 $X=5635 $Y=31685
X13850 271 502 509 38 975 271 ICV_34 $T=8790 34600 0 0 $X=8675 $Y=34485
X13851 271 502 968 15 205 1265 ICV_34 $T=11450 1000 0 0 $X=11335 $Y=885
X13852 271 502 1130 24 1036 271 ICV_34 $T=35200 57000 1 0 $X=35085 $Y=55485
X13853 271 502 1133 24 899 271 ICV_34 $T=40140 54200 0 0 $X=40025 $Y=54085
X13854 271 502 1236 24 1084 271 ICV_34 $T=53060 34600 1 0 $X=52945 $Y=33085
X13855 271 502 1213 24 754 271 ICV_34 $T=53060 40200 1 0 $X=52945 $Y=38685
X13856 91 271 766 964 502 NAND2_X1 $T=8600 48600 1 180 $X=7915 $Y=48485
X13857 55 271 67 529 502 NAND2_X1 $T=9740 20600 1 0 $X=9625 $Y=19085
X13858 524 271 83 767 502 NAND2_X1 $T=10500 48600 0 180 $X=9815 $Y=47085
X13859 55 271 526 113 502 NAND2_X1 $T=10310 20600 1 0 $X=10195 $Y=19085
X13860 55 271 179 68 502 NAND2_X1 $T=10500 17800 0 0 $X=10385 $Y=17685
X13861 969 271 770 536 502 NAND2_X1 $T=11830 26200 1 0 $X=11715 $Y=24685
X13862 1155 271 94 784 502 NAND2_X1 $T=12780 40200 0 0 $X=12665 $Y=40085
X13863 75 271 106 1242 502 NAND2_X1 $T=14110 20600 0 180 $X=13425 $Y=19085
X13864 788 271 96 93 502 NAND2_X1 $T=13920 23400 0 0 $X=13805 $Y=23285
X13865 790 271 101 95 502 NAND2_X1 $T=14110 31800 0 0 $X=13995 $Y=31685
X13866 986 271 980 796 502 NAND2_X1 $T=16200 37400 0 0 $X=16085 $Y=37285
X13867 118 271 207 799 502 NAND2_X1 $T=16580 9400 1 0 $X=16465 $Y=7885
X13868 986 271 803 126 502 NAND2_X1 $T=17150 37400 0 0 $X=17035 $Y=37285
X13869 194 271 134 804 502 NAND2_X1 $T=17530 51400 0 0 $X=17415 $Y=51285
X13870 75 271 128 988 502 NAND2_X1 $T=19240 9400 0 180 $X=18555 $Y=7885
X13871 109 271 121 159 502 NAND2_X1 $T=18860 23400 0 0 $X=18745 $Y=23285
X13872 557 271 121 565 502 NAND2_X1 $T=19430 17800 0 0 $X=19315 $Y=17685
X13873 821 271 146 999 502 NAND2_X1 $T=22850 37400 1 180 $X=22165 $Y=37285
X13874 98 271 90 263 502 NAND2_X1 $T=23040 45800 0 0 $X=22925 $Y=45685
X13875 210 271 178 1001 502 NAND2_X1 $T=23610 51400 0 180 $X=22925 $Y=49885
X13876 1005 271 823 1183 502 NAND2_X1 $T=24180 45800 1 180 $X=23495 $Y=45685
X13877 1012 271 590 229 502 NAND2_X1 $T=26650 48600 1 0 $X=26535 $Y=47085
X13878 256 271 1017 251 502 NAND2_X1 $T=27790 48600 0 0 $X=27675 $Y=48485
X13879 845 271 261 841 502 NAND2_X1 $T=28930 34600 1 0 $X=28815 $Y=33085
X13880 361 271 371 1018 502 NAND2_X1 $T=31210 9400 0 180 $X=30525 $Y=7885
X13881 281 271 328 612 502 NAND2_X1 $T=30640 23400 1 0 $X=30525 $Y=21885
X13882 361 271 221 619 502 NAND2_X1 $T=31780 23400 0 180 $X=31095 $Y=21885
X13883 278 271 290 260 502 NAND2_X1 $T=31970 15000 1 0 $X=31855 $Y=13485
X13884 290 271 1008 300 502 NAND2_X1 $T=32350 17800 1 0 $X=32235 $Y=16285
X13885 638 271 356 1022 502 NAND2_X1 $T=33110 12200 1 180 $X=32425 $Y=12085
X13886 322 271 670 637 502 NAND2_X1 $T=35200 40200 1 180 $X=34515 $Y=40085
X13887 1165 271 353 345 502 NAND2_X1 $T=36910 26200 1 180 $X=36225 $Y=26085
X13888 479 271 665 354 502 NAND2_X1 $T=36530 48600 0 0 $X=36415 $Y=48485
X13889 667 271 269 1025 502 NAND2_X1 $T=37670 17800 0 180 $X=36985 $Y=16285
X13890 884 271 373 877 502 NAND2_X1 $T=39760 37400 1 180 $X=39075 $Y=37285
X13891 890 271 315 893 502 NAND2_X1 $T=40710 45800 0 0 $X=40595 $Y=45685
X13892 1169 271 401 897 502 NAND2_X1 $T=43370 26200 1 180 $X=42685 $Y=26085
X13893 1052 271 1053 413 502 NAND2_X1 $T=43750 51400 1 0 $X=43635 $Y=49885
X13894 703 271 710 1140 502 NAND2_X1 $T=44320 20600 0 0 $X=44205 $Y=20485
X13895 407 271 702 708 502 NAND2_X1 $T=44320 23400 1 0 $X=44205 $Y=21885
X13896 1055 271 707 431 502 NAND2_X1 $T=45460 51400 0 180 $X=44775 $Y=49885
X13897 1051 271 702 908 502 NAND2_X1 $T=45080 29000 1 0 $X=44965 $Y=27485
X13898 420 271 1057 437 502 NAND2_X1 $T=45840 48600 1 0 $X=45725 $Y=47085
X13899 912 271 1058 459 502 NAND2_X1 $T=46980 48600 0 180 $X=46295 $Y=47085
X13900 724 271 421 447 502 NAND2_X1 $T=48310 29000 0 180 $X=47625 $Y=27485
X13901 725 271 365 466 502 NAND2_X1 $T=47930 48600 1 0 $X=47815 $Y=47085
X13902 1063 271 737 480 502 NAND2_X1 $T=48500 37400 1 0 $X=48385 $Y=35885
X13903 732 271 393 921 502 NAND2_X1 $T=48690 40200 0 0 $X=48575 $Y=40085
X13904 1224 271 738 481 502 NAND2_X1 $T=48690 45800 1 0 $X=48575 $Y=44285
X13905 933 271 744 490 502 NAND2_X1 $T=51540 43000 1 180 $X=50855 $Y=42885
X13906 1070 271 1072 485 502 NAND2_X1 $T=51350 40200 1 0 $X=51235 $Y=38685
X13907 938 271 483 939 502 NAND2_X1 $T=53060 20600 0 0 $X=52945 $Y=20485
X14045 49 271 502 517 ICV_39 $T=11260 45800 0 180 $X=10765 $Y=44285
X14046 113 271 502 522 ICV_39 $T=11640 15000 0 180 $X=11145 $Y=13485
X14047 559 271 502 135 ICV_39 $T=19050 54200 0 180 $X=18555 $Y=52685
X14048 860 271 502 847 ICV_39 $T=30070 45800 1 180 $X=29575 $Y=45685
X14049 645 271 502 1127 ICV_39 $T=33870 34600 0 180 $X=33375 $Y=33085
X14050 653 271 502 321 ICV_39 $T=35010 37400 0 180 $X=34515 $Y=35885
X14051 1045 271 502 1134 ICV_39 $T=41090 31800 0 180 $X=40595 $Y=30285
X14052 414 271 502 436 ICV_39 $T=45270 15000 1 180 $X=44775 $Y=14885
X14053 730 271 502 439 ICV_39 $T=47930 15000 1 180 $X=47435 $Y=14885
X14054 1148 271 502 935 ICV_39 $T=52680 26200 0 180 $X=52185 $Y=24685
X14055 507 22 271 502 30 OR2_X1 $T=2330 43000 0 0 $X=2215 $Y=42885
X14056 507 22 271 502 47 OR2_X1 $T=5750 48600 1 180 $X=4875 $Y=48485
X14057 507 22 271 502 610 OR2_X1 $T=5940 48600 0 180 $X=5065 $Y=47085
X14058 626 287 271 502 268 OR2_X1 $T=31970 29000 1 180 $X=31095 $Y=28885
X14059 345 309 271 502 626 OR2_X1 $T=33870 29000 0 180 $X=32995 $Y=27485
X14060 69 331 271 502 655 OR2_X1 $T=34630 15000 1 0 $X=34515 $Y=13485
X14061 1140 880 271 502 681 OR2_X1 $T=39190 23400 1 0 $X=39075 $Y=21885
X14062 430 389 271 502 397 OR2_X1 $T=40330 34600 0 0 $X=40215 $Y=34485
X14063 1061 452 271 502 920 OR2_X1 $T=47930 23400 0 0 $X=47815 $Y=23285
X14064 920 458 271 502 463 OR2_X1 $T=48690 20600 1 0 $X=48575 $Y=19085
X14065 1069 929 271 502 488 OR2_X1 $T=52300 15000 0 0 $X=52185 $Y=14885
X14159 531 72 502 74 75 142 271 204 571 AOI222_X1 $T=12210 12200 1 0 $X=12095 $Y=10685
X14160 515 72 502 81 75 142 271 112 538 AOI222_X1 $T=13160 12200 0 0 $X=13045 $Y=12085
X14161 971 83 502 86 53 91 271 540 1154 AOI222_X1 $T=13350 48600 0 0 $X=13235 $Y=48485
X14162 791 83 502 108 53 91 271 552 982 AOI222_X1 $T=15250 45800 0 0 $X=15135 $Y=45685
X14163 104 72 502 207 75 142 271 224 127 AOI222_X1 $T=15440 12200 0 0 $X=15325 $Y=12085
X14164 555 83 502 116 53 91 271 1111 966 AOI222_X1 $T=17150 48600 1 180 $X=15515 $Y=48485
X14165 75 112 502 577 109 118 271 119 152 AOI222_X1 $T=15820 20600 1 0 $X=15705 $Y=19085
X14166 118 225 502 128 109 75 271 204 572 AOI222_X1 $T=17340 20600 1 0 $X=17225 $Y=19085
X14167 806 83 502 141 53 91 271 563 991 AOI222_X1 $T=18100 48600 1 0 $X=17985 $Y=47085
X14168 1180 83 502 144 53 91 271 814 559 AOI222_X1 $T=18290 51400 1 0 $X=18175 $Y=49885
X14169 1159 164 502 166 151 170 271 191 482 AOI222_X1 $T=20380 15000 1 0 $X=20265 $Y=13485
X14170 176 191 502 164 170 151 271 995 477 AOI222_X1 $T=23610 15000 1 180 $X=21975 $Y=14885
X14171 213 191 502 185 151 176 271 164 442 AOI222_X1 $T=23800 12200 1 180 $X=22165 $Y=12085
X14172 1182 164 502 92 151 192 271 191 404 AOI222_X1 $T=22280 17800 0 0 $X=22165 $Y=17685
X14173 1182 191 502 128 151 1179 271 164 1035 AOI222_X1 $T=22280 20600 1 0 $X=22165 $Y=19085
X14174 271 191 502 164 186 151 271 577 372 AOI222_X1 $T=22280 20600 0 0 $X=22165 $Y=20485
X14175 573 164 502 179 151 186 271 191 346 AOI222_X1 $T=22280 23400 1 0 $X=22165 $Y=21885
X14176 153 191 502 180 164 151 271 112 282 AOI222_X1 $T=22280 23400 0 0 $X=22165 $Y=23285
X14177 1159 191 502 74 151 206 271 164 496 AOI222_X1 $T=23610 15000 0 0 $X=23495 $Y=14885
X14178 579 191 502 201 151 213 271 164 465 AOI222_X1 $T=23800 12200 0 0 $X=23685 $Y=12085
X14179 217 191 502 81 151 192 271 164 583 AOI222_X1 $T=23800 17800 0 0 $X=23685 $Y=17685
X14180 1179 191 502 202 151 271 271 164 396 AOI222_X1 $T=23800 20600 1 0 $X=23685 $Y=19085
X14181 573 191 502 204 151 214 271 164 203 AOI222_X1 $T=23800 23400 1 0 $X=23685 $Y=21885
X14182 206 191 502 207 151 217 271 164 493 AOI222_X1 $T=23990 17800 1 0 $X=23875 $Y=16285
X14183 215 219 502 594 182 177 271 1011 826 AOI222_X1 $T=24940 31800 1 0 $X=24825 $Y=30285
X14184 153 164 502 224 151 214 271 191 301 AOI222_X1 $T=25320 23400 0 0 $X=25205 $Y=23285
X14185 362 620 502 285 278 293 271 252 622 AOI222_X1 $T=31020 9400 0 0 $X=30905 $Y=9285
X14186 1163 304 502 308 146 313 271 357 854 AOI222_X1 $T=32920 23400 1 0 $X=32805 $Y=21885
X14187 462 320 502 316 203 301 271 644 279 AOI222_X1 $T=34820 26200 0 180 $X=33185 $Y=24685
X14188 629 314 502 317 322 271 271 603 649 AOI222_X1 $T=33490 40200 1 0 $X=33375 $Y=38685
X14189 370 697 502 326 323 318 271 639 632 AOI222_X1 $T=35200 43000 1 180 $X=33565 $Y=42885
X14190 312 69 502 683 328 330 271 243 658 AOI222_X1 $T=33870 6600 0 0 $X=33755 $Y=6485
X14191 313 304 502 247 146 333 271 357 627 AOI222_X1 $T=34440 23400 1 0 $X=34325 $Y=21885
X14192 361 247 502 303 330 328 271 366 686 AOI222_X1 $T=35580 15000 0 0 $X=35465 $Y=14885
X14193 1028 357 502 356 146 350 271 304 1220 AOI222_X1 $T=37860 20600 0 180 $X=36225 $Y=19085
X14194 333 304 502 344 146 350 271 357 654 AOI222_X1 $T=36340 20600 0 0 $X=36225 $Y=20485
X14195 629 393 502 359 322 271 271 295 664 AOI222_X1 $T=36720 40200 1 0 $X=36605 $Y=38685
X14196 661 290 502 247 355 361 271 679 896 AOI222_X1 $T=37100 6600 1 0 $X=36985 $Y=5085
X14197 361 356 502 300 362 328 271 274 691 AOI222_X1 $T=37290 15000 1 0 $X=37175 $Y=13485
X14198 318 653 502 365 323 370 271 680 647 AOI222_X1 $T=37670 40200 0 0 $X=37555 $Y=40085
X14199 1028 304 502 357 369 146 271 620 671 AOI222_X1 $T=37860 20600 1 0 $X=37745 $Y=19085
X14200 361 366 502 667 362 328 271 679 898 AOI222_X1 $T=38050 12200 1 0 $X=37935 $Y=10685
X14201 330 368 502 371 328 361 271 344 379 AOI222_X1 $T=38240 12200 0 0 $X=38125 $Y=12085
X14202 355 377 502 274 361 334 271 290 694 AOI222_X1 $T=39950 9400 1 180 $X=38315 $Y=9285
X14203 370 378 502 380 323 318 271 665 648 AOI222_X1 $T=39190 40200 0 0 $X=39075 $Y=40085
X14204 312 290 502 243 361 355 271 344 1050 AOI222_X1 $T=39380 6600 0 0 $X=39265 $Y=6485
X14205 364 391 502 393 322 271 271 359 400 AOI222_X1 $T=40330 43000 1 0 $X=40215 $Y=41485
X14206 1039 357 502 366 146 369 271 304 682 AOI222_X1 $T=40710 17800 0 0 $X=40595 $Y=17685
X14207 364 389 502 365 322 271 271 680 689 AOI222_X1 $T=42230 40200 1 180 $X=40595 $Y=40085
X14208 382 304 502 274 146 409 271 357 1048 AOI222_X1 $T=42230 15000 0 0 $X=42115 $Y=14885
X14209 364 314 502 380 322 271 271 378 699 AOI222_X1 $T=42230 40200 1 0 $X=42115 $Y=38685
X14210 364 430 502 326 322 271 271 697 405 AOI222_X1 $T=42230 43000 0 0 $X=42115 $Y=42885
X14211 690 357 502 304 411 146 271 242 706 AOI222_X1 $T=43180 9400 0 0 $X=43065 $Y=9285
X14212 701 357 502 304 409 146 271 335 1146 AOI222_X1 $T=44320 15000 1 0 $X=44205 $Y=13485
X14213 435 304 502 423 146 425 271 357 721 AOI222_X1 $T=44510 9400 1 0 $X=44395 $Y=7885
X14214 435 357 502 190 146 712 271 304 730 AOI222_X1 $T=46030 9400 1 0 $X=45915 $Y=7885
X14215 438 304 502 243 146 446 271 357 454 AOI222_X1 $T=46410 12200 0 0 $X=46295 $Y=12085
X14216 712 357 502 285 146 448 271 304 320 AOI222_X1 $T=46790 9400 0 0 $X=46675 $Y=9285
X14217 446 304 502 453 146 448 271 357 924 AOI222_X1 $T=47740 12200 1 0 $X=47625 $Y=10685
X14218 743 718 502 314 479 478 271 389 1074 AOI222_X1 $T=52870 40200 1 180 $X=51235 $Y=40085
X14291 553 802 271 130 133 502 987 801 OAI221_X1 $T=17720 31800 1 0 $X=17605 $Y=30285
X14292 423 60 271 175 99 502 190 189 OAI221_X1 $T=22280 6600 0 0 $X=22165 $Y=6485
X14293 1004 995 271 189 185 502 276 197 OAI221_X1 $T=23800 6600 0 180 $X=22545 $Y=5085
X14294 285 61 271 197 198 502 453 576 OAI221_X1 $T=23420 9400 1 0 $X=23305 $Y=7885
X14295 298 201 271 212 205 502 200 175 OAI221_X1 $T=25320 6600 0 180 $X=24065 $Y=5085
X14296 589 836 271 238 157 502 387 245 OAI221_X1 $T=27030 6600 0 0 $X=26915 $Y=6485
X14297 1007 840 271 245 242 502 1122 212 OAI221_X1 $T=28360 6600 0 180 $X=27105 $Y=5085
X14298 237 620 271 248 593 502 356 1219 OAI221_X1 $T=27980 15000 0 0 $X=27865 $Y=14885
X14299 81 602 271 249 92 502 277 1124 OAI221_X1 $T=28170 12200 1 0 $X=28055 $Y=10685
X14300 254 623 271 279 265 502 261 449 OAI221_X1 $T=30260 26200 1 0 $X=30145 $Y=24685
X14301 636 263 271 284 289 502 291 299 OAI221_X1 $T=31020 51400 1 0 $X=30905 $Y=49885
X14302 636 291 271 324 327 502 263 306 OAI221_X1 $T=33870 51400 0 0 $X=33755 $Y=51285
X14303 342 263 271 862 327 502 291 343 OAI221_X1 $T=35010 51400 0 0 $X=34895 $Y=51285
X14304 1041 263 271 374 375 502 291 381 OAI221_X1 $T=38620 51400 1 0 $X=38505 $Y=49885
X14305 216 403 271 406 407 502 702 688 OAI221_X1 $T=42420 23400 1 0 $X=42305 $Y=21885
X14306 436 418 271 415 414 502 410 700 OAI221_X1 $T=44890 15000 1 180 $X=43635 $Y=14885
X14307 466 263 271 467 468 502 291 476 OAI221_X1 $T=49830 48600 1 0 $X=49715 $Y=47085
X14308 468 263 271 470 474 502 291 486 OAI221_X1 $T=50400 45800 1 0 $X=50285 $Y=44285
X14320 512 528 271 770 958 765 502 OAI22_X1 $T=8600 26200 1 0 $X=8485 $Y=24685
X14321 523 771 271 532 528 765 502 OAI22_X1 $T=11070 23400 0 0 $X=10955 $Y=23285
X14322 537 72 271 543 76 73 502 OAI22_X1 $T=13160 15000 0 0 $X=13045 $Y=14885
X14323 76 224 271 544 762 72 502 OAI22_X1 $T=14680 20600 0 0 $X=14565 $Y=20485
X14324 543 121 271 170 117 809 502 OAI22_X1 $T=17910 15000 0 0 $X=17795 $Y=14885
X14325 811 121 271 153 187 159 502 OAI22_X1 $T=19430 23400 0 0 $X=19315 $Y=23285
X14326 121 187 271 815 566 117 502 OAI22_X1 $T=20000 26200 0 0 $X=19885 $Y=26085
X14327 566 252 271 820 303 138 502 OAI22_X1 $T=20950 26200 0 0 $X=20835 $Y=26085
X14328 818 817 271 131 305 144 502 OAI22_X1 $T=20950 43000 1 0 $X=20835 $Y=41485
X14329 820 822 271 574 234 119 502 OAI22_X1 $T=22280 26200 0 0 $X=22165 $Y=26085
X14330 832 123 271 238 568 683 502 OAI22_X1 $T=26080 6600 0 0 $X=25965 $Y=6485
X14331 221 227 271 281 267 269 502 OAI22_X1 $T=29120 20600 0 0 $X=29005 $Y=20485
X14332 260 836 271 338 290 622 502 OAI22_X1 $T=33110 9400 0 180 $X=32045 $Y=7885
X14333 634 290 271 857 69 622 502 OAI22_X1 $T=33490 9400 1 180 $X=32425 $Y=9285
X14334 657 305 271 635 339 632 502 OAI22_X1 $T=32540 45800 0 0 $X=32425 $Y=45685
X14335 858 292 271 860 315 659 502 OAI22_X1 $T=33490 45800 0 0 $X=33375 $Y=45685
X14336 329 315 271 289 292 659 502 OAI22_X1 $T=33680 48600 1 0 $X=33565 $Y=47085
X14337 352 269 271 1028 319 1025 502 OAI22_X1 $T=37100 17800 0 180 $X=36035 $Y=16285
X14338 871 305 271 660 339 648 502 OAI22_X1 $T=37100 45800 1 180 $X=36035 $Y=45685
X14339 896 269 271 435 221 694 502 OAI22_X1 $T=42230 6600 0 0 $X=42115 $Y=6485
X14340 666 221 271 712 269 687 502 OAI22_X1 $T=43180 9400 1 180 $X=42115 $Y=9285
X14341 689 315 271 714 292 400 502 OAI22_X1 $T=43180 45800 0 180 $X=42115 $Y=44285
X14342 699 315 271 901 292 405 502 OAI22_X1 $T=44130 45800 0 180 $X=43065 $Y=44285
X14343 689 292 271 434 315 422 502 OAI22_X1 $T=43750 43000 0 0 $X=43635 $Y=42885
X14344 428 315 271 713 292 699 502 OAI22_X1 $T=44510 40200 0 0 $X=44395 $Y=40085
X14345 1054 315 271 716 292 428 502 OAI22_X1 $T=44700 40200 1 0 $X=44585 $Y=38685
X14346 722 315 271 909 292 422 502 OAI22_X1 $T=46220 43000 0 180 $X=45155 $Y=41485
X14347 929 483 271 925 924 482 502 OAI22_X1 $T=50970 12200 1 180 $X=49905 $Y=12085
X14386 965 271 502 789 ICV_53 $T=12590 31800 1 0 $X=12475 $Y=30285
X14387 1109 271 502 985 ICV_53 $T=15440 17800 1 0 $X=15325 $Y=16285
X14388 282 271 502 258 ICV_53 $T=28550 29000 1 0 $X=28435 $Y=27485
X14389 842 271 502 616 ICV_53 $T=30260 37400 0 0 $X=30145 $Y=37285
X14390 301 271 502 287 ICV_53 $T=31970 26200 0 0 $X=31855 $Y=26085
X14391 627 271 502 644 ICV_53 $T=32540 26200 1 0 $X=32425 $Y=24685
X14392 372 271 502 676 ICV_53 $T=37860 26200 0 0 $X=37745 $Y=26085
X14393 742 271 502 475 ICV_53 $T=49830 51400 0 0 $X=49715 $Y=51285
X14413 151 959 502 62 564 130 271 151 89 965 71 130 ICV_55 $T=10690 31800 0 0 $X=10575 $Y=31685
X14414 543 121 502 117 213 127 271 127 121 117 136 549 ICV_55 $T=16960 12200 0 0 $X=16845 $Y=12085
X14415 158 121 502 117 176 538 271 538 121 117 579 571 ICV_55 $T=20000 12200 0 0 $X=19885 $Y=12085
X14416 479 250 502 456 256 843 271 843 718 603 259 479 ICV_55 $T=28360 48600 0 0 $X=28245 $Y=48485
X14417 1043 269 502 221 446 666 271 898 269 221 448 694 ICV_55 $T=42230 12200 1 0 $X=42115 $Y=10685
X14418 687 269 502 221 425 1050 271 411 357 304 902 425 ICV_55 $T=42610 9400 1 0 $X=42495 $Y=7885
X14419 434 718 502 680 1224 479 271 725 393 365 474 732 ICV_55 $T=46790 45800 1 0 $X=46675 $Y=44285
X14420 478 326 502 365 922 918 271 478 365 380 742 918 ICV_55 $T=48690 48600 0 0 $X=48575 $Y=48485
X14421 478 391 502 456 1170 916 271 916 718 430 1072 478 ICV_55 $T=49640 37400 0 0 $X=49525 $Y=37285
X14430 271 502 124 650 827 ICV_57 $T=23990 26200 1 0 $X=23875 $Y=24685
X14431 271 502 453 198 585 ICV_57 $T=24370 6600 0 0 $X=24255 $Y=6485
X14432 271 502 478 250 844 ICV_57 $T=28170 51400 1 0 $X=28055 $Y=49885
X14433 271 502 280 842 1014 ICV_57 $T=28550 37400 0 0 $X=28435 $Y=37285
X14434 271 502 253 124 604 ICV_57 $T=28740 23400 0 0 $X=28625 $Y=23285
X14435 271 502 638 607 662 ICV_57 $T=33300 12200 1 0 $X=33185 $Y=10685
X14436 271 502 479 888 887 ICV_57 $T=39950 48600 0 0 $X=39835 $Y=48485
X14437 271 502 685 315 271 ICV_57 $T=41090 48600 1 0 $X=40975 $Y=47085
X14438 271 502 436 410 906 ICV_57 $T=43750 31800 1 0 $X=43635 $Y=30285
X14439 271 502 725 380 1066 ICV_57 $T=47930 48600 0 0 $X=47815 $Y=48485
X14440 271 502 1225 1170 469 ICV_57 $T=49450 37400 1 0 $X=49335 $Y=35885
X14457 271 502 511 225 128 514 516 ICV_58 $T=9170 15000 1 0 $X=9055 $Y=13485
X14458 271 502 151 794 541 70 130 ICV_58 $T=15440 40200 1 0 $X=15325 $Y=38685
X14459 271 502 1108 117 121 168 549 ICV_58 $T=17150 12200 1 0 $X=17035 $Y=10685
X14460 271 502 141 315 292 567 564 ICV_58 $T=20760 43000 0 0 $X=20645 $Y=42885
X14461 271 502 478 653 456 1030 1034 ICV_58 $T=37100 51400 1 0 $X=36985 $Y=49885
X14462 271 502 364 680 365 677 663 ICV_58 $T=39760 45800 1 0 $X=39645 $Y=44285
X14463 271 502 478 888 718 1053 1047 ICV_58 $T=41660 51400 1 0 $X=41545 $Y=49885
X14464 271 502 478 670 456 707 714 ICV_58 $T=43940 48600 0 0 $X=43825 $Y=48485
X14465 271 502 434 456 697 912 479 ICV_58 $T=45650 45800 1 0 $X=45535 $Y=44285
X14466 271 502 479 326 393 467 478 ICV_58 $T=48690 48600 1 0 $X=48575 $Y=47085
X14467 271 502 736 1067 915 923 739 ICV_58 $T=49260 29000 0 0 $X=49145 $Y=28885
X14554 963 49 767 502 964 46 271 OAI211_X1 $T=7650 48600 1 0 $X=7535 $Y=47085
X14555 289 263 844 502 259 264 271 OAI211_X1 $T=29880 51400 0 180 $X=28815 $Y=49885
X14556 647 305 637 502 302 858 271 OAI211_X1 $T=33870 43000 0 180 $X=32805 $Y=41485
X14557 342 291 1030 502 354 360 271 OAI211_X1 $T=36150 51400 0 0 $X=36035 $Y=51285
X14558 1041 291 887 502 1136 399 271 OAI211_X1 $T=39760 51400 1 0 $X=39645 $Y=49885
X14559 451 454 1147 502 457 443 271 OAI211_X1 $T=47930 17800 1 0 $X=47815 $Y=16285
X14560 970 83 502 53 91 271 57 520 AOI221_X1 $T=9550 48600 0 0 $X=9435 $Y=48485
X14561 118 74 502 534 97 271 204 556 AOI221_X1 $T=14300 9400 1 0 $X=14185 $Y=7885
X14562 97 224 502 100 104 271 76 1108 AOI221_X1 $T=14680 9400 0 0 $X=14565 $Y=9285
X14563 97 106 502 105 109 271 205 549 AOI221_X1 $T=15250 15000 1 0 $X=15135 $Y=13485
X14564 97 112 502 107 109 271 589 140 AOI221_X1 $T=15440 9400 1 0 $X=15325 $Y=7885
X14565 109 207 502 978 75 271 202 809 AOI221_X1 $T=15630 15000 0 0 $X=15515 $Y=14885
X14566 544 117 502 113 115 271 121 214 AOI221_X1 $T=15820 23400 1 0 $X=15705 $Y=21885
X14567 142 119 502 985 109 271 81 561 AOI221_X1 $T=16770 15000 0 0 $X=16655 $Y=14885
X14568 556 117 502 137 140 271 121 165 AOI221_X1 $T=18100 9400 0 0 $X=17985 $Y=9285
X14569 118 204 502 129 142 271 225 158 AOI221_X1 $T=18290 15000 1 0 $X=18175 $Y=13485
X14570 151 764 502 165 168 271 164 414 AOI221_X1 $T=20570 12200 1 0 $X=20455 $Y=10685
X14571 180 191 502 173 151 271 106 265 AOI221_X1 $T=22470 26200 0 180 $X=21215 $Y=24685
X14572 138 303 502 181 187 271 368 822 AOI221_X1 $T=22470 26200 1 0 $X=22355 $Y=24685
X14573 106 1008 502 222 225 271 227 181 AOI221_X1 $T=25320 20600 0 0 $X=25205 $Y=20485
X14574 587 377 502 231 233 271 308 222 AOI221_X1 $T=26460 20600 0 0 $X=26345 $Y=20485
X14575 143 366 502 232 237 271 620 246 AOI221_X1 $T=26650 15000 0 0 $X=26535 $Y=14885
X14576 132 243 502 239 235 271 679 241 AOI221_X1 $T=27980 9400 0 180 $X=26725 $Y=7885
X14577 207 837 502 241 81 271 602 240 AOI221_X1 $T=27030 12200 1 0 $X=26915 $Y=10685
X14578 224 1125 502 1216 112 271 267 231 AOI221_X1 $T=27030 20600 1 0 $X=26915 $Y=19085
X14579 221 852 502 260 269 271 267 611 AOI221_X1 $T=29690 20600 1 0 $X=29575 $Y=19085
X14580 617 315 502 291 296 271 292 1021 AOI221_X1 $T=31400 45800 0 0 $X=31285 $Y=45685
X14581 1163 357 502 307 146 271 377 623 AOI221_X1 $T=33110 20600 0 0 $X=32995 $Y=20485
X14582 287 627 502 310 309 271 654 1033 AOI221_X1 $T=33300 26200 0 0 $X=33185 $Y=26085
X14583 1240 221 502 319 325 271 269 333 AOI221_X1 $T=33870 20600 1 0 $X=33755 $Y=19085
X14584 658 336 502 604 332 271 650 384 AOI221_X1 $T=35960 12200 1 180 $X=34705 $Y=12085
X14585 341 247 502 340 328 271 832 656 AOI221_X1 $T=36530 6600 1 180 $X=35275 $Y=6485
X14586 334 69 502 337 341 271 377 891 AOI221_X1 $T=35390 9400 1 0 $X=35275 $Y=7885
X14587 330 335 502 338 341 271 308 332 AOI221_X1 $T=35390 12200 1 0 $X=35275 $Y=10685
X14588 330 344 502 351 355 271 368 666 AOI221_X1 $T=36530 9400 1 0 $X=36415 $Y=7885
X14589 361 377 502 330 328 271 356 352 AOI221_X1 $T=37100 15000 0 0 $X=36985 $Y=14885
X14590 146 683 502 384 388 271 304 418 AOI221_X1 $T=39760 12200 0 0 $X=39645 $Y=12085
X14591 386 682 502 394 396 271 692 1137 AOI221_X1 $T=40710 20600 1 0 $X=40595 $Y=19085
X14592 493 720 502 440 450 271 421 715 AOI221_X1 $T=46980 17800 0 180 $X=45725 $Y=16285
X14593 461 730 502 443 442 271 439 415 AOI221_X1 $T=47550 15000 1 180 $X=46295 $Y=14885
X14594 583 915 502 449 451 271 454 457 AOI221_X1 $T=47550 20600 1 0 $X=47435 $Y=19085
X14595 972 70 1102 973 271 502 972 70 973 ICV_64 $T=12020 45800 1 0 $X=11905 $Y=44285
X14596 85 90 791 793 271 502 85 90 793 ICV_64 $T=13920 45800 1 0 $X=13805 $Y=44285
X14597 211 226 829 834 271 502 211 226 834 ICV_64 $T=25700 51400 1 0 $X=25585 $Y=49885
X14598 218 228 1120 833 271 502 218 228 833 ICV_64 $T=25890 48600 0 0 $X=25775 $Y=48485
X14599 296 292 843 297 271 502 635 292 297 ICV_64 $T=31400 48600 1 0 $X=31285 $Y=47085
X14600 260 200 337 861 271 502 330 274 861 ICV_64 $T=33110 9400 1 0 $X=32995 $Y=7885
X14601 1026 349 870 875 271 502 1026 349 875 ICV_64 $T=36340 31800 1 0 $X=36225 $Y=30285
X14602 722 292 916 921 271 502 732 326 1062 ICV_64 $T=47360 40200 0 0 $X=47245 $Y=40085
X14689 548 271 517 525 161 120 502 NAND4_X1 $T=15630 43000 1 180 $X=14565 $Y=42885
X14690 873 271 1033 1029 1020 672 502 NAND4_X1 $T=37290 26200 1 0 $X=37175 $Y=24685
X14691 711 271 1137 715 925 704 502 NAND4_X1 $T=45650 17800 1 180 $X=44585 $Y=17685
X14714 76 502 55 67 271 97 NOR3_X1 $T=12780 17800 0 180 $X=11905 $Y=16285
X14715 1232 502 517 525 271 546 NOR3_X1 $T=14870 48600 0 0 $X=14755 $Y=48485
X14716 542 502 794 980 271 1107 NOR3_X1 $T=16010 34600 0 180 $X=15135 $Y=33085
X14717 117 502 544 113 271 797 NOR3_X1 $T=15630 20600 0 0 $X=15515 $Y=20485
X14718 796 502 541 111 271 554 NOR3_X1 $T=16390 34600 0 0 $X=16275 $Y=34485
X14719 601 502 250 283 271 218 NOR3_X1 $T=28930 45800 0 180 $X=28055 $Y=44285
X14720 339 502 273 798 271 629 NOR3_X1 $T=29690 40200 1 180 $X=28815 $Y=40085
X14721 124 502 269 303 271 849 NOR3_X1 $T=29500 26200 1 0 $X=29385 $Y=24685
X14722 1019 502 295 603 271 601 NOR3_X1 $T=30830 45800 0 180 $X=29955 $Y=44285
X14723 260 502 221 852 271 615 NOR3_X1 $T=30260 17800 0 0 $X=30145 $Y=17685
X14724 305 502 575 288 271 663 NOR3_X1 $T=32160 43000 1 0 $X=32045 $Y=41485
X14725 640 502 653 639 271 1019 NOR3_X1 $T=33300 37400 1 180 $X=32425 $Y=37285
X14726 69 502 638 607 271 341 NOR3_X1 $T=33110 12200 0 0 $X=32995 $Y=12085
X14727 868 502 347 665 271 640 NOR3_X1 $T=36910 37400 1 180 $X=36035 $Y=37285
X14728 1166 502 670 888 271 868 NOR3_X1 $T=37670 37400 1 180 $X=36795 $Y=37285
X14729 314 502 397 393 271 363 NOR3_X1 $T=39570 37400 0 180 $X=38695 $Y=35885
X14730 676 502 386 681 271 353 NOR3_X1 $T=39190 26200 1 0 $X=39075 $Y=24685
X14731 1049 502 393 314 271 900 NOR3_X1 $T=42990 37400 1 0 $X=42875 $Y=35885
X14741 763 24 271 502 1230 1101 24 1174 ICV_72 $T=1000 54200 0 0 $X=885 $Y=54085
X14742 949 15 271 502 128 1097 15 202 ICV_72 $T=1760 9400 1 0 $X=1645 $Y=7885
X14743 503 15 271 502 762 1090 15 179 ICV_72 $T=2330 20600 0 0 $X=2215 $Y=20485
X14744 1086 15 271 502 960 758 15 94 ICV_72 $T=2330 40200 1 0 $X=2215 $Y=38685
X14745 955 15 271 502 794 48 15 101 ICV_72 $T=3850 34600 1 0 $X=3735 $Y=33085
X14746 518 24 271 502 530 786 24 547 ICV_72 $T=8980 57000 1 0 $X=8865 $Y=55485
X14747 521 15 271 502 157 785 15 589 ICV_72 $T=10310 6600 0 0 $X=10195 $Y=6485
X14748 1114 15 271 502 166 810 38 303 ICV_72 $T=15440 3800 0 0 $X=15325 $Y=3685
X14749 997 38 271 502 840 1187 38 832 ICV_72 $T=22280 3800 1 0 $X=22165 $Y=2285
X14750 835 24 271 502 584 1192 24 1190 ICV_72 $T=22280 57000 1 0 $X=22165 $Y=55485
X14751 1201 24 271 502 1142 1223 24 1064 ICV_72 $T=42230 54200 1 0 $X=42115 $Y=52685
X14752 976 502 70 979 108 548 271 NOR4_X1 $T=14680 43000 1 0 $X=14565 $Y=41485
X14753 295 502 603 250 283 842 271 NOR4_X1 $T=29310 37400 0 0 $X=29195 $Y=37285
X14754 347 502 665 653 639 280 271 NOR4_X1 $T=36150 37400 1 180 $X=35085 $Y=37285
X14755 359 502 317 670 888 674 271 NOR4_X1 $T=39190 40200 0 180 $X=38125 $Y=38685
X14756 672 502 904 688 1044 711 271 NOR4_X1 $T=43180 23400 1 180 $X=42115 $Y=23285
X14757 507 29 759 271 22 1227 502 AOI211_X1 $T=2330 48600 0 0 $X=2215 $Y=48485
X14758 507 40 961 271 22 1172 502 AOI211_X1 $T=4800 45800 1 0 $X=4685 $Y=44285
X14759 541 111 783 271 550 802 502 AOI211_X1 $T=15630 37400 1 0 $X=15515 $Y=35885
X14760 154 171 169 271 553 570 502 AOI211_X1 $T=21900 31800 0 180 $X=20835 $Y=30285
X14761 208 234 260 271 117 1121 502 AOI211_X1 $T=27600 26200 1 180 $X=26535 $Y=26085
X14762 600 124 260 271 849 1188 502 AOI211_X1 $T=28550 26200 1 0 $X=28435 $Y=24685
X14763 325 221 319 271 631 1163 502 AOI211_X1 $T=33870 17800 1 180 $X=32805 $Y=17685
X14764 373 398 359 271 317 1166 502 AOI211_X1 $T=40900 37400 0 0 $X=40785 $Y=37285
X14778 802 271 160 562 502 169 NAND3_X1 $T=17910 31800 0 0 $X=17795 $Y=31685
X14779 141 271 144 116 502 979 NAND3_X1 $T=19430 43000 1 180 $X=18555 $Y=42885
X14780 156 271 210 194 502 539 NAND3_X1 $T=21900 40200 1 180 $X=21025 $Y=40085
X14781 826 271 570 1003 502 310 NAND3_X1 $T=24180 29000 1 180 $X=23305 $Y=28885
X14782 328 271 221 223 502 586 NAND3_X1 $T=25320 29000 1 0 $X=25205 $Y=27485
X14783 884 271 373 674 502 1015 NAND3_X1 $T=39190 37400 1 180 $X=38315 $Y=37285
X14784 78 271 502 537 ICV_73 $T=12780 15000 1 0 $X=12665 $Y=13485
X14785 541 271 502 542 ICV_73 $T=13540 34600 0 0 $X=13425 $Y=34485
X14786 539 271 502 53 ICV_73 $T=13540 45800 0 0 $X=13425 $Y=45685
X14787 977 271 502 545 ICV_73 $T=14300 17800 1 0 $X=14185 $Y=16285
X14788 762 271 502 138 ICV_73 $T=18290 26200 1 0 $X=18175 $Y=24685
X14789 106 271 502 587 ICV_73 $T=25320 20600 1 0 $X=25205 $Y=19085
X14790 246 271 502 248 ICV_73 $T=27980 15000 1 0 $X=27865 $Y=13485
X14791 368 271 502 227 ICV_73 $T=27980 20600 0 0 $X=27865 $Y=20485
X14792 190 271 502 276 ICV_73 $T=28930 6600 0 0 $X=28815 $Y=6485
X14793 600 271 502 605 ICV_73 $T=29500 23400 1 0 $X=29385 $Y=21885
X14794 859 271 502 296 ICV_73 $T=31590 45800 1 0 $X=31475 $Y=44285
X14795 286 271 502 350 ICV_73 $T=34630 20600 0 0 $X=34515 $Y=20485
X14796 1164 271 502 340 ICV_73 $T=35770 6600 1 0 $X=35655 $Y=5085
X14797 662 271 502 362 ICV_73 $T=36530 12200 1 0 $X=36415 $Y=10685
X14816 161 91 120 271 502 478 AND3_X1 $T=17530 40200 0 180 $X=16465 $Y=38685
X14817 109 815 164 271 502 173 AND3_X1 $T=20380 26200 1 0 $X=20265 $Y=24685
X14818 1015 280 842 271 502 210 AND3_X1 $T=28360 40200 1 0 $X=28245 $Y=38685
X14819 328 605 304 271 502 307 AND3_X1 $T=32160 20600 0 0 $X=32045 $Y=20485
X14820 76 109 113 271 502 NOR2_X2 $T=14300 23400 0 180 $X=13235 $Y=21885
X14821 124 164 801 271 502 NOR2_X2 $T=18290 26200 0 180 $X=17225 $Y=24685
X14822 208 191 801 271 502 NOR2_X2 $T=17530 26200 0 0 $X=17415 $Y=26085
X14823 90 718 1158 271 502 NOR2_X2 $T=23420 48600 0 180 $X=22355 $Y=47085
X14824 290 361 319 271 502 NOR2_X2 $T=31400 17800 1 0 $X=31285 $Y=16285
X14825 288 364 273 305 271 502 NOR3_X2 $T=31020 40200 1 180 $X=29575 $Y=40085
X14826 288 322 575 339 271 502 NOR3_X2 $T=32350 40200 1 180 $X=30905 $Y=40085
X14829 504 271 502 51 CLKBUF_X1 $T=8600 48600 0 0 $X=8485 $Y=48485
X14830 1156 271 502 117 CLKBUF_X1 $T=14490 29000 1 0 $X=14375 $Y=27485
X14831 1160 271 502 339 CLKBUF_X1 $T=23610 45800 0 180 $X=22925 $Y=44285
X14832 591 271 502 288 CLKBUF_X1 $T=26270 40200 1 0 $X=26155 $Y=38685
X14833 592 271 502 292 CLKBUF_X1 $T=27220 45800 1 0 $X=27105 $Y=44285
X14834 539 271 161 479 693 502 OAI21_X2 $T=21140 40200 1 180 $X=19695 $Y=40085
X14835 827 271 124 269 121 502 OAI21_X2 $T=24750 26200 1 0 $X=24635 $Y=24685
X14836 766 519 517 271 502 63 HA_X1 $T=7840 51400 0 0 $X=7725 $Y=51285
X14837 781 776 58 271 502 519 HA_X1 $T=11640 51400 1 180 $X=9625 $Y=51285
X14838 540 1177 86 271 502 776 HA_X1 $T=14110 51400 1 0 $X=13995 $Y=49885
X14839 1111 819 116 271 502 1177 HA_X1 $T=16390 51400 1 0 $X=16275 $Y=49885
X14840 552 108 161 271 502 807 HA_X1 $T=16770 45800 0 0 $X=16655 $Y=45685
X14841 563 807 141 271 502 996 HA_X1 $T=19620 48600 1 0 $X=19505 $Y=47085
X14842 814 996 144 271 502 819 HA_X1 $T=20000 48600 0 0 $X=19885 $Y=48485
X14843 273 1006 210 271 502 581 HA_X1 $T=23610 43000 1 0 $X=23495 $Y=41485
X14844 1160 1241 211 271 502 1006 HA_X1 $T=25700 43000 1 180 $X=23685 $Y=42885
X14845 1243 1120 1183 271 502 184 HA_X1 $T=25700 48600 0 180 $X=23685 $Y=47085
X14846 591 581 194 271 502 1244 HA_X1 $T=26270 40200 0 180 $X=24255 $Y=38685
X14847 592 1005 218 271 502 1241 HA_X1 $T=26270 45800 0 180 $X=24255 $Y=44285
X14848 191 502 168 157 151 164 582 407 271 AOI222_X2 $T=23610 9400 0 0 $X=23495 $Y=9285
X14849 164 502 136 589 151 191 582 216 271 AOI222_X2 $T=26650 12200 0 180 $X=23875 $Y=10685
X14850 191 502 136 205 151 164 579 450 271 AOI222_X2 $T=23990 15000 1 0 $X=23875 $Y=13485
X14851 1232 114 804 58 502 271 FA_X1 $T=15630 54200 1 0 $X=15515 $Y=52685
X14852 114 147 808 1001 502 271 FA_X1 $T=18860 51400 0 0 $X=18745 $Y=51285
X14853 147 172 1002 834 502 271 FA_X1 $T=21140 54200 1 0 $X=21025 $Y=52685
X14854 172 184 829 833 502 271 FA_X1 $T=22280 51400 0 0 $X=22165 $Y=51285
X14855 796 542 794 271 111 541 1157 133 502 OAI33_X1 $T=16010 34600 1 0 $X=15895 $Y=33085
X14856 121 115 113 271 117 560 138 180 502 OAI33_X1 $T=17530 23400 0 0 $X=17415 $Y=23285
X14857 271 30 23 502 271 15 271 CLKGATETST_X1 $T=2900 37400 1 0 $X=2785 $Y=35885
X14858 271 47 51 502 271 24 271 CLKGATETST_X1 $T=7080 51400 1 0 $X=6965 $Y=49885
.ENDS
***************************************
