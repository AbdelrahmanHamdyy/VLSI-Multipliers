/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Jan  4 01:36:47 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3422931764 */

/* blackbox module unsigned_seq_multiplier_bbox */

module fp_mul(clk, rst, a_s, b_s, c_out, overflow);
   input clk;
   input rst;
   input [31:0]a_s;
   input [31:0]b_s;
   output [31:0]c_out;
   output overflow;

   wire [25:0]res_mant;
   wire mul_start;
   wire n_0_1;
   wire b;
   wire a;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire [4:0]counter;
   wire n_0_50;
   wire n_0_0;
   wire n_0_0_18;
   wire n_0_0_2;
   wire n_0_0_19;
   wire n_0_0_3;
   wire n_0_0_20;
   wire n_0_0_4;
   wire n_0_0_21;
   wire n_0_0_5;
   wire n_0_0_22;
   wire n_0_0_6;
   wire n_0_0_23;
   wire n_0_0_7;
   wire n_0_0_24;
   wire n_0_0_8;
   wire n_0_0_25;
   wire n_0_0_0;
   wire n_0_0_26;
   wire n_0_0_1;
   wire n_0_0_27;
   wire n_0_0_9;
   wire n_0_0_28;
   wire n_0_0_10;
   wire n_0_0_29;
   wire n_0_0_11;
   wire n_0_0_30;
   wire n_0_0_12;
   wire n_0_0_31;
   wire n_0_0_13;
   wire n_0_0_32;
   wire n_0_0_14;
   wire n_0_0_33;
   wire n_0_0_15;
   wire n_0_18;
   wire n_0_0_34;
   wire n_0_19;
   wire n_0_0_35;
   wire n_0_20;
   wire n_0_0_36;
   wire n_0_21;
   wire n_0_0_37;
   wire n_0_22;
   wire n_0_0_38;
   wire n_0_23;
   wire n_0_0_39;
   wire n_0_24;
   wire n_0_0_40;
   wire n_0_25;
   wire n_0_0_41;
   wire n_0_26;
   wire n_0_0_42;
   wire n_0_27;
   wire n_0_0_43;
   wire n_0_28;
   wire n_0_0_44;
   wire n_0_29;
   wire n_0_0_45;
   wire n_0_30;
   wire n_0_0_46;
   wire n_0_31;
   wire n_0_0_47;
   wire n_0_32;
   wire n_0_0_48;
   wire n_0_33;
   wire n_0_0_49;
   wire n_0_34;
   wire n_0_0_50;
   wire n_0_35;
   wire n_0_0_51;
   wire n_0_36;
   wire n_0_0_52;
   wire n_0_37;
   wire n_0_0_53;
   wire n_0_38;
   wire n_0_0_54;
   wire n_0_39;
   wire n_0_0_55;
   wire n_0_40;
   wire n_0_0_56;
   wire n_0_41;
   wire n_0_42;
   wire n_0_0_57;
   wire n_0_43;
   wire n_0_0_58;
   wire n_0_44;
   wire n_0_0_59;
   wire n_0_45;
   wire n_0_0_60;
   wire n_0_46;
   wire n_0_0_61;
   wire n_0_47;
   wire n_0_0_62;
   wire n_0_48;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_49;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_0_76;
   wire n_0_58;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_16;
   wire n_0_0_81;
   wire n_0_59;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire start;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_57;
   wire n_0_0_17;

   unsigned_seq_multiplier_bbox unsigned_seq_multiplier_dut (.start_s(mul_start), 
      .clk(clk), .rst(rst), .a({1'b1, n_23, n_24, n_25, n_26, n_27, n_28, n_29, 
      n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, 
      n_42, n_43, n_44, n_45}), .b({1'b1, n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, 
      n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, 
      n_21, n_22}), .c({res_mant[25], res_mant[24], res_mant[23], res_mant[22], 
      res_mant[21], res_mant[20], res_mant[19], res_mant[18], res_mant[17], 
      res_mant[16], res_mant[15], res_mant[14], res_mant[13], res_mant[12], 
      res_mant[11], res_mant[10], res_mant[9], res_mant[8], res_mant[7], 
      res_mant[6], res_mant[5], res_mant[4], res_mant[3], res_mant[2], 
      res_mant[1], res_mant[0], uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, 
      uc_19, uc_20, uc_21}));
   DFF_X1 overflow_reg (.D(n_0_58), .CK(n_0_50), .Q(overflow), .QN());
   DFF_X1 \c_out_reg[31]  (.D(n_0_49), .CK(n_0_50), .Q(c_out[31]), .QN());
   DFF_X1 \c_out_reg[30]  (.D(n_0_48), .CK(n_0_50), .Q(c_out[30]), .QN());
   DFF_X1 \c_out_reg[29]  (.D(n_0_47), .CK(n_0_50), .Q(c_out[29]), .QN());
   DFF_X1 \c_out_reg[28]  (.D(n_0_46), .CK(n_0_50), .Q(c_out[28]), .QN());
   DFF_X1 \c_out_reg[27]  (.D(n_0_45), .CK(n_0_50), .Q(c_out[27]), .QN());
   DFF_X1 \c_out_reg[26]  (.D(n_0_44), .CK(n_0_50), .Q(c_out[26]), .QN());
   DFF_X1 \c_out_reg[25]  (.D(n_0_43), .CK(n_0_50), .Q(c_out[25]), .QN());
   DFF_X1 \c_out_reg[24]  (.D(n_0_42), .CK(n_0_50), .Q(c_out[24]), .QN());
   DFF_X1 \c_out_reg[23]  (.D(n_0_41), .CK(n_0_50), .Q(c_out[23]), .QN());
   DFF_X1 \c_out_reg[22]  (.D(n_0_40), .CK(n_0_50), .Q(c_out[22]), .QN());
   DFF_X1 \c_out_reg[21]  (.D(n_0_39), .CK(n_0_50), .Q(c_out[21]), .QN());
   DFF_X1 \c_out_reg[20]  (.D(n_0_38), .CK(n_0_50), .Q(c_out[20]), .QN());
   DFF_X1 \c_out_reg[19]  (.D(n_0_37), .CK(n_0_50), .Q(c_out[19]), .QN());
   DFF_X1 \c_out_reg[18]  (.D(n_0_36), .CK(n_0_50), .Q(c_out[18]), .QN());
   DFF_X1 \c_out_reg[17]  (.D(n_0_35), .CK(n_0_50), .Q(c_out[17]), .QN());
   DFF_X1 \c_out_reg[16]  (.D(n_0_34), .CK(n_0_50), .Q(c_out[16]), .QN());
   DFF_X1 \c_out_reg[15]  (.D(n_0_33), .CK(n_0_50), .Q(c_out[15]), .QN());
   DFF_X1 \c_out_reg[14]  (.D(n_0_32), .CK(n_0_50), .Q(c_out[14]), .QN());
   DFF_X1 \c_out_reg[13]  (.D(n_0_31), .CK(n_0_50), .Q(c_out[13]), .QN());
   DFF_X1 \c_out_reg[12]  (.D(n_0_30), .CK(n_0_50), .Q(c_out[12]), .QN());
   DFF_X1 \c_out_reg[11]  (.D(n_0_29), .CK(n_0_50), .Q(c_out[11]), .QN());
   DFF_X1 \c_out_reg[10]  (.D(n_0_28), .CK(n_0_50), .Q(c_out[10]), .QN());
   DFF_X1 \c_out_reg[9]  (.D(n_0_27), .CK(n_0_50), .Q(c_out[9]), .QN());
   DFF_X1 \c_out_reg[8]  (.D(n_0_26), .CK(n_0_50), .Q(c_out[8]), .QN());
   DFF_X1 \c_out_reg[7]  (.D(n_0_25), .CK(n_0_50), .Q(c_out[7]), .QN());
   DFF_X1 \c_out_reg[6]  (.D(n_0_24), .CK(n_0_50), .Q(c_out[6]), .QN());
   DFF_X1 \c_out_reg[5]  (.D(n_0_23), .CK(n_0_50), .Q(c_out[5]), .QN());
   DFF_X1 \c_out_reg[4]  (.D(n_0_22), .CK(n_0_50), .Q(c_out[4]), .QN());
   DFF_X1 \c_out_reg[3]  (.D(n_0_21), .CK(n_0_50), .Q(c_out[3]), .QN());
   DFF_X1 \c_out_reg[2]  (.D(n_0_20), .CK(n_0_50), .Q(c_out[2]), .QN());
   DFF_X1 \c_out_reg[1]  (.D(n_0_19), .CK(n_0_50), .Q(c_out[1]), .QN());
   DFF_X1 \c_out_reg[0]  (.D(n_0_18), .CK(n_0_50), .Q(c_out[0]), .QN());
   DFF_X1 \b_reg[22]  (.D(b_s[22]), .CK(n_0_0), .Q(n_0), .QN());
   DFF_X1 \b_reg[21]  (.D(b_s[21]), .CK(n_0_0), .Q(n_1), .QN());
   DFF_X1 \b_reg[20]  (.D(b_s[20]), .CK(n_0_0), .Q(n_2), .QN());
   DFF_X1 \b_reg[19]  (.D(b_s[19]), .CK(n_0_0), .Q(n_3), .QN());
   DFF_X1 \b_reg[18]  (.D(b_s[18]), .CK(n_0_0), .Q(n_4), .QN());
   DFF_X1 \b_reg[17]  (.D(b_s[17]), .CK(n_0_0), .Q(n_5), .QN());
   DFF_X1 \b_reg[16]  (.D(b_s[16]), .CK(n_0_0), .Q(n_6), .QN());
   DFF_X1 \b_reg[15]  (.D(b_s[15]), .CK(n_0_0), .Q(n_7), .QN());
   DFF_X1 \b_reg[14]  (.D(b_s[14]), .CK(n_0_0), .Q(n_8), .QN());
   DFF_X1 \b_reg[13]  (.D(b_s[13]), .CK(n_0_0), .Q(n_9), .QN());
   DFF_X1 \b_reg[12]  (.D(b_s[12]), .CK(n_0_0), .Q(n_10), .QN());
   DFF_X1 \b_reg[11]  (.D(b_s[11]), .CK(n_0_0), .Q(n_11), .QN());
   DFF_X1 \b_reg[10]  (.D(b_s[10]), .CK(n_0_0), .Q(n_12), .QN());
   DFF_X1 \b_reg[9]  (.D(b_s[9]), .CK(n_0_0), .Q(n_13), .QN());
   DFF_X1 \b_reg[8]  (.D(b_s[8]), .CK(n_0_0), .Q(n_14), .QN());
   DFF_X1 \b_reg[7]  (.D(b_s[7]), .CK(n_0_0), .Q(n_15), .QN());
   DFF_X1 \b_reg[6]  (.D(b_s[6]), .CK(n_0_0), .Q(n_16), .QN());
   DFF_X1 \b_reg[5]  (.D(b_s[5]), .CK(n_0_0), .Q(n_17), .QN());
   DFF_X1 \b_reg[4]  (.D(b_s[4]), .CK(n_0_0), .Q(n_18), .QN());
   DFF_X1 \b_reg[3]  (.D(b_s[3]), .CK(n_0_0), .Q(n_19), .QN());
   DFF_X1 \b_reg[2]  (.D(b_s[2]), .CK(n_0_0), .Q(n_20), .QN());
   DFF_X1 \b_reg[1]  (.D(b_s[1]), .CK(n_0_0), .Q(n_21), .QN());
   DFF_X1 \b_reg[0]  (.D(b_s[0]), .CK(n_0_0), .Q(n_22), .QN());
   DFF_X1 \a_reg[22]  (.D(a_s[22]), .CK(n_0_0), .Q(n_23), .QN());
   DFF_X1 \a_reg[21]  (.D(a_s[21]), .CK(n_0_0), .Q(n_24), .QN());
   DFF_X1 \a_reg[20]  (.D(a_s[20]), .CK(n_0_0), .Q(n_25), .QN());
   DFF_X1 \a_reg[19]  (.D(a_s[19]), .CK(n_0_0), .Q(n_26), .QN());
   DFF_X1 \a_reg[18]  (.D(a_s[18]), .CK(n_0_0), .Q(n_27), .QN());
   DFF_X1 \a_reg[17]  (.D(a_s[17]), .CK(n_0_0), .Q(n_28), .QN());
   DFF_X1 \a_reg[16]  (.D(a_s[16]), .CK(n_0_0), .Q(n_29), .QN());
   DFF_X1 \a_reg[15]  (.D(a_s[15]), .CK(n_0_0), .Q(n_30), .QN());
   DFF_X1 \a_reg[14]  (.D(a_s[14]), .CK(n_0_0), .Q(n_31), .QN());
   DFF_X1 \a_reg[13]  (.D(a_s[13]), .CK(n_0_0), .Q(n_32), .QN());
   DFF_X1 \a_reg[12]  (.D(a_s[12]), .CK(n_0_0), .Q(n_33), .QN());
   DFF_X1 \a_reg[11]  (.D(a_s[11]), .CK(n_0_0), .Q(n_34), .QN());
   DFF_X1 \a_reg[10]  (.D(a_s[10]), .CK(n_0_0), .Q(n_35), .QN());
   DFF_X1 \a_reg[9]  (.D(a_s[9]), .CK(n_0_0), .Q(n_36), .QN());
   DFF_X1 \a_reg[8]  (.D(a_s[8]), .CK(n_0_0), .Q(n_37), .QN());
   DFF_X1 \a_reg[7]  (.D(a_s[7]), .CK(n_0_0), .Q(n_38), .QN());
   DFF_X1 \a_reg[6]  (.D(a_s[6]), .CK(n_0_0), .Q(n_39), .QN());
   DFF_X1 \a_reg[5]  (.D(a_s[5]), .CK(n_0_0), .Q(n_40), .QN());
   DFF_X1 \a_reg[4]  (.D(a_s[4]), .CK(n_0_0), .Q(n_41), .QN());
   DFF_X1 \a_reg[3]  (.D(a_s[3]), .CK(n_0_0), .Q(n_42), .QN());
   DFF_X1 \a_reg[2]  (.D(a_s[2]), .CK(n_0_0), .Q(n_43), .QN());
   DFF_X1 \a_reg[1]  (.D(a_s[1]), .CK(n_0_0), .Q(n_44), .QN());
   DFF_X1 \a_reg[0]  (.D(a_s[0]), .CK(n_0_0), .Q(n_45), .QN());
   DFF_X1 mul_start_reg (.D(n_0_1), .CK(clk), .Q(mul_start), .QN());
   MUX2_X1 mul_start_reg_enable_mux_0 (.A(mul_start), .B(start), .S(n_0_57), 
      .Z(n_0_1));
   DFF_X1 \b_reg[31]  (.D(b_s[31]), .CK(n_0_0), .Q(b), .QN());
   DFF_X1 \a_reg[31]  (.D(a_s[31]), .CK(n_0_0), .Q(a), .QN());
   DFF_X1 \b_reg[30]  (.D(b_s[30]), .CK(n_0_0), .Q(n_0_2), .QN());
   DFF_X1 \b_reg[29]  (.D(b_s[29]), .CK(n_0_0), .Q(n_0_3), .QN());
   DFF_X1 \b_reg[28]  (.D(b_s[28]), .CK(n_0_0), .Q(n_0_4), .QN());
   DFF_X1 \b_reg[27]  (.D(b_s[27]), .CK(n_0_0), .Q(n_0_5), .QN());
   DFF_X1 \b_reg[26]  (.D(b_s[26]), .CK(n_0_0), .Q(n_0_6), .QN());
   DFF_X1 \b_reg[25]  (.D(b_s[25]), .CK(n_0_0), .Q(n_0_7), .QN());
   DFF_X1 \b_reg[24]  (.D(b_s[24]), .CK(n_0_0), .Q(n_0_8), .QN());
   DFF_X1 \b_reg[23]  (.D(b_s[23]), .CK(n_0_0), .Q(n_0_9), .QN());
   DFF_X1 \a_reg[30]  (.D(a_s[30]), .CK(n_0_0), .Q(n_0_10), .QN());
   DFF_X1 \a_reg[29]  (.D(a_s[29]), .CK(n_0_0), .Q(n_0_11), .QN());
   DFF_X1 \a_reg[28]  (.D(a_s[28]), .CK(n_0_0), .Q(n_0_12), .QN());
   DFF_X1 \a_reg[27]  (.D(a_s[27]), .CK(n_0_0), .Q(n_0_13), .QN());
   DFF_X1 \a_reg[26]  (.D(a_s[26]), .CK(n_0_0), .Q(n_0_14), .QN());
   DFF_X1 \a_reg[25]  (.D(a_s[25]), .CK(n_0_0), .Q(n_0_15), .QN());
   DFF_X1 \a_reg[24]  (.D(a_s[24]), .CK(n_0_0), .Q(n_0_16), .QN());
   DFF_X1 \a_reg[23]  (.D(a_s[23]), .CK(n_0_0), .Q(n_0_17), .QN());
   DFF_X1 \counter_reg[4]  (.D(n_0_56), .CK(clk), .Q(counter[4]), .QN());
   DFF_X1 \counter_reg[3]  (.D(n_0_55), .CK(clk), .Q(counter[3]), .QN());
   DFF_X1 \counter_reg[2]  (.D(n_0_54), .CK(clk), .Q(counter[2]), .QN());
   DFF_X1 \counter_reg[1]  (.D(n_0_53), .CK(clk), .Q(counter[1]), .QN());
   DFF_X1 \counter_reg[0]  (.D(n_0_52), .CK(clk), .Q(counter[0]), .QN());
   CLKGATETST_X1 clk_gate_overflow_reg (.CK(clk), .E(n_0_59), .SE(1'b0), 
      .GCK(n_0_50));
   CLKGATETST_X1 clk_gate_b_reg (.CK(clk), .E(n_0_51), .SE(1'b0), .GCK(n_0_0));
   FA_X1 i_0_0_0 (.A(n_0_8), .B(n_0_16), .CI(n_0_0_16), .CO(n_0_0_2), .S(
      n_0_0_18));
   FA_X1 i_0_0_1 (.A(n_0_7), .B(n_0_15), .CI(n_0_0_2), .CO(n_0_0_3), .S(n_0_0_19));
   FA_X1 i_0_0_2 (.A(n_0_6), .B(n_0_14), .CI(n_0_0_3), .CO(n_0_0_4), .S(n_0_0_20));
   FA_X1 i_0_0_3 (.A(n_0_5), .B(n_0_13), .CI(n_0_0_4), .CO(n_0_0_5), .S(n_0_0_21));
   FA_X1 i_0_0_4 (.A(n_0_4), .B(n_0_12), .CI(n_0_0_5), .CO(n_0_0_6), .S(n_0_0_22));
   FA_X1 i_0_0_5 (.A(n_0_3), .B(n_0_11), .CI(n_0_0_6), .CO(n_0_0_7), .S(n_0_0_23));
   FA_X1 i_0_0_6 (.A(n_0_10), .B(n_0_0_17), .CI(n_0_0_7), .CO(n_0_0_8), .S(
      n_0_0_24));
   HA_X1 i_0_0_7 (.A(n_0_0_18), .B(n_0_0_80), .CO(n_0_0_0), .S(n_0_0_25));
   HA_X1 i_0_0_8 (.A(n_0_0_19), .B(n_0_0_0), .CO(n_0_0_1), .S(n_0_0_26));
   HA_X1 i_0_0_9 (.A(n_0_0_20), .B(n_0_0_1), .CO(n_0_0_9), .S(n_0_0_27));
   HA_X1 i_0_0_10 (.A(n_0_0_21), .B(n_0_0_9), .CO(n_0_0_10), .S(n_0_0_28));
   HA_X1 i_0_0_11 (.A(n_0_0_22), .B(n_0_0_10), .CO(n_0_0_11), .S(n_0_0_29));
   HA_X1 i_0_0_12 (.A(n_0_0_23), .B(n_0_0_11), .CO(n_0_0_12), .S(n_0_0_30));
   HA_X1 i_0_0_13 (.A(counter[1]), .B(counter[0]), .CO(n_0_0_13), .S(n_0_0_31));
   HA_X1 i_0_0_14 (.A(counter[2]), .B(n_0_0_13), .CO(n_0_0_14), .S(n_0_0_32));
   HA_X1 i_0_0_15 (.A(counter[3]), .B(n_0_0_14), .CO(n_0_0_15), .S(n_0_0_33));
   INV_X1 i_0_0_16 (.A(n_0_0_34), .ZN(n_0_18));
   AOI22_X1 i_0_0_17 (.A1(res_mant[1]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[2]), .ZN(n_0_0_34));
   INV_X1 i_0_0_18 (.A(n_0_0_35), .ZN(n_0_19));
   AOI22_X1 i_0_0_19 (.A1(res_mant[2]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[3]), .ZN(n_0_0_35));
   INV_X1 i_0_0_20 (.A(n_0_0_36), .ZN(n_0_20));
   AOI22_X1 i_0_0_21 (.A1(res_mant[3]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[4]), .ZN(n_0_0_36));
   INV_X1 i_0_0_22 (.A(n_0_0_37), .ZN(n_0_21));
   AOI22_X1 i_0_0_23 (.A1(res_mant[4]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[5]), .ZN(n_0_0_37));
   INV_X1 i_0_0_24 (.A(n_0_0_38), .ZN(n_0_22));
   AOI22_X1 i_0_0_25 (.A1(res_mant[5]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[6]), .ZN(n_0_0_38));
   INV_X1 i_0_0_26 (.A(n_0_0_39), .ZN(n_0_23));
   AOI22_X1 i_0_0_27 (.A1(res_mant[6]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[7]), .ZN(n_0_0_39));
   INV_X1 i_0_0_28 (.A(n_0_0_40), .ZN(n_0_24));
   AOI22_X1 i_0_0_29 (.A1(res_mant[7]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[8]), .ZN(n_0_0_40));
   INV_X1 i_0_0_30 (.A(n_0_0_41), .ZN(n_0_25));
   AOI22_X1 i_0_0_31 (.A1(res_mant[8]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[9]), .ZN(n_0_0_41));
   INV_X1 i_0_0_32 (.A(n_0_0_42), .ZN(n_0_26));
   AOI22_X1 i_0_0_33 (.A1(res_mant[9]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[10]), .ZN(n_0_0_42));
   INV_X1 i_0_0_34 (.A(n_0_0_43), .ZN(n_0_27));
   AOI22_X1 i_0_0_35 (.A1(res_mant[10]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[11]), .ZN(n_0_0_43));
   INV_X1 i_0_0_36 (.A(n_0_0_44), .ZN(n_0_28));
   AOI22_X1 i_0_0_37 (.A1(res_mant[11]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[12]), .ZN(n_0_0_44));
   INV_X1 i_0_0_38 (.A(n_0_0_45), .ZN(n_0_29));
   AOI22_X1 i_0_0_39 (.A1(res_mant[12]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[13]), .ZN(n_0_0_45));
   INV_X1 i_0_0_40 (.A(n_0_0_46), .ZN(n_0_30));
   AOI22_X1 i_0_0_41 (.A1(res_mant[13]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[14]), .ZN(n_0_0_46));
   INV_X1 i_0_0_42 (.A(n_0_0_47), .ZN(n_0_31));
   AOI22_X1 i_0_0_43 (.A1(res_mant[14]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[15]), .ZN(n_0_0_47));
   INV_X1 i_0_0_44 (.A(n_0_0_48), .ZN(n_0_32));
   AOI22_X1 i_0_0_45 (.A1(res_mant[15]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[16]), .ZN(n_0_0_48));
   INV_X1 i_0_0_46 (.A(n_0_0_49), .ZN(n_0_33));
   AOI22_X1 i_0_0_47 (.A1(res_mant[16]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[17]), .ZN(n_0_0_49));
   INV_X1 i_0_0_48 (.A(n_0_0_50), .ZN(n_0_34));
   AOI22_X1 i_0_0_49 (.A1(res_mant[17]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[18]), .ZN(n_0_0_50));
   INV_X1 i_0_0_50 (.A(n_0_0_51), .ZN(n_0_35));
   AOI22_X1 i_0_0_51 (.A1(res_mant[18]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[19]), .ZN(n_0_0_51));
   INV_X1 i_0_0_52 (.A(n_0_0_52), .ZN(n_0_36));
   AOI22_X1 i_0_0_53 (.A1(res_mant[19]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[20]), .ZN(n_0_0_52));
   INV_X1 i_0_0_54 (.A(n_0_0_53), .ZN(n_0_37));
   AOI22_X1 i_0_0_55 (.A1(res_mant[20]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[21]), .ZN(n_0_0_53));
   INV_X1 i_0_0_56 (.A(n_0_0_54), .ZN(n_0_38));
   AOI22_X1 i_0_0_57 (.A1(res_mant[21]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[22]), .ZN(n_0_0_54));
   INV_X1 i_0_0_58 (.A(n_0_0_55), .ZN(n_0_39));
   AOI22_X1 i_0_0_59 (.A1(res_mant[22]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[23]), .ZN(n_0_0_55));
   INV_X1 i_0_0_60 (.A(n_0_0_56), .ZN(n_0_40));
   AOI22_X1 i_0_0_61 (.A1(res_mant[23]), .A2(n_0_0_64), .B1(n_0_0_63), .B2(
      res_mant[24]), .ZN(n_0_0_56));
   MUX2_X1 i_0_0_62 (.A(n_0_0_63), .B(n_0_0_64), .S(n_0_0_80), .Z(n_0_41));
   INV_X1 i_0_0_63 (.A(n_0_0_57), .ZN(n_0_42));
   AOI22_X1 i_0_0_64 (.A1(n_0_0_18), .A2(n_0_0_64), .B1(n_0_0_63), .B2(n_0_0_25), 
      .ZN(n_0_0_57));
   INV_X1 i_0_0_65 (.A(n_0_0_58), .ZN(n_0_43));
   AOI22_X1 i_0_0_66 (.A1(n_0_0_19), .A2(n_0_0_64), .B1(n_0_0_63), .B2(n_0_0_26), 
      .ZN(n_0_0_58));
   INV_X1 i_0_0_67 (.A(n_0_0_59), .ZN(n_0_44));
   AOI22_X1 i_0_0_68 (.A1(n_0_0_20), .A2(n_0_0_64), .B1(n_0_0_63), .B2(n_0_0_27), 
      .ZN(n_0_0_59));
   INV_X1 i_0_0_69 (.A(n_0_0_60), .ZN(n_0_45));
   AOI22_X1 i_0_0_70 (.A1(n_0_0_21), .A2(n_0_0_64), .B1(n_0_0_63), .B2(n_0_0_28), 
      .ZN(n_0_0_60));
   INV_X1 i_0_0_71 (.A(n_0_0_61), .ZN(n_0_46));
   AOI22_X1 i_0_0_72 (.A1(n_0_0_22), .A2(n_0_0_64), .B1(n_0_0_63), .B2(n_0_0_29), 
      .ZN(n_0_0_61));
   INV_X1 i_0_0_73 (.A(n_0_0_62), .ZN(n_0_47));
   AOI22_X1 i_0_0_74 (.A1(n_0_0_23), .A2(n_0_0_64), .B1(n_0_0_63), .B2(n_0_0_30), 
      .ZN(n_0_0_62));
   NOR2_X1 i_0_0_75 (.A1(n_0_0_67), .A2(n_0_0_65), .ZN(n_0_48));
   NOR2_X1 i_0_0_76 (.A1(n_0_0_86), .A2(n_0_0_67), .ZN(n_0_0_63));
   NOR2_X1 i_0_0_77 (.A1(n_0_0_67), .A2(res_mant[25]), .ZN(n_0_0_64));
   XOR2_X1 i_0_0_78 (.A(n_0_0_24), .B(n_0_0_66), .Z(n_0_0_65));
   NAND2_X1 i_0_0_79 (.A1(res_mant[25]), .A2(n_0_0_12), .ZN(n_0_0_66));
   NAND3_X1 i_0_0_80 (.A1(n_0_57), .A2(n_0_0_73), .A3(n_0_0_70), .ZN(n_0_0_67));
   AND2_X1 i_0_0_81 (.A1(n_0_0_68), .A2(n_0_57), .ZN(n_0_49));
   XNOR2_X1 i_0_0_82 (.A(a), .B(n_0_0_69), .ZN(n_0_0_68));
   NAND3_X1 i_0_0_83 (.A1(n_0_0_73), .A2(n_0_0_70), .A3(b), .ZN(n_0_0_69));
   NAND2_X1 i_0_0_84 (.A1(n_0_0_72), .A2(n_0_0_71), .ZN(n_0_0_70));
   NOR4_X1 i_0_0_85 (.A1(n_0_10), .A2(n_0_11), .A3(n_0_12), .A4(n_0_13), 
      .ZN(n_0_0_71));
   NOR4_X1 i_0_0_86 (.A1(n_0_14), .A2(n_0_15), .A3(n_0_16), .A4(n_0_17), 
      .ZN(n_0_0_72));
   NAND2_X1 i_0_0_87 (.A1(n_0_0_75), .A2(n_0_0_74), .ZN(n_0_0_73));
   NOR4_X1 i_0_0_88 (.A1(n_0_2), .A2(n_0_3), .A3(n_0_4), .A4(n_0_5), .ZN(
      n_0_0_74));
   NOR4_X1 i_0_0_89 (.A1(n_0_6), .A2(n_0_7), .A3(n_0_8), .A4(n_0_9), .ZN(
      n_0_0_75));
   AND2_X1 i_0_0_90 (.A1(start), .A2(n_0_57), .ZN(n_0_51));
   NOR2_X1 i_0_0_91 (.A1(rst), .A2(counter[0]), .ZN(n_0_52));
   AND2_X1 i_0_0_92 (.A1(n_0_0_31), .A2(n_0_0_82), .ZN(n_0_53));
   AND2_X1 i_0_0_93 (.A1(n_0_0_32), .A2(n_0_0_82), .ZN(n_0_54));
   AND2_X1 i_0_0_94 (.A1(n_0_0_33), .A2(n_0_0_82), .ZN(n_0_55));
   NOR2_X1 i_0_0_95 (.A1(n_0_59), .A2(n_0_0_76), .ZN(n_0_56));
   XNOR2_X1 i_0_0_96 (.A(counter[4]), .B(n_0_0_15), .ZN(n_0_0_76));
   AOI21_X1 i_0_0_97 (.A(rst), .B1(n_0_0_81), .B2(n_0_0_77), .ZN(n_0_58));
   NAND3_X1 i_0_0_98 (.A1(n_0_0_80), .A2(n_0_0_79), .A3(n_0_0_78), .ZN(n_0_0_77));
   AND4_X1 i_0_0_99 (.A1(res_mant[25]), .A2(n_0_0_18), .A3(n_0_0_19), .A4(
      n_0_0_20), .ZN(n_0_0_78));
   AND4_X1 i_0_0_100 (.A1(n_0_0_21), .A2(n_0_0_22), .A3(n_0_0_23), .A4(n_0_0_24), 
      .ZN(n_0_0_79));
   XNOR2_X1 i_0_0_101 (.A(n_0_9), .B(n_0_17), .ZN(n_0_0_80));
   OR2_X1 i_0_0_102 (.A1(n_0_9), .A2(n_0_17), .ZN(n_0_0_16));
   XNOR2_X1 i_0_0_103 (.A(n_0_0_17), .B(n_0_0_8), .ZN(n_0_0_81));
   INV_X1 i_0_0_104 (.A(n_0_0_82), .ZN(n_0_59));
   AOI21_X1 i_0_0_105 (.A(rst), .B1(counter[3]), .B2(n_0_0_83), .ZN(n_0_0_82));
   NOR2_X1 i_0_0_106 (.A1(n_0_0_85), .A2(n_0_0_84), .ZN(n_0_0_83));
   NAND2_X1 i_0_0_107 (.A1(counter[4]), .A2(counter[0]), .ZN(n_0_0_84));
   NOR4_X1 i_0_0_108 (.A1(n_0_0_85), .A2(counter[0]), .A3(counter[3]), .A4(
      counter[4]), .ZN(start));
   OR2_X1 i_0_0_109 (.A1(counter[2]), .A2(counter[1]), .ZN(n_0_0_85));
   INV_X1 i_0_0_110 (.A(res_mant[25]), .ZN(n_0_0_86));
   INV_X1 i_0_0_111 (.A(rst), .ZN(n_0_57));
   INV_X1 i_0_0_112 (.A(n_0_2), .ZN(n_0_0_17));
endmodule
