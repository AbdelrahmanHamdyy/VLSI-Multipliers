* SPICE NETLIST
***************************************

.SUBCKT MGC_via2_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X2
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_2
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X4
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_5
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MUX2_X1 A S B VSS VDD Z 7 8
** N=14 EP=8 IP=0 FDC=12
M0 VSS S 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 13 A VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 10 9 13 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 14 S 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=715 $Y=90 $D=1
M4 VSS B 14 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=905 $Y=90 $D=1
M5 Z 10 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1095 $Y=90 $D=1
M6 VDD S 9 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M7 11 A VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M8 10 S 11 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M9 12 9 10 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=715 $Y=995 $D=0
M10 VDD B 12 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=905 $Y=995 $D=0
M11 Z 10 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1095 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X8
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT DFF_X1 D CK VSS VDD Q 6 7
** N=22 EP=7 IP=0 FDC=28
M0 VSS 11 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=160 $Y=180 $D=1
M1 19 10 VSS 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=350 $Y=300 $D=1
M2 9 8 19 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.6e-14 AS=1.26e-14 PD=8.4e-07 PS=4.6e-07 $X=540 $Y=300 $D=1
M3 20 11 9 6 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=2.6e-14 PD=8.3e-07 PS=8.4e-07 $X=735 $Y=180 $D=1
M4 VSS D 20 6 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.395e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=925 $Y=180 $D=1
M5 10 9 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=3.395e-14 PD=6.3e-07 PS=8.3e-07 $X=1115 $Y=180 $D=1
M6 VSS CK 11 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1530 $Y=255 $D=1
M7 21 9 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1720 $Y=255 $D=1
M8 12 8 21 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1910 $Y=255 $D=1
M9 22 11 12 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.1e-14 PD=4.7e-07 PS=7e-07 $X=2100 $Y=300 $D=1
M10 VSS 14 22 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.305e-14 PD=7e-07 PS=4.7e-07 $X=2295 $Y=300 $D=1
M11 14 12 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.1e-14 PD=6.3e-07 PS=7e-07 $X=2485 $Y=255 $D=1
M12 VSS 12 QN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=2825 $Y=90 $D=1
M13 Q 14 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=3015 $Y=90 $D=1
M14 VDD 11 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=160 $Y=785 $D=0
M15 15 10 VDD 7 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=350 $Y=1010 $D=0
M16 9 11 15 7 PMOS_VTL L=5e-08 W=9e-08 AD=3.615e-14 AS=1.26e-14 PD=1.13e-06 PS=4.6e-07 $X=540 $Y=1010 $D=0
M17 16 8 9 7 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=3.615e-14 PD=1.12e-06 PS=1.13e-06 $X=735 $Y=765 $D=0
M18 VDD D 16 7 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.145e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=925 $Y=765 $D=0
M19 10 9 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=5.145e-14 PD=9.9e-07 PS=1.12e-06 $X=1115 $Y=870 $D=0
M20 VDD CK 11 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1530 $Y=870 $D=0
M21 17 9 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1720 $Y=870 $D=0
M22 12 11 17 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1910 $Y=870 $D=0
M23 18 8 12 7 PMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.835e-14 PD=4.7e-07 PS=9.1e-07 $X=2100 $Y=1095 $D=0
M24 VDD 14 18 7 PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.305e-14 PD=9.1e-07 PS=4.7e-07 $X=2295 $Y=1095 $D=0
M25 14 12 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=2.835e-14 PD=8.4e-07 PS=9.1e-07 $X=2485 $Y=870 $D=0
M26 VDD 12 QN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=2825 $Y=680 $D=0
M27 Q 14 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3015 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4 5 6 7
** N=7 EP=7 IP=11 FDC=28
X1 3 4 1 2 5 6 7 DFF_X1 $T=190 0 0 0 $X=75 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_19
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X16
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_21
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN 6 7
** N=9 EP=7 IP=0 FDC=6
M0 9 A1 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 9 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 8 A1 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT MGC_AUTO_NDR_MGC_CLK_NDR_1.0w2.0s_via2_single_MA_north
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4_X1 A4 VDD A3 A2 A1 ZN VSS 8 9
** N=12 EP=9 IP=0 FDC=8
M0 ZN A4 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A3 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A2 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A1 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 10 A4 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 11 A3 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 12 A2 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 ZN A1 12 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FILLCELL_X32
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FA_X1 CO CI B A VDD VSS S 8 9
** N=21 EP=9 IP=0 FDC=28
M0 VSS 10 CO 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 19 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=360 $Y=215 $D=1
M2 10 A 19 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=550 $Y=215 $D=1
M3 11 CI 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07 $X=740 $Y=215 $D=1
M4 VSS A 11 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=935 $Y=215 $D=1
M5 11 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1125 $Y=215 $D=1
M6 13 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1465 $Y=90 $D=1
M7 VSS CI 13 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1655 $Y=90 $D=1
M8 13 A VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1845 $Y=90 $D=1
M9 15 10 13 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07 $X=2035 $Y=90 $D=1
M10 20 CI 15 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07 $X=2235 $Y=90 $D=1
M11 21 B 20 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2425 $Y=90 $D=1
M12 VSS A 21 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=2615 $Y=90 $D=1
M13 S 15 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M14 VDD 10 CO 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M15 16 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=360 $Y=870 $D=0
M16 10 A 16 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=550 $Y=870 $D=0
M17 12 CI 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06 PS=9.1e-07 $X=740 $Y=870 $D=0
M18 VDD A 12 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06 $X=935 $Y=945 $D=0
M19 12 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1125 $Y=945 $D=0
M20 14 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1465 $Y=995 $D=0
M21 VDD CI 14 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1655 $Y=995 $D=0
M22 14 A VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1845 $Y=995 $D=0
M23 15 10 14 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07 $X=2035 $Y=995 $D=0
M24 17 CI 15 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07 $X=2235 $Y=995 $D=0
M25 18 B 17 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2425 $Y=995 $D=0
M26 VDD A 18 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2615 $Y=995 $D=0
M27 S 15 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=14 FDC=56
X0 1 2 3 4 5 9 10 DFF_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 6 7 3 4 8 9 10 DFF_X1 $T=3230 0 0 0 $X=3115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_28
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT INV_X1 A VSS VDD ZN 5 6
** N=6 EP=6 IP=0 FDC=2
M0 ZN A VSS 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI21_X1 B2 B1 ZN A VSS VDD 7 8
** N=10 EP=8 IP=0 FDC=6
M0 10 B2 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN B1 10 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS A ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B2 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 9 B1 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD A 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI21_X1 B2 B1 ZN A VSS VDD 7 8
** N=10 EP=8 IP=0 FDC=6
M0 ZN B2 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 9 B1 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS A 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 10 B2 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M4 ZN B1 10 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M5 VDD A ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT CLKGATETST_X8 SE E CK GCK VSS VDD 7 8
** N=23 EP=8 IP=0 FDC=52
M0 9 SE VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=170 $Y=90 $D=1
M1 VSS E 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=360 $Y=90 $D=1
M2 VSS 12 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.205e-14 PD=8.3e-07 PS=6.3e-07 $X=700 $Y=90 $D=1
M3 18 9 VSS 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=8.3e-07 $X=890 $Y=90 $D=1
M4 13 12 18 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.0125e-14 AS=3.85e-14 PD=8.7e-07 PS=8.3e-07 $X=1080 $Y=90 $D=1
M5 19 10 13 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.0125e-14 PD=4.6e-07 PS=8.7e-07 $X=1290 $Y=160 $D=1
M6 VSS 11 19 7 NMOS_VTL L=5e-08 W=9e-08 AD=3.58e-14 AS=1.26e-14 PD=1.12e-06 PS=4.6e-07 $X=1480 $Y=160 $D=1
M7 11 13 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.58e-14 PD=1.11e-06 PS=1.12e-06 $X=1675 $Y=90 $D=1
M8 VSS 13 11 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1865 $Y=90 $D=1
M9 VSS CK 12 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.69e-14 AS=3.36e-14 PD=1.14e-06 PS=7.4e-07 $X=2260 $Y=90 $D=1
M10 20 CK VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.69e-14 PD=1.11e-06 PS=1.14e-06 $X=2465 $Y=90 $D=1
M11 14 13 20 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2655 $Y=90 $D=1
M12 21 13 14 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2845 $Y=90 $D=1
M13 VSS CK 21 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=3035 $Y=90 $D=1
M14 22 CK VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=3225 $Y=90 $D=1
M15 14 13 22 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=3415 $Y=90 $D=1
M16 23 13 14 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=3605 $Y=90 $D=1
M17 VSS CK 23 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.27e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=3795 $Y=90 $D=1
M18 GCK 14 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.27e-14 PD=6.7e-07 PS=1.11e-06 $X=3985 $Y=90 $D=1
M19 VSS 14 GCK 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=4175 $Y=90 $D=1
M20 GCK 14 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=4365 $Y=90 $D=1
M21 VSS 14 GCK 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=4555 $Y=90 $D=1
M22 GCK 14 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=4745 $Y=90 $D=1
M23 VSS 14 GCK 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=4935 $Y=90 $D=1
M24 GCK 14 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=5125 $Y=90 $D=1
M25 VSS 14 GCK 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=5315 $Y=90 $D=1
M26 15 SE 9 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=170 $Y=995 $D=0
M27 VDD E 15 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=360 $Y=995 $D=0
M28 VDD 12 10 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=3.3075e-14 PD=1.12e-06 PS=8.4e-07 $X=700 $Y=995 $D=0
M29 16 9 VDD 8 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=890 $Y=890 $D=0
M30 13 10 16 8 PMOS_VTL L=5e-08 W=4.2e-07 AD=4.245e-14 AS=5.88e-14 PD=1.16e-06 PS=1.12e-06 $X=1080 $Y=890 $D=0
M31 17 12 13 8 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=4.245e-14 PD=4.6e-07 PS=1.16e-06 $X=1290 $Y=1080 $D=0
M32 VDD 11 17 8 PMOS_VTL L=5e-08 W=9e-08 AD=5.085e-14 AS=1.26e-14 PD=1.55e-06 PS=4.6e-07 $X=1480 $Y=1080 $D=0
M33 11 13 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=5.085e-14 PD=1.54e-06 PS=1.55e-06 $X=1675 $Y=680 $D=0
M34 VDD 13 11 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1865 $Y=680 $D=0
M35 VDD CK 12 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=5.04e-14 PD=1.57e-06 PS=9.5e-07 $X=2260 $Y=790 $D=0
M36 14 CK VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06 PS=1.57e-06 $X=2465 $Y=680 $D=0
M37 VDD 13 14 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2655 $Y=680 $D=0
M38 14 13 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2845 $Y=680 $D=0
M39 VDD CK 14 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3035 $Y=680 $D=0
M40 14 CK VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3225 $Y=680 $D=0
M41 VDD 13 14 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3415 $Y=680 $D=0
M42 14 13 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3605 $Y=680 $D=0
M43 VDD CK 14 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3795 $Y=680 $D=0
M44 GCK 14 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3985 $Y=680 $D=0
M45 VDD 14 GCK 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4175 $Y=680 $D=0
M46 GCK 14 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4365 $Y=680 $D=0
M47 VDD 14 GCK 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4555 $Y=680 $D=0
M48 GCK 14 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4745 $Y=680 $D=0
M49 VDD 14 GCK 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4935 $Y=680 $D=0
M50 GCK 14 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=5125 $Y=680 $D=0
M51 VDD 14 GCK 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=5315 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2_X1 VSS A ZN B VDD 6 7
** N=11 EP=7 IP=0 FDC=10
M0 11 A 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=155 $Y=90 $D=1
M1 VSS B 11 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=345 $Y=90 $D=1
M2 9 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=540 $Y=90 $D=1
M3 ZN A 9 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 9 B ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 8 A VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=155 $Y=995 $D=0
M6 VDD B 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=345 $Y=995 $D=0
M7 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=540 $Y=680 $D=0
M8 10 A ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M9 VDD B 10 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_31
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT NOR2_X1 A2 VDD A1 ZN VSS 6 7
** N=8 EP=7 IP=0 FDC=4
M0 ZN A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A1 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 8 A2 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 ZN A1 8 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND3_X1 A3 VSS A2 A1 VDD ZN 7 8
** N=10 EP=8 IP=0 FDC=6
M0 9 A3 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 10 A2 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 10 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A3 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 VDD A2 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND2_X1 A2 VSS A1 ZN VDD 6 7
** N=8 EP=7 IP=0 FDC=4
M0 8 A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN A1 8 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A2 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A1 ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI211_X1 C2 C1 B VSS A ZN VDD 8 9
** N=12 EP=9 IP=0 FDC=8
M0 12 C2 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN C1 12 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS B ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN A VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 ZN C2 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 10 C1 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 11 B 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT HA_X1 S B A VSS VDD CO 7 8
** N=14 EP=8 IP=0 FDC=16
M0 13 B VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 S A 13 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 10 S 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.48e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 10 B VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.48e-14 PD=7e-07 PS=1.12e-06 $X=760 $Y=90 $D=1
M4 VSS A 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=950 $Y=90 $D=1
M5 14 A 11 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1320 $Y=90 $D=1
M6 VSS B 14 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=1510 $Y=90 $D=1
M7 CO 11 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1700 $Y=90 $D=1
M8 S B 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 9 A S 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 VDD 10 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.7725e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 12 B VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.7725e-14 PD=9.1e-07 PS=1.55e-06 $X=760 $Y=870 $D=0
M12 10 A 12 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=950 $Y=870 $D=0
M13 11 A VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1320 $Y=870 $D=0
M14 VDD B 11 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=1510 $Y=870 $D=0
M15 CO 11 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1700 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT CLKBUF_X3 A VSS VDD Z 5 6
** N=7 EP=6 IP=0 FDC=8
M0 VSS A 7 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=145 $Y=90 $D=1
M1 Z 7 VSS 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=335 $Y=90 $D=1
M2 VSS 7 Z 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=525 $Y=90 $D=1
M3 Z 7 VSS 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=715 $Y=90 $D=1
M4 VDD A 7 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 Z 7 VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 VDD 7 Z 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 Z 7 VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT via1_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT OR2_X1 A1 A2 VSS VDD ZN 6 7
** N=9 EP=7 IP=0 FDC=6
M0 8 A1 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 9 A1 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 9 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_34
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFFR_X1 CK D RN VSS VDD Q 7 8
** N=25 EP=8 IP=0 FDC=32
M0 VSS CK 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=140 $D=1
M1 13 9 VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=335 $Y=140 $D=1
M2 20 D VSS 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=2.8875e-14 PD=8.3e-07 PS=7.6e-07 $X=675 $Y=215 $D=1
M3 10 9 20 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=2.555e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=865 $Y=215 $D=1
M4 21 13 10 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.555e-14 PD=4.6e-07 PS=8.3e-07 $X=1055 $Y=305 $D=1
M5 22 12 21 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=1245 $Y=305 $D=1
M6 VSS RN 22 7 NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14 PD=3.9e-07 PS=4.6e-07 $X=1435 $Y=305 $D=1
M7 VSS 10 12 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.41e-14 AS=2.205e-14 PD=8.4e-07 PS=6.3e-07 $X=1790 $Y=215 $D=1
M8 23 10 VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.41e-14 PD=7e-07 PS=8.4e-07 $X=2050 $Y=215 $D=1
M9 14 13 23 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2240 $Y=215 $D=1
M10 24 9 14 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=2430 $Y=215 $D=1
M11 VSS 16 24 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.26e-14 PD=7e-07 PS=4.6e-07 $X=2620 $Y=215 $D=1
M12 25 RN VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.1e-14 PD=7e-07 PS=7e-07 $X=2810 $Y=215 $D=1
M13 16 14 25 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=3000 $Y=215 $D=1
M14 VSS 14 QN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=3385 $Y=90 $D=1
M15 Q 16 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=3575 $Y=90 $D=1
M16 VDD CK 9 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M17 13 9 VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M18 17 D VDD 8 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=4.41e-14 PD=1.12e-06 PS=1.05e-06 $X=675 $Y=840 $D=0
M19 10 13 17 8 PMOS_VTL L=5e-08 W=4.2e-07 AD=3.57e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=865 $Y=840 $D=0
M20 11 9 10 8 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.57e-14 PD=4.6e-07 PS=1.12e-06 $X=1055 $Y=1020 $D=0
M21 VDD 12 11 8 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=1245 $Y=1020 $D=0
M22 11 RN VDD 8 PMOS_VTL L=5e-08 W=9e-08 AD=1.035e-14 AS=1.26e-14 PD=4.1e-07 PS=4.6e-07 $X=1435 $Y=1020 $D=0
M23 VDD 10 12 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.465e-14 PD=1.05e-06 PS=8.5e-07 $X=1790 $Y=855 $D=0
M24 18 10 VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.05e-06 $X=2050 $Y=855 $D=0
M25 14 9 18 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2240 $Y=855 $D=0
M26 19 13 14 8 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=2430 $Y=995 $D=0
M27 VDD 16 19 8 PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.26e-14 PD=9.1e-07 PS=4.6e-07 $X=2620 $Y=995 $D=0
M28 16 RN VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=2.835e-14 PD=9.1e-07 PS=9.1e-07 $X=2810 $Y=995 $D=0
M29 VDD 14 16 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=3000 $Y=995 $D=0
M30 VDD 14 QN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=3385 $Y=680 $D=0
M31 Q 16 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3575 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI22_X1 B2 B1 VDD A1 ZN A2 VSS 8 9
** N=12 EP=9 IP=0 FDC=8
M0 11 B2 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN B1 11 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 12 A1 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 VSS A2 12 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 VDD B2 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 10 B1 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 ZN A1 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 10 A2 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS 6 7
** N=11 EP=7 IP=0 FDC=10
M0 8 A VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 11 A Z 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 11 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 10 A 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 10 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 9 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 9 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 9 B Z 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUF_X1 A VSS VDD Z 5 6
** N=7 EP=6 IP=0 FDC=4
M0 VSS A 7 5 NMOS_VTL L=5e-08 W=9.5e-08 AD=2.03e-14 AS=9.975e-15 PD=6.7e-07 PS=4e-07 $X=165 $Y=160 $D=1
M1 Z 7 VSS 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.03e-14 PD=6e-07 PS=6.7e-07 $X=355 $Y=160 $D=1
M2 VDD A 7 6 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=165 $Y=995 $D=0
M3 Z 7 VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=355 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI22_X1 B2 B1 VSS ZN A1 A2 VDD 8 9
** N=12 EP=9 IP=0 FDC=8
M0 VSS B2 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 10 B1 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A1 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 10 A2 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 11 B2 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 ZN B1 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 12 A1 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 VDD A2 12 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR3_X1 A1 A2 A3 VSS VDD ZN 7 8
** N=11 EP=8 IP=0 FDC=8
M0 VSS A1 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 9 A2 VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 VSS A3 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=525 $Y=90 $D=1
M3 ZN 9 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 10 A1 9 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M5 11 A2 10 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M6 VDD A3 11 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=525 $Y=995 $D=0
M7 ZN 9 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR3_X1 A3 VDD A2 A1 VSS ZN 7 8
** N=10 EP=8 IP=0 FDC=6
M0 ZN A3 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A2 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 9 A3 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 10 A2 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 10 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT fp_mul
** N=668 EP=0 IP=11415 FDC=7576
M0 205 171 171 634 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=5325 $Y=34690 $D=1
M1 171 204 205 634 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=5515 $Y=34690 $D=1
M2 171 215 209 634 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.205e-14 PD=8.3e-07 PS=6.3e-07 $X=5855 $Y=34690 $D=1
M3 628 205 171 634 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=8.3e-07 $X=6045 $Y=34690 $D=1
M4 217 215 628 634 NMOS_VTL L=5e-08 W=2.75e-07 AD=2.555e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=6235 $Y=34690 $D=1
M5 629 209 217 634 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.555e-14 PD=4.6e-07 PS=8.3e-07 $X=6425 $Y=34765 $D=1
M6 171 214 629 634 NMOS_VTL L=5e-08 W=9e-08 AD=3.58e-14 AS=1.26e-14 PD=1.12e-06 PS=4.6e-07 $X=6615 $Y=34765 $D=1
M7 214 217 171 634 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=3.58e-14 PD=1.04e-06 PS=1.12e-06 $X=6810 $Y=34690 $D=1
M8 171 1 215 634 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.69e-14 AS=2.31e-14 PD=1.14e-06 PS=6.4e-07 $X=7210 $Y=34690 $D=1
M9 630 1 171 634 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.69e-14 PD=1.11e-06 PS=1.14e-06 $X=7415 $Y=34690 $D=1
M10 219 217 630 634 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7605 $Y=34690 $D=1
M11 631 217 219 634 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7795 $Y=34690 $D=1
M12 171 1 631 634 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.27e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7985 $Y=34690 $D=1
M13 223 219 171 634 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.27e-14 PD=6.7e-07 PS=1.11e-06 $X=8175 $Y=34690 $D=1
M14 171 219 223 634 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=8365 $Y=34690 $D=1
M15 223 219 171 634 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=8555 $Y=34690 $D=1
M16 171 219 223 634 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=8745 $Y=34690 $D=1
M17 632 232 171 635 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=14825 $Y=11695 $D=1
M18 241 59 632 635 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=15015 $Y=11695 $D=1
M19 171 63 241 635 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=15205 $Y=11695 $D=1
M20 633 67 171 635 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=15395 $Y=11695 $D=1
M21 241 239 633 635 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=15585 $Y=11695 $D=1
M22 10 279 171 636 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=35915 $Y=14495 $D=1
M23 171 278 10 636 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=36105 $Y=14495 $D=1
M24 10 278 171 636 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=36295 $Y=14495 $D=1
M25 171 279 10 636 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=36485 $Y=14495 $D=1
M26 623 171 205 652 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=5325 $Y=35595 $D=0
M27 203 204 623 652 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=5515 $Y=35595 $D=0
M28 203 215 209 652 PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=3.3075e-14 PD=1.12e-06 PS=8.4e-07 $X=5855 $Y=35520 $D=0
M29 624 205 203 652 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=6045 $Y=35490 $D=0
M30 217 209 624 652 PMOS_VTL L=5e-08 W=4.2e-07 AD=3.6075e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=6235 $Y=35490 $D=0
M31 625 215 217 652 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.6075e-14 PD=4.6e-07 PS=1.12e-06 $X=6425 $Y=35745 $D=0
M32 203 214 625 652 PMOS_VTL L=5e-08 W=9e-08 AD=5.085e-14 AS=1.26e-14 PD=1.55e-06 PS=4.6e-07 $X=6615 $Y=35745 $D=0
M33 214 217 203 652 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=5.085e-14 PD=1.47e-06 PS=1.55e-06 $X=6810 $Y=35280 $D=0
M34 203 1 215 652 PMOS_VTL L=5e-08 W=3.15e-07 AD=7.5425e-14 AS=4.5675e-14 PD=1.57e-06 PS=9.2e-07 $X=7210 $Y=35465 $D=0
M35 219 1 203 652 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=7.5425e-14 PD=1.54e-06 PS=1.57e-06 $X=7415 $Y=35280 $D=0
M36 203 217 219 652 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7605 $Y=35280 $D=0
M37 219 217 203 652 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7795 $Y=35280 $D=0
M38 203 1 219 652 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7985 $Y=35280 $D=0
M39 223 219 203 652 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=8175 $Y=35280 $D=0
M40 203 219 223 652 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=8365 $Y=35280 $D=0
M41 223 219 203 652 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=8555 $Y=35280 $D=0
M42 203 219 223 652 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=8745 $Y=35280 $D=0
M43 203 232 235 653 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=14825 $Y=10890 $D=0
M44 235 59 203 653 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=15015 $Y=10890 $D=0
M45 240 63 235 653 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=15205 $Y=10890 $D=0
M46 241 67 240 653 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=15395 $Y=10890 $D=0
M47 240 239 241 653 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=15585 $Y=10890 $D=0
M48 626 279 203 654 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=35915 $Y=13690 $D=0
M49 10 278 626 654 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=36105 $Y=13690 $D=0
M50 627 278 10 654 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=36295 $Y=13690 $D=0
M51 203 279 627 654 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=36485 $Y=13690 $D=0
X4452 6 245 7 171 203 532 650 665 MUX2_X1 $T=4230 43000 1 0 $X=4115 $Y=41485
X4453 411 245 8 171 203 291 646 662 MUX2_X1 $T=4230 45800 1 0 $X=4115 $Y=44285
X4454 17 245 13 171 203 478 635 654 MUX2_X1 $T=7460 12200 1 180 $X=6015 $Y=12085
X4455 14 245 18 171 203 533 643 664 MUX2_X1 $T=6320 26200 1 0 $X=6205 $Y=24685
X4456 480 245 20 171 203 24 640 657 MUX2_X1 $T=6510 29000 1 0 $X=6395 $Y=27485
X4457 16 245 21 171 203 534 648 660 MUX2_X1 $T=6700 17800 1 0 $X=6585 $Y=16285
X4458 23 245 27 171 203 39 635 653 MUX2_X1 $T=7460 12200 1 0 $X=7345 $Y=10685
X4459 28 245 33 171 203 421 636 660 MUX2_X1 $T=8030 15000 0 0 $X=7915 $Y=14885
X4460 34 245 30 171 203 210 642 658 MUX2_X1 $T=9360 23400 0 180 $X=7915 $Y=21885
X4461 35 245 31 171 203 218 650 662 MUX2_X1 $T=9360 43000 1 180 $X=7915 $Y=42885
X4462 41 245 44 171 203 314 636 654 MUX2_X1 $T=10120 15000 1 0 $X=10005 $Y=13485
X4463 46 245 49 171 203 535 650 662 MUX2_X1 $T=11070 43000 0 0 $X=10955 $Y=42885
X4464 66 245 62 171 203 506 650 665 MUX2_X1 $T=15440 43000 0 180 $X=13995 $Y=41485
X4465 73 245 64 171 203 433 636 660 MUX2_X1 $T=16010 15000 1 180 $X=14565 $Y=14885
X4466 80 245 82 171 203 342 638 656 MUX2_X1 $T=17150 40200 1 0 $X=17035 $Y=38685
X4467 85 245 87 171 203 94 640 667 MUX2_X1 $T=18480 29000 0 0 $X=18365 $Y=28885
X4468 88 245 92 171 203 511 646 662 MUX2_X1 $T=19050 45800 1 0 $X=18935 $Y=44285
X4469 100 245 96 171 203 91 648 660 MUX2_X1 $T=21710 17800 0 180 $X=20265 $Y=16285
X4470 102 245 105 171 203 512 638 656 MUX2_X1 $T=21710 40200 1 0 $X=21595 $Y=38685
X4471 356 245 107 171 203 353 635 654 MUX2_X1 $T=22090 12200 0 0 $X=21975 $Y=12085
X4472 108 245 113 171 203 536 640 667 MUX2_X1 $T=23040 29000 0 0 $X=22925 $Y=28885
X4473 118 245 120 171 203 123 650 662 MUX2_X1 $T=23990 43000 0 0 $X=23875 $Y=42885
X4474 133 245 128 171 203 537 646 668 MUX2_X1 $T=28170 45800 1 180 $X=26725 $Y=45685
X4475 137 245 139 171 203 516 650 665 MUX2_X1 $T=27980 43000 1 0 $X=27865 $Y=41485
X4476 140 245 142 171 203 144 648 660 MUX2_X1 $T=28740 17800 1 0 $X=28625 $Y=16285
X4477 145 245 141 171 203 135 641 652 MUX2_X1 $T=30070 37400 0 180 $X=28625 $Y=35885
X4478 370 245 143 171 203 538 636 654 MUX2_X1 $T=28930 15000 1 0 $X=28815 $Y=13485
X4479 147 245 148 171 203 539 646 668 MUX2_X1 $T=29880 45800 0 0 $X=29765 $Y=45685
X4480 158 245 155 171 203 540 638 665 MUX2_X1 $T=34820 40200 1 180 $X=33375 $Y=40085
X4481 159 245 276 171 203 541 638 665 MUX2_X1 $T=34820 40200 0 0 $X=34705 $Y=40085
X4482 381 161 160 171 203 542 648 663 MUX2_X1 $T=35200 17800 0 0 $X=35085 $Y=17685
X4483 162 245 166 171 203 165 634 659 MUX2_X1 $T=36530 34600 1 0 $X=36415 $Y=33085
X4484 168 245 167 171 203 530 646 662 MUX2_X1 $T=38810 45800 0 180 $X=37365 $Y=44285
X4485 173 245 175 171 203 543 646 668 MUX2_X1 $T=39380 45800 0 0 $X=39265 $Y=45685
X4486 179 245 176 171 203 522 650 665 MUX2_X1 $T=41660 43000 0 180 $X=40215 $Y=41485
X4487 177 245 181 171 203 282 643 664 MUX2_X1 $T=41090 26200 1 0 $X=40975 $Y=24685
X4488 178 245 182 171 203 544 647 667 MUX2_X1 $T=41090 31800 1 0 $X=40975 $Y=30285
X4489 183 245 180 171 203 469 641 652 MUX2_X1 $T=42420 37400 0 180 $X=40975 $Y=35885
X4490 184 245 188 171 203 397 646 662 MUX2_X1 $T=42040 45800 1 0 $X=41925 $Y=44285
X4491 187 245 190 171 203 284 634 652 MUX2_X1 $T=42610 34600 0 0 $X=42495 $Y=34485
X4492 191 245 189 171 203 395 640 667 MUX2_X1 $T=44320 29000 1 180 $X=42875 $Y=28885
X4493 197 245 194 171 203 473 642 664 MUX2_X1 $T=45080 23400 1 180 $X=43635 $Y=23285
X4494 192 245 195 171 203 531 641 656 MUX2_X1 $T=43750 37400 0 0 $X=43635 $Y=37285
X4495 193 245 196 171 203 545 650 665 MUX2_X1 $T=43750 43000 1 0 $X=43635 $Y=41485
X4496 198 245 200 171 203 406 643 657 MUX2_X1 $T=46980 26200 0 0 $X=46865 $Y=26085
X4497 201 245 199 171 203 496 650 662 MUX2_X1 $T=48310 43000 1 180 $X=46865 $Y=42885
X5337 564 3 171 203 44 635 653 DFF_X1 $T=1000 12200 1 0 $X=885 $Y=10685
X5338 565 3 171 203 13 635 654 DFF_X1 $T=1000 12200 0 0 $X=885 $Y=12085
X5339 566 3 171 203 64 636 660 DFF_X1 $T=1000 15000 0 0 $X=885 $Y=14885
X5340 567 3 171 203 21 648 660 DFF_X1 $T=1000 17800 1 0 $X=885 $Y=16285
X5341 318 2 171 203 409 645 658 DFF_X1 $T=1000 20600 0 0 $X=885 $Y=20485
X5342 568 3 171 203 30 642 658 DFF_X1 $T=1000 23400 1 0 $X=885 $Y=21885
X5343 569 3 171 203 18 642 664 DFF_X1 $T=1000 23400 0 0 $X=885 $Y=23285
X5344 315 2 171 203 477 643 664 DFF_X1 $T=1000 26200 1 0 $X=885 $Y=24685
X5345 551 2 171 203 288 640 657 DFF_X1 $T=1000 29000 1 0 $X=885 $Y=27485
X5346 301 2 171 203 410 640 667 DFF_X1 $T=1000 29000 0 0 $X=885 $Y=28885
X5347 299 2 171 203 289 634 659 DFF_X1 $T=1000 34600 1 0 $X=885 $Y=33085
X5348 570 3 171 203 7 638 665 DFF_X1 $T=1000 40200 0 0 $X=885 $Y=40085
X5349 532 4 171 203 6 650 665 DFF_X1 $T=1000 43000 1 0 $X=885 $Y=41485
X5350 291 4 171 203 411 646 662 DFF_X1 $T=1000 45800 1 0 $X=885 $Y=44285
X5351 571 3 171 203 8 651 668 DFF_X1 $T=1000 48600 1 0 $X=885 $Y=47085
X5352 572 3 171 203 27 637 653 DFF_X1 $T=1950 9400 0 0 $X=1835 $Y=9285
X5353 478 4 171 203 17 636 654 DFF_X1 $T=5560 15000 1 0 $X=5445 $Y=13485
X5354 218 4 171 203 35 646 662 DFF_X1 $T=5560 45800 1 0 $X=5445 $Y=44285
X5355 24 4 171 203 480 643 657 DFF_X1 $T=6890 26200 0 0 $X=6775 $Y=26085
X5356 533 4 171 203 14 642 664 DFF_X1 $T=7270 23400 0 0 $X=7155 $Y=23285
X5357 534 4 171 203 16 648 663 DFF_X1 $T=7460 17800 0 0 $X=7345 $Y=17685
X5358 529 2 171 203 305 647 667 DFF_X1 $T=11450 31800 0 180 $X=8105 $Y=30285
X5359 432 2 171 203 419 647 659 DFF_X1 $T=11830 31800 1 180 $X=8485 $Y=31685
X5360 39 4 171 203 23 635 653 DFF_X1 $T=8790 12200 1 0 $X=8675 $Y=10685
X5361 421 4 171 203 28 636 660 DFF_X1 $T=9360 15000 0 0 $X=9245 $Y=14885
X5362 505 2 171 203 507 649 661 DFF_X1 $T=11260 1000 0 0 $X=11145 $Y=885
X5363 314 4 171 203 41 636 654 DFF_X1 $T=11450 15000 1 0 $X=11335 $Y=13485
X5364 577 3 171 203 87 640 667 DFF_X1 $T=11830 29000 0 0 $X=11715 $Y=28885
X5365 506 4 171 203 66 638 665 DFF_X1 $T=12970 40200 0 0 $X=12855 $Y=40085
X5366 510 2 171 203 610 649 661 DFF_X1 $T=17720 1000 1 180 $X=14375 $Y=885
X5367 247 3 171 203 96 644 661 DFF_X1 $T=16390 3800 1 0 $X=16275 $Y=2285
X5368 342 4 171 203 80 638 656 DFF_X1 $T=18480 40200 1 0 $X=18365 $Y=38685
X5369 91 4 171 203 100 648 663 DFF_X1 $T=19050 17800 0 0 $X=18935 $Y=17685
X5370 94 4 171 203 85 640 667 DFF_X1 $T=19810 29000 0 0 $X=19695 $Y=28885
X5371 581 3 171 203 107 639 655 DFF_X1 $T=21140 6600 0 0 $X=21025 $Y=6485
X5372 537 4 171 203 88 646 662 DFF_X1 $T=22090 45800 1 0 $X=21975 $Y=44285
X5373 512 4 171 203 102 641 656 DFF_X1 $T=23040 37400 0 0 $X=22925 $Y=37285
X5374 353 4 171 203 356 635 654 DFF_X1 $T=23420 12200 0 0 $X=23305 $Y=12085
X5375 125 2 171 203 354 641 652 DFF_X1 $T=26840 37400 0 180 $X=23495 $Y=35885
X5376 528 3 171 203 363 644 666 DFF_X1 $T=23990 3800 0 0 $X=23875 $Y=3685
X5377 122 3 171 203 143 637 653 DFF_X1 $T=24370 9400 0 0 $X=24255 $Y=9285
X5378 452 2 171 203 515 649 661 DFF_X1 $T=24560 1000 0 0 $X=24445 $Y=885
X5379 123 4 171 203 137 650 665 DFF_X1 $T=24750 43000 1 0 $X=24635 $Y=41485
X5380 262 3 171 203 139 650 662 DFF_X1 $T=25320 43000 0 0 $X=25205 $Y=42885
X5381 611 3 171 203 153 637 655 DFF_X1 $T=25890 9400 1 0 $X=25775 $Y=7885
X5382 134 3 171 203 375 644 666 DFF_X1 $T=27220 3800 0 0 $X=27105 $Y=3685
X5383 135 4 171 203 145 641 656 DFF_X1 $T=27220 37400 0 0 $X=27105 $Y=37285
X5384 138 3 171 203 371 644 661 DFF_X1 $T=27790 3800 1 0 $X=27675 $Y=2285
X5385 266 2 171 203 489 634 652 DFF_X1 $T=31210 34600 1 180 $X=27865 $Y=34485
X5386 490 115 171 203 151 640 657 DFF_X1 $T=28360 29000 1 0 $X=28245 $Y=27485
X5387 516 4 171 203 127 638 656 DFF_X1 $T=28550 40200 1 0 $X=28435 $Y=38685
X5388 144 4 171 203 140 645 663 DFF_X1 $T=28930 20600 1 0 $X=28815 $Y=19085
X5389 268 3 171 203 155 650 665 DFF_X1 $T=29310 43000 1 0 $X=29195 $Y=41485
X5390 517 115 171 203 164 642 658 DFF_X1 $T=29500 23400 1 0 $X=29385 $Y=21885
X5391 149 3 171 203 166 641 652 DFF_X1 $T=30070 37400 1 0 $X=29955 $Y=35885
X5392 606 3 171 203 378 636 654 DFF_X1 $T=30260 15000 1 0 $X=30145 $Y=13485
X5393 559 4 171 203 162 634 659 DFF_X1 $T=30640 34600 1 0 $X=30525 $Y=33085
X5394 540 4 171 203 159 638 656 DFF_X1 $T=31780 40200 1 0 $X=31665 $Y=38685
X5395 519 115 171 203 379 645 663 DFF_X1 $T=32160 20600 1 0 $X=32045 $Y=19085
X5396 274 2 171 203 373 635 653 DFF_X1 $T=35580 12200 0 180 $X=32235 $Y=10685
X5397 469 4 171 203 158 641 652 DFF_X1 $T=33300 37400 1 0 $X=33185 $Y=35885
X5398 530 4 171 203 147 646 662 DFF_X1 $T=37480 45800 0 180 $X=34135 $Y=44285
X5399 165 4 171 203 177 640 667 DFF_X1 $T=36530 29000 0 0 $X=36415 $Y=28885
X5400 543 4 171 203 168 650 665 DFF_X1 $T=37100 43000 1 0 $X=36985 $Y=41485
X5401 369 2 171 203 390 643 664 DFF_X1 $T=37860 26200 1 0 $X=37745 $Y=24685
X5402 281 3 171 203 185 637 653 DFF_X1 $T=38050 9400 0 0 $X=37935 $Y=9285
X5403 382 2 171 203 562 647 659 DFF_X1 $T=38620 31800 0 0 $X=38505 $Y=31685
X5404 589 3 171 203 275 637 655 DFF_X1 $T=38810 9400 1 0 $X=38695 $Y=7885
X5405 397 4 171 203 173 646 662 DFF_X1 $T=42040 45800 0 180 $X=38695 $Y=44285
X5406 395 4 171 203 178 640 667 DFF_X1 $T=42990 29000 1 180 $X=39645 $Y=28885
X5407 560 2 171 203 494 648 660 DFF_X1 $T=40520 17800 1 0 $X=40405 $Y=16285
X5408 531 4 171 203 183 641 656 DFF_X1 $T=43750 37400 1 180 $X=40405 $Y=37285
X5409 544 4 171 203 187 647 659 DFF_X1 $T=41850 31800 0 0 $X=41735 $Y=31685
X5410 592 3 171 203 188 651 668 DFF_X1 $T=41850 48600 1 0 $X=41735 $Y=47085
X5411 545 4 171 203 201 650 662 DFF_X1 $T=43750 43000 0 0 $X=43635 $Y=42885
X5412 563 2 171 203 474 649 661 DFF_X1 $T=45080 1000 0 0 $X=44965 $Y=885
X5413 593 3 171 203 497 644 666 DFF_X1 $T=45080 3800 0 0 $X=44965 $Y=3685
X5414 398 2 171 203 475 639 655 DFF_X1 $T=45080 6600 0 0 $X=44965 $Y=6485
X5415 594 3 171 203 396 637 655 DFF_X1 $T=45080 9400 1 0 $X=44965 $Y=7885
X5416 399 2 171 203 525 635 654 DFF_X1 $T=45080 12200 0 0 $X=44965 $Y=12085
X5417 596 3 171 203 476 636 660 DFF_X1 $T=45080 15000 0 0 $X=44965 $Y=14885
X5418 401 2 171 203 404 648 663 DFF_X1 $T=45080 17800 0 0 $X=44965 $Y=17685
X5419 609 3 171 203 181 642 664 DFF_X1 $T=45080 23400 0 0 $X=44965 $Y=23285
X5420 598 3 171 203 182 647 667 DFF_X1 $T=45080 31800 1 0 $X=44965 $Y=30285
X5421 599 3 171 203 189 647 659 DFF_X1 $T=45080 31800 0 0 $X=44965 $Y=31685
X5422 600 3 171 203 190 634 659 DFF_X1 $T=45080 34600 1 0 $X=44965 $Y=33085
X5423 601 3 171 203 180 641 652 DFF_X1 $T=45080 37400 1 0 $X=44965 $Y=35885
X5424 602 3 171 203 195 641 656 DFF_X1 $T=45080 37400 0 0 $X=44965 $Y=37285
X5425 604 3 171 203 176 650 665 DFF_X1 $T=45080 43000 1 0 $X=44965 $Y=41485
X5426 496 4 171 203 184 646 662 DFF_X1 $T=48310 45800 0 180 $X=44965 $Y=44285
X5427 605 3 171 203 199 651 668 DFF_X1 $T=45080 48600 1 0 $X=44965 $Y=47085
X5630 171 203 573 3 33 648 663 ICV_18 $T=4040 17800 0 0 $X=3925 $Y=17685
X5631 171 203 574 3 20 647 667 ICV_18 $T=4040 31800 1 0 $X=3925 $Y=30285
X5632 171 203 535 4 46 650 665 ICV_18 $T=10690 43000 1 0 $X=10575 $Y=41485
X5633 171 203 578 3 62 646 662 ICV_18 $T=12970 45800 1 0 $X=12855 $Y=44285
X5634 171 203 433 4 73 648 660 ICV_18 $T=14110 17800 1 0 $X=13995 $Y=16285
X5635 171 203 579 3 79 651 668 ICV_18 $T=14490 48600 1 0 $X=14375 $Y=47085
X5636 171 203 557 2 257 649 661 ICV_18 $T=21140 1000 0 0 $X=21025 $Y=885
X5637 171 203 582 3 141 638 665 ICV_18 $T=24180 40200 0 0 $X=24065 $Y=40085
X5638 171 203 536 4 108 640 657 ICV_18 $T=24940 29000 1 0 $X=24825 $Y=27485
X5639 171 203 459 4 154 647 659 ICV_18 $T=30260 31800 0 0 $X=30145 $Y=31685
X5640 171 203 376 115 152 640 667 ICV_18 $T=30830 29000 0 0 $X=30715 $Y=28885
X5641 171 203 542 115 381 648 663 ICV_18 $T=31780 17800 0 0 $X=31665 $Y=17685
X5642 171 203 520 1 163 642 658 ICV_18 $T=38430 23400 1 0 $X=38315 $Y=21885
X5643 171 203 541 4 179 638 656 ICV_18 $T=38430 40200 1 0 $X=38315 $Y=38685
X5644 171 203 284 4 192 634 652 ICV_18 $T=39190 34600 0 0 $X=39075 $Y=34485
X5645 171 203 386 2 283 645 658 ICV_18 $T=39950 20600 0 0 $X=39835 $Y=20485
X5646 171 203 473 4 198 643 657 ICV_18 $T=43560 26200 0 0 $X=43445 $Y=26085
X5647 171 203 595 3 403 637 653 ICV_18 $T=44890 9400 0 0 $X=44775 $Y=9285
X5648 171 203 393 2 405 645 663 ICV_18 $T=44890 20600 1 0 $X=44775 $Y=19085
X5926 40 10 171 203 292 644 661 AND2_X1 $T=6320 3800 0 180 $X=5445 $Y=2285
X5927 29 10 171 203 296 634 659 AND2_X1 $T=5560 34600 1 0 $X=5445 $Y=33085
X5928 233 11 171 203 413 639 666 AND2_X1 $T=6510 6600 0 180 $X=5635 $Y=5085
X5929 233 12 171 203 302 641 656 AND2_X1 $T=6130 37400 0 0 $X=6015 $Y=37285
X5930 12 10 171 203 547 634 659 AND2_X1 $T=6320 34600 1 0 $X=6205 $Y=33085
X5931 233 15 171 203 304 639 666 AND2_X1 $T=6510 6600 1 0 $X=6395 $Y=5085
X5932 15 10 171 203 415 644 666 AND2_X1 $T=6700 3800 0 0 $X=6585 $Y=3685
X5933 32 10 171 203 301 647 667 AND2_X1 $T=8220 31800 0 180 $X=7345 $Y=30285
X5934 233 29 171 203 227 641 656 AND2_X1 $T=8030 37400 0 0 $X=7915 $Y=37285
X5935 233 32 171 203 37 634 659 AND2_X1 $T=8980 34600 0 180 $X=8105 $Y=33085
X5936 216 37 171 203 308 634 659 AND2_X1 $T=8980 34600 1 0 $X=8865 $Y=33085
X5937 72 10 171 203 310 634 659 AND2_X1 $T=10500 34600 0 180 $X=9625 $Y=33085
X5938 233 40 171 203 226 639 666 AND2_X1 $T=9930 6600 1 0 $X=9815 $Y=5085
X5939 45 10 171 203 312 645 663 AND2_X1 $T=10880 20600 0 180 $X=10005 $Y=19085
X5940 52 10 171 203 551 643 657 AND2_X1 $T=10880 26200 1 180 $X=10005 $Y=26085
X5941 43 10 171 203 315 643 664 AND2_X1 $T=10690 26200 1 0 $X=10575 $Y=24685
X5942 233 45 171 203 228 645 658 AND2_X1 $T=11640 20600 1 180 $X=10765 $Y=20485
X5943 74 10 171 203 48 645 663 AND2_X1 $T=12780 20600 0 180 $X=11905 $Y=19085
X5944 233 52 171 203 320 643 657 AND2_X1 $T=12590 26200 0 0 $X=12475 $Y=26085
X5945 55 10 171 203 431 644 661 AND2_X1 $T=14110 3800 0 180 $X=13235 $Y=2285
X5946 233 55 171 203 232 639 655 AND2_X1 $T=13350 6600 0 0 $X=13235 $Y=6485
X5947 328 10 171 203 432 647 659 AND2_X1 $T=13350 31800 0 0 $X=13235 $Y=31685
X5948 233 328 171 203 321 634 659 AND2_X1 $T=14110 34600 0 180 $X=13235 $Y=33085
X5949 233 72 171 203 78 634 659 AND2_X1 $T=15250 34600 1 0 $X=15135 $Y=33085
X5950 233 74 171 203 326 645 663 AND2_X1 $T=16200 20600 0 180 $X=15325 $Y=19085
X5951 75 10 171 203 616 644 661 AND2_X1 $T=15630 3800 1 0 $X=15515 $Y=2285
X5952 233 75 171 203 336 639 666 AND2_X1 $T=15630 6600 1 0 $X=15515 $Y=5085
X5953 243 78 171 203 335 634 659 AND2_X1 $T=16770 34600 0 180 $X=15895 $Y=33085
X5954 90 10 171 203 529 647 667 AND2_X1 $T=16200 31800 1 0 $X=16085 $Y=30285
X5955 245 79 171 203 206 646 662 AND2_X1 $T=17150 45800 0 180 $X=16275 $Y=44285
X5956 233 43 171 203 83 643 657 AND2_X1 $T=17530 26200 0 0 $X=17415 $Y=26085
X5957 341 83 171 203 439 643 664 AND2_X1 $T=17910 26200 1 0 $X=17795 $Y=24685
X5958 233 90 171 203 252 647 659 AND2_X1 $T=19430 31800 0 0 $X=19315 $Y=31685
X5959 233 95 171 203 248 639 655 AND2_X1 $T=21140 6600 1 180 $X=20265 $Y=6485
X5960 95 10 171 203 449 644 666 AND2_X1 $T=21520 3800 0 0 $X=21405 $Y=3685
X5961 233 103 171 203 249 635 653 AND2_X1 $T=22660 12200 0 180 $X=21785 $Y=10685
X5962 233 104 171 203 106 636 660 AND2_X1 $T=22090 15000 0 0 $X=21975 $Y=14885
X5963 348 106 171 203 450 648 660 AND2_X1 $T=22280 17800 1 0 $X=22165 $Y=16285
X5964 104 10 171 203 357 637 653 AND2_X1 $T=23610 9400 0 0 $X=23495 $Y=9285
X5965 103 10 171 203 259 639 666 AND2_X1 $T=23990 6600 1 0 $X=23875 $Y=5085
X5966 233 121 171 203 116 634 652 AND2_X1 $T=25320 34600 1 180 $X=24445 $Y=34485
X5967 121 10 171 203 125 634 652 AND2_X1 $T=26650 34600 1 180 $X=25775 $Y=34485
X5968 233 127 171 203 224 641 656 AND2_X1 $T=26270 37400 0 0 $X=26155 $Y=37285
X5969 233 129 171 203 453 648 660 AND2_X1 $T=27790 17800 0 180 $X=26915 $Y=16285
X5970 233 131 171 203 126 642 658 AND2_X1 $T=27980 23400 0 180 $X=27105 $Y=21885
X5971 233 132 171 203 364 643 664 AND2_X1 $T=27980 26200 0 180 $X=27105 $Y=24685
X5972 233 136 171 203 367 647 659 AND2_X1 $T=28550 31800 1 180 $X=27675 $Y=31685
X5973 129 10 171 203 368 636 654 AND2_X1 $T=28170 15000 1 0 $X=28055 $Y=13485
X5974 132 10 171 203 369 643 664 AND2_X1 $T=28740 26200 1 0 $X=28625 $Y=24685
X5975 460 146 171 203 490 643 657 AND2_X1 $T=30450 26200 1 180 $X=29575 $Y=26085
X5976 136 10 171 203 266 634 659 AND2_X1 $T=30640 34600 0 180 $X=29765 $Y=33085
X5977 372 146 171 203 517 643 664 AND2_X1 $T=31020 26200 0 180 $X=30145 $Y=24685
X5978 462 146 171 203 376 643 657 AND2_X1 $T=32350 26200 0 0 $X=32235 $Y=26085
X5979 377 10 171 203 273 644 666 AND2_X1 $T=33490 3800 0 0 $X=33375 $Y=3685
X5980 154 10 171 203 382 647 659 AND2_X1 $T=34440 31800 0 0 $X=34325 $Y=31685
X5981 160 161 171 203 465 648 663 AND2_X1 $T=36530 17800 0 0 $X=36415 $Y=17685
X5982 131 10 171 203 386 645 658 AND2_X1 $T=36530 20600 0 0 $X=36415 $Y=20485
X5983 272 10 171 203 172 644 666 AND2_X1 $T=37100 3800 0 0 $X=36985 $Y=3685
X5984 467 161 171 203 560 648 663 AND2_X1 $T=38050 17800 0 0 $X=37935 $Y=17685
X5985 280 10 171 203 524 644 661 AND2_X1 $T=41280 3800 1 0 $X=41165 $Y=2285
X5986 472 10 171 203 398 639 655 AND2_X1 $T=43180 6600 0 0 $X=43065 $Y=6485
X5987 471 10 171 203 399 635 654 AND2_X1 $T=43180 12200 0 0 $X=43065 $Y=12085
X5988 400 10 171 203 401 648 660 AND2_X1 $T=43750 17800 1 0 $X=43635 $Y=16285
X5989 470 10 171 203 563 644 666 AND2_X1 $T=44320 3800 0 0 $X=44205 $Y=3685
X6285 230 203 621 422 308 69 171 641 652 NOR4_X1 $T=12970 37400 1 0 $X=12855 $Y=35885
X6286 331 203 620 438 439 101 171 642 664 NOR4_X1 $T=17150 23400 0 0 $X=17035 $Y=23285
X6287 255 203 513 351 450 256 171 648 663 NOR4_X1 $T=23230 17800 1 180 $X=22165 $Y=17685
X6288 153 203 461 363 275 385 171 637 655 NOR4_X1 $T=33870 9400 1 0 $X=33755 $Y=7885
X6289 163 203 164 379 156 160 171 642 658 NOR4_X1 $T=34060 23400 1 0 $X=33945 $Y=21885
X6290 375 203 371 380 277 622 171 639 666 NOR4_X1 $T=34250 6600 1 0 $X=34135 $Y=5085
X6291 495 203 403 185 392 391 171 637 653 NOR4_X1 $T=42230 9400 1 180 $X=41165 $Y=9285
X6292 497 203 396 394 476 383 171 635 653 NOR4_X1 $T=43560 12200 0 180 $X=42495 $Y=10685
X6326 170 518 363 380 203 171 377 644 666 FA_X1 $T=30450 3800 0 0 $X=30335 $Y=3685
X6327 518 150 461 371 203 171 272 639 655 FA_X1 $T=30830 6600 0 0 $X=30715 $Y=6485
X6328 561 170 275 277 203 171 280 639 666 FA_X1 $T=39380 6600 0 180 $X=36225 $Y=5085
X6329 468 561 497 495 203 171 470 639 655 FA_X1 $T=40140 6600 0 0 $X=40025 $Y=6485
X6330 186 402 394 185 203 171 471 635 654 FA_X1 $T=40140 12200 0 0 $X=40025 $Y=12085
X6331 402 468 396 403 203 171 472 637 655 FA_X1 $T=45080 9400 0 180 $X=41925 $Y=7885
X6332 389 186 174 476 203 171 400 636 660 FA_X1 $T=42040 15000 0 0 $X=41925 $Y=14885
X6333 503 2 171 203 498 548 2 221 649 661 ICV_27 $T=1000 1000 0 0 $X=885 $Y=885
X6334 425 2 171 203 287 210 4 34 645 663 ICV_27 $T=1000 20600 1 0 $X=885 $Y=19085
X6335 549 2 171 203 499 310 2 479 647 659 ICV_27 $T=1000 31800 0 0 $X=885 $Y=31685
X6336 575 3 171 203 31 576 3 49 651 668 ICV_27 $T=4230 48600 1 0 $X=4115 $Y=47085
X6337 231 3 171 203 82 511 4 118 650 662 ICV_27 $T=17530 43000 0 0 $X=17415 $Y=42885
X6338 580 3 171 203 92 251 3 120 651 668 ICV_27 $T=17910 48600 1 0 $X=17795 $Y=47085
X6339 250 3 171 203 105 253 3 113 650 665 ICV_27 $T=18290 43000 1 0 $X=18175 $Y=41485
X6340 260 2 171 203 264 584 3 461 639 655 ICV_27 $T=24370 6600 0 0 $X=24255 $Y=6485
X6341 583 3 171 203 128 585 3 148 651 668 ICV_27 $T=24370 48600 1 0 $X=24255 $Y=47085
X6342 263 3 171 203 142 368 2 267 635 653 ICV_27 $T=25890 12200 1 0 $X=25775 $Y=10685
X6343 539 4 171 203 133 269 3 276 650 662 ICV_27 $T=28550 43000 0 0 $X=28435 $Y=42885
X6344 538 4 171 203 370 157 3 463 636 660 ICV_27 $T=30450 15000 0 0 $X=30335 $Y=14885
X6345 586 3 171 203 380 273 2 521 649 661 ICV_27 $T=32160 1000 0 0 $X=32045 $Y=885
X6346 587 3 171 203 167 588 3 175 651 668 ICV_27 $T=35390 48600 1 0 $X=35275 $Y=47085
X6347 169 3 171 203 277 590 3 495 644 666 ICV_27 $T=37860 3800 0 0 $X=37745 $Y=3685
X6348 172 2 171 203 523 524 2 615 649 661 ICV_27 $T=38620 1000 0 0 $X=38505 $Y=885
X6349 591 3 171 203 394 607 3 392 636 654 ICV_27 $T=41850 15000 1 0 $X=41735 $Y=13485
X6350 282 4 171 203 197 608 3 194 642 658 ICV_27 $T=41850 23400 1 0 $X=41735 $Y=21885
X6351 406 4 171 203 191 597 3 200 640 657 ICV_27 $T=41850 29000 1 0 $X=41735 $Y=27485
X6352 522 4 171 203 193 603 3 196 638 656 ICV_27 $T=41850 40200 1 0 $X=41735 $Y=38685
X6368 295 171 203 500 637 655 INV_X1 $T=4230 9400 1 0 $X=4115 $Y=7885
X6369 208 171 203 9 637 653 INV_X1 $T=6130 9400 1 180 $X=5635 $Y=9285
X6370 207 171 203 25 650 665 INV_X1 $T=6890 43000 1 0 $X=6775 $Y=41485
X6371 300 171 203 216 650 665 INV_X1 $T=7270 43000 1 0 $X=7155 $Y=41485
X6372 418 171 203 26 637 653 INV_X1 $T=7460 9400 0 0 $X=7345 $Y=9285
X6373 303 171 203 414 638 665 INV_X1 $T=8030 40200 1 180 $X=7535 $Y=40085
X6374 38 171 203 213 637 655 INV_X1 $T=9740 9400 0 180 $X=9245 $Y=7885
X6375 311 171 203 526 638 665 INV_X1 $T=9550 40200 0 0 $X=9435 $Y=40085
X6376 309 171 203 307 637 655 INV_X1 $T=10120 9400 0 180 $X=9625 $Y=7885
X6377 36 171 203 423 636 654 INV_X1 $T=9740 15000 1 0 $X=9625 $Y=13485
X6378 423 171 203 47 637 653 INV_X1 $T=10120 9400 0 0 $X=10005 $Y=9285
X6379 527 171 203 324 642 664 INV_X1 $T=10500 23400 0 0 $X=10385 $Y=23285
X6380 612 171 203 50 642 658 INV_X1 $T=10690 23400 1 0 $X=10575 $Y=21885
X6381 226 171 203 426 637 655 INV_X1 $T=10880 9400 1 0 $X=10765 $Y=7885
X6382 483 171 203 481 641 656 INV_X1 $T=11450 37400 1 180 $X=10955 $Y=37285
X6383 313 171 203 70 643 657 INV_X1 $T=12210 26200 0 0 $X=12095 $Y=26085
X6384 434 171 203 504 643 664 INV_X1 $T=12590 26200 1 0 $X=12475 $Y=24685
X6385 430 171 203 61 638 665 INV_X1 $T=12590 40200 0 0 $X=12475 $Y=40085
X6386 613 171 203 59 635 653 INV_X1 $T=12970 12200 1 0 $X=12855 $Y=10685
X6387 435 171 203 77 635 654 INV_X1 $T=15820 12200 0 0 $X=15705 $Y=12085
X6388 330 171 203 243 638 656 INV_X1 $T=16010 40200 1 0 $X=15895 $Y=38685
X6389 337 171 203 236 645 658 INV_X1 $T=16770 20600 1 180 $X=16275 $Y=20485
X6390 437 171 203 89 635 654 INV_X1 $T=16960 12200 0 0 $X=16845 $Y=12085
X6391 256 171 203 239 635 653 INV_X1 $T=17530 12200 0 180 $X=17035 $Y=10685
X6392 442 171 203 341 643 657 INV_X1 $T=18670 26200 1 180 $X=18175 $Y=26085
X6393 553 171 203 86 636 660 INV_X1 $T=19810 15000 0 0 $X=19695 $Y=14885
X6394 245 171 203 233 640 657 INV_X1 $T=20570 29000 1 0 $X=20455 $Y=27485
X6395 554 171 203 99 641 652 INV_X1 $T=20570 37400 1 0 $X=20455 $Y=35885
X6396 447 171 203 98 643 657 INV_X1 $T=21330 26200 1 180 $X=20835 $Y=26085
X6397 448 171 203 119 641 652 INV_X1 $T=22470 37400 1 0 $X=22355 $Y=35885
X6398 558 171 203 348 636 660 INV_X1 $T=23230 15000 1 180 $X=22735 $Y=14885
X6399 110 171 203 488 642 658 INV_X1 $T=23420 23400 1 0 $X=23305 $Y=21885
X6400 254 171 203 361 645 663 INV_X1 $T=25890 20600 1 0 $X=25775 $Y=19085
X6401 458 171 203 130 634 652 INV_X1 $T=27600 34600 0 0 $X=27485 $Y=34485
X6402 366 171 203 365 648 660 INV_X1 $T=28170 17800 0 180 $X=27675 $Y=16285
X6403 265 171 203 124 645 658 INV_X1 $T=29120 20600 1 180 $X=28625 $Y=20485
X6404 456 171 203 459 647 659 INV_X1 $T=29120 31800 0 0 $X=29005 $Y=31685
X6405 279 171 203 204 648 660 INV_X1 $T=31780 17800 1 0 $X=31665 $Y=16285
X6406 374 171 203 146 643 664 INV_X1 $T=32920 26200 0 180 $X=32425 $Y=24685
X6407 279 171 203 161 648 663 INV_X1 $T=37670 17800 0 0 $X=37555 $Y=17685
X6408 392 171 203 174 636 654 INV_X1 $T=41470 15000 1 0 $X=41355 $Y=13485
X6409 413 9 501 294 171 203 639 655 AOI21_X1 $T=4800 6600 0 0 $X=4685 $Y=6485
X6410 481 225 211 42 171 203 638 656 AOI21_X1 $T=9360 40200 1 0 $X=9245 $Y=38685
X6411 227 526 617 42 171 203 638 656 AOI21_X1 $T=10880 40200 0 180 $X=10005 $Y=38685
X6412 228 50 429 65 171 203 642 664 AOI21_X1 $T=11640 23400 0 0 $X=11525 $Y=23285
X6413 225 322 621 54 171 203 638 656 AOI21_X1 $T=12400 40200 1 0 $X=12285 $Y=38685
X6414 504 57 482 65 171 203 642 658 AOI21_X1 $T=13730 23400 1 0 $X=13615 $Y=21885
X6415 232 59 508 234 171 203 637 653 AOI21_X1 $T=13920 9400 0 0 $X=13805 $Y=9285
X6416 57 60 620 329 171 203 642 664 AOI21_X1 $T=13920 23400 0 0 $X=13805 $Y=23285
X6417 322 58 483 56 171 203 641 652 AOI21_X1 $T=14680 37400 0 180 $X=13805 $Y=35885
X6418 60 69 434 327 171 203 643 664 AOI21_X1 $T=14870 26200 1 0 $X=14755 $Y=24685
X6419 320 70 71 327 171 203 643 657 AOI21_X1 $T=15820 26200 1 180 $X=14945 $Y=26085
X6420 248 89 345 344 171 203 637 655 AOI21_X1 $T=20000 9400 0 180 $X=19125 $Y=7885
X6421 256 93 484 485 171 203 635 653 AOI21_X1 $T=19620 12200 1 0 $X=19505 $Y=10685
X6422 248 89 242 484 171 203 637 653 AOI21_X1 $T=19810 9400 0 0 $X=19695 $Y=9285
X6423 109 101 110 556 171 203 642 658 AOI21_X1 $T=21140 23400 1 0 $X=21025 $Y=21885
X6424 114 109 513 258 171 203 645 658 AOI21_X1 $T=23040 20600 0 0 $X=22925 $Y=20485
X6425 488 114 514 112 171 203 645 658 AOI21_X1 $T=24560 20600 1 180 $X=23685 $Y=20485
X6426 358 117 346 355 171 203 647 659 AOI21_X1 $T=24750 31800 1 180 $X=23875 $Y=31685
X6427 126 124 618 112 171 203 642 658 AOI21_X1 $T=25510 23400 1 0 $X=25395 $Y=21885
X6428 174 389 393 493 171 203 636 660 AOI21_X1 $T=41280 15000 0 0 $X=41165 $Y=14885
X6429 213 19 298 212 171 203 639 655 OAI21_X1 $T=6890 6600 0 0 $X=6775 $Y=6485
X6430 304 26 417 212 171 203 639 655 OAI21_X1 $T=7650 6600 0 0 $X=7535 $Y=6485
X6431 304 26 19 307 171 203 637 655 OAI21_X1 $T=8030 9400 1 0 $X=7915 $Y=7885
X6432 426 47 316 307 171 203 637 655 OAI21_X1 $T=11260 9400 1 0 $X=11145 $Y=7885
X6433 426 47 38 241 171 203 637 653 OAI21_X1 $T=11260 9400 0 0 $X=11145 $Y=9285
X6434 321 61 509 322 171 203 638 656 OAI21_X1 $T=15060 40200 0 180 $X=14185 $Y=38685
X6435 242 76 332 238 171 203 637 655 OAI21_X1 $T=16010 9400 1 0 $X=15895 $Y=7885
X6436 336 77 340 238 171 203 639 655 OAI21_X1 $T=16960 6600 1 180 $X=16085 $Y=6485
X6437 249 86 343 93 171 203 635 654 OAI21_X1 $T=18860 12200 0 0 $X=18745 $Y=12085
X6438 364 98 446 109 171 203 642 664 OAI21_X1 $T=20760 23400 0 0 $X=20645 $Y=23285
X6439 252 99 555 346 171 203 634 659 OAI21_X1 $T=20760 34600 1 0 $X=20645 $Y=33085
X6440 252 99 486 97 171 203 634 652 OAI21_X1 $T=21710 34600 1 180 $X=20835 $Y=34485
X6441 116 119 619 358 171 203 634 659 OAI21_X1 $T=24180 34600 1 0 $X=24065 $Y=33085
X6442 367 130 456 117 171 203 647 659 OAI21_X1 $T=27030 31800 0 0 $X=26915 $Y=31685
X6443 270 156 374 161 171 203 642 664 OAI21_X1 $T=33680 23400 0 0 $X=33565 $Y=23285
X6444 389 174 493 161 171 203 648 660 OAI21_X1 $T=40520 17800 0 180 $X=39645 $Y=16285
X6445 171 374 115 2 171 203 642 664 CLKGATETST_X8 $T=27600 23400 0 0 $X=27485 $Y=23285
X6446 171 465 1 261 171 203 648 663 CLKGATETST_X8 $T=38810 17800 0 0 $X=38695 $Y=17685
X6512 171 500 285 5 203 639 655 XNOR2_X1 $T=3280 6600 1 180 $X=2025 $Y=6485
X6513 171 420 286 297 203 641 656 XNOR2_X1 $T=8030 37400 1 180 $X=6775 $Y=37285
X6514 171 417 222 22 203 639 666 XNOR2_X1 $T=7270 6600 1 0 $X=7155 $Y=5085
X6515 171 69 436 71 203 640 667 XNOR2_X1 $T=15060 29000 0 0 $X=14945 $Y=28885
X6516 171 340 338 81 203 639 655 XNOR2_X1 $T=18100 6600 1 180 $X=16845 $Y=6485
X6517 171 441 440 84 203 642 658 XNOR2_X1 $T=18860 23400 0 180 $X=17605 $Y=21885
X6518 171 346 352 486 203 634 659 XNOR2_X1 $T=22470 34600 1 0 $X=22355 $Y=33085
X6519 171 614 359 454 203 648 660 XNOR2_X1 $T=24560 17800 1 0 $X=24445 $Y=16285
X6520 171 463 467 492 203 648 660 XNOR2_X1 $T=39000 17800 0 180 $X=37745 $Y=16285
X6531 413 203 9 294 171 639 655 NOR2_X1 $T=6130 6600 1 180 $X=5445 $Y=6485
X6532 212 203 294 502 171 637 655 NOR2_X1 $T=6510 9400 0 180 $X=5825 $Y=7885
X6533 224 203 206 295 171 635 653 NOR2_X1 $T=6510 12200 0 180 $X=5825 $Y=10685
X6534 414 203 416 546 171 638 665 NOR2_X1 $T=7080 40200 1 180 $X=6395 $Y=40085
X6535 302 203 25 416 171 638 665 NOR2_X1 $T=7650 40200 1 180 $X=6965 $Y=40085
X6536 37 203 216 306 171 641 652 NOR2_X1 $T=8220 37400 1 0 $X=8105 $Y=35885
X6537 308 203 306 420 171 641 652 NOR2_X1 $T=8790 37400 1 0 $X=8675 $Y=35885
X6538 213 203 309 22 171 639 655 NOR2_X1 $T=9550 6600 1 180 $X=8865 $Y=6485
X6539 226 203 423 309 171 637 653 NOR2_X1 $T=9550 9400 0 0 $X=9435 $Y=9285
X6540 303 203 306 422 171 641 652 NOR2_X1 $T=10120 37400 0 180 $X=9435 $Y=35885
X6541 227 203 526 42 171 638 665 NOR2_X1 $T=10500 40200 0 0 $X=10385 $Y=40085
X6542 228 203 50 65 171 642 658 NOR2_X1 $T=11640 23400 1 0 $X=11525 $Y=21885
X6543 321 203 61 56 171 638 656 NOR2_X1 $T=13160 40200 1 0 $X=13045 $Y=38685
X6544 236 203 68 323 171 645 658 NOR2_X1 $T=14490 20600 1 180 $X=13805 $Y=20485
X6545 232 203 59 234 171 635 653 NOR2_X1 $T=14110 12200 1 0 $X=13995 $Y=10685
X6546 320 203 70 327 171 643 657 NOR2_X1 $T=14490 26200 0 0 $X=14375 $Y=26085
X6547 326 203 324 68 171 642 658 NOR2_X1 $T=16010 23400 0 180 $X=15325 $Y=21885
X6548 485 203 334 67 171 635 653 NOR2_X1 $T=17150 12200 0 180 $X=16465 $Y=10685
X6549 337 203 339 438 171 642 658 NOR2_X1 $T=17150 23400 1 0 $X=17035 $Y=21885
X6550 83 203 341 339 171 643 664 NOR2_X1 $T=17340 26200 1 0 $X=17225 $Y=24685
X6551 439 203 339 441 171 642 664 NOR2_X1 $T=18100 23400 0 0 $X=17985 $Y=23285
X6552 242 203 344 81 171 639 655 NOR2_X1 $T=19240 6600 1 180 $X=18555 $Y=6485
X6553 248 203 89 344 171 637 655 NOR2_X1 $T=18670 9400 1 0 $X=18555 $Y=7885
X6554 249 203 86 485 171 635 654 NOR2_X1 $T=19620 12200 0 0 $X=19505 $Y=12085
X6555 106 203 348 347 171 648 660 NOR2_X1 $T=21710 17800 1 0 $X=21595 $Y=16285
X6556 364 203 98 556 171 642 664 NOR2_X1 $T=22660 23400 1 180 $X=21975 $Y=23285
X6557 254 203 347 351 171 645 663 NOR2_X1 $T=22850 20600 1 0 $X=22735 $Y=19085
X6558 450 203 347 614 171 648 660 NOR2_X1 $T=23040 17800 1 0 $X=22925 $Y=16285
X6559 116 203 119 355 171 634 659 NOR2_X1 $T=23610 34600 1 0 $X=23495 $Y=33085
X6560 126 203 124 112 171 645 658 NOR2_X1 $T=25700 20600 0 0 $X=25585 $Y=20485
X6561 453 203 365 111 171 648 663 NOR2_X1 $T=26270 17800 0 0 $X=26155 $Y=17685
X6562 361 203 111 455 171 645 663 NOR2_X1 $T=26270 20600 1 0 $X=26155 $Y=19085
X6563 379 203 279 519 171 645 658 NOR2_X1 $T=34060 20600 1 180 $X=33375 $Y=20485
X6564 466 203 163 388 171 642 664 NOR2_X1 $T=37860 23400 1 180 $X=37175 $Y=23285
X6565 379 171 164 163 203 270 642 658 NAND3_X1 $T=34060 23400 0 180 $X=33185 $Y=21885
X6566 378 171 464 387 203 492 635 654 NAND3_X1 $T=38050 12200 1 180 $X=37175 $Y=12085
X6567 302 171 25 303 203 638 656 NAND2_X1 $T=7460 40200 1 0 $X=7345 $Y=38685
X6568 304 171 26 212 203 637 653 NAND2_X1 $T=8410 9400 1 180 $X=7725 $Y=9285
X6569 227 171 526 225 203 638 665 NAND2_X1 $T=10500 40200 1 180 $X=9815 $Y=40085
X6570 228 171 50 57 203 642 658 NAND2_X1 $T=12210 23400 1 0 $X=12095 $Y=21885
X6571 321 171 61 322 203 638 656 NAND2_X1 $T=13730 40200 1 0 $X=13615 $Y=38685
X6572 320 171 70 60 203 643 664 NAND2_X1 $T=14300 26200 1 0 $X=14185 $Y=24685
X6573 336 171 77 238 203 639 655 NAND2_X1 $T=15630 6600 0 0 $X=15515 $Y=6485
X6574 326 171 324 337 203 642 658 NAND2_X1 $T=16580 23400 1 0 $X=16465 $Y=21885
X6575 555 171 97 244 203 634 652 NAND2_X1 $T=20380 34600 1 180 $X=19695 $Y=34485
X6576 249 171 86 93 203 635 654 NAND2_X1 $T=20760 12200 1 180 $X=20075 $Y=12085
X6577 252 171 99 97 203 634 652 NAND2_X1 $T=20950 34600 1 180 $X=20265 $Y=34485
X6578 364 171 98 109 203 642 664 NAND2_X1 $T=21520 23400 0 0 $X=21405 $Y=23285
X6579 116 171 119 358 203 634 652 NAND2_X1 $T=23990 34600 0 0 $X=23875 $Y=34485
X6580 453 171 365 254 203 648 660 NAND2_X1 $T=26270 17800 0 180 $X=25585 $Y=16285
X6581 126 171 124 114 203 642 658 NAND2_X1 $T=26270 23400 1 0 $X=26155 $Y=21885
X6582 367 171 130 117 203 634 659 NAND2_X1 $T=28170 34600 0 180 $X=27485 $Y=33085
X6583 153 171 375 271 203 637 655 NAND2_X1 $T=32540 9400 1 0 $X=32425 $Y=7885
X6584 391 171 622 464 203 637 653 NAND2_X1 $T=36530 9400 0 0 $X=36415 $Y=9285
X6585 383 171 385 387 203 635 653 NAND2_X1 $T=36720 12200 1 0 $X=36605 $Y=10685
X6586 464 171 387 278 203 635 654 NAND2_X1 $T=37290 12200 1 180 $X=36605 $Y=12085
X6587 413 9 293 171 502 5 203 637 655 AOI211_X1 $T=4990 9400 1 0 $X=4875 $Y=7885
X6588 271 150 278 171 279 274 203 635 654 AOI211_X1 $T=33680 12200 0 0 $X=33565 $Y=12085
X6589 466 163 374 171 388 520 203 642 664 AOI211_X1 $T=37290 23400 1 180 $X=36225 $Y=23285
X6590 460 379 151 171 203 491 643 657 HA_X1 $T=30450 26200 0 0 $X=30335 $Y=26085
X6591 462 491 152 171 203 384 640 657 HA_X1 $T=33490 29000 0 180 $X=31475 $Y=27485
X6592 372 384 164 171 203 466 643 664 HA_X1 $T=35960 26200 1 0 $X=35845 $Y=24685
X6593 202 171 203 1 637 653 CLKBUF_X3 $T=1000 9400 0 0 $X=885 $Y=9285
X6594 223 171 203 4 647 659 CLKBUF_X3 $T=24750 31800 0 0 $X=24635 $Y=31685
X6595 261 171 203 3 643 657 CLKBUF_X3 $T=26270 26200 0 0 $X=26155 $Y=26085
X6596 381 171 203 245 648 660 CLKBUF_X3 $T=35200 17800 1 0 $X=35085 $Y=16285
X6634 234 76 171 203 334 635 653 OR2_X1 $T=15820 12200 1 0 $X=15705 $Y=10685
X6635 375 153 171 203 150 637 655 OR2_X1 $T=33870 9400 0 180 $X=32995 $Y=7885
X6636 152 151 171 203 156 643 657 OR2_X1 $T=33680 26200 0 0 $X=33565 $Y=26085
X6637 245 154 171 203 559 647 659 OR2_X1 $T=33680 31800 0 0 $X=33565 $Y=31685
X6654 1 407 204 171 203 15 644 666 DFFR_X1 $T=1000 3800 0 0 $X=885 $Y=3685
X6655 1 285 204 171 203 11 639 666 DFFR_X1 $T=1000 6600 1 0 $X=885 $Y=5085
X6656 1 286 204 171 203 12 641 652 DFFR_X1 $T=1000 37400 1 0 $X=885 $Y=35885
X6657 1 408 204 171 203 29 641 656 DFFR_X1 $T=1000 37400 0 0 $X=885 $Y=37285
X6658 1 222 204 171 203 40 644 666 DFFR_X1 $T=7460 3800 0 0 $X=7345 $Y=3685
X6659 1 424 204 171 203 55 639 655 DFFR_X1 $T=9550 6600 0 0 $X=9435 $Y=6485
X6660 1 427 204 171 203 45 648 663 DFFR_X1 $T=10690 17800 0 0 $X=10575 $Y=17685
X6661 1 428 204 171 203 75 644 666 DFFR_X1 $T=11260 3800 0 0 $X=11145 $Y=3685
X6662 51 53 204 171 203 328 634 652 DFFR_X1 $T=12210 34600 0 0 $X=12095 $Y=34485
X6663 51 317 204 171 203 52 640 657 DFFR_X1 $T=13540 29000 1 0 $X=13425 $Y=27485
X6664 1 325 204 171 203 104 636 654 DFFR_X1 $T=14680 15000 1 0 $X=14565 $Y=13485
X6665 51 436 204 171 203 32 647 659 DFFR_X1 $T=15630 31800 0 0 $X=15515 $Y=31685
X6666 1 338 204 171 203 95 639 666 DFFR_X1 $T=16390 6600 1 0 $X=16275 $Y=5085
X6667 51 333 204 171 203 72 641 652 DFFR_X1 $T=16770 37400 1 0 $X=16655 $Y=35885
X6668 1 440 204 171 203 74 645 658 DFFR_X1 $T=17530 20600 0 0 $X=17415 $Y=20485
X6669 51 445 204 171 203 90 647 659 DFFR_X1 $T=20190 31800 0 0 $X=20075 $Y=31685
X6670 51 444 204 171 203 43 643 657 DFFR_X1 $T=21330 26200 0 0 $X=21215 $Y=26085
X6671 1 350 204 171 203 103 637 655 DFFR_X1 $T=22090 9400 1 0 $X=21975 $Y=7885
X6672 51 352 204 171 203 121 647 667 DFFR_X1 $T=22470 31800 1 0 $X=22355 $Y=30285
X6673 115 360 204 171 203 132 642 664 DFFR_X1 $T=23800 23400 0 0 $X=23685 $Y=23285
X6674 115 359 204 171 203 129 636 654 DFFR_X1 $T=24370 15000 1 0 $X=24255 $Y=13485
X6675 115 362 204 171 203 136 647 667 DFFR_X1 $T=26270 31800 1 0 $X=26155 $Y=30285
X6676 115 457 204 171 203 131 645 658 DFFR_X1 $T=29690 20600 0 0 $X=29575 $Y=20485
X6677 224 6 203 7 300 206 171 650 665 AOI22_X1 $T=5560 43000 1 0 $X=5445 $Y=41485
X6678 224 16 203 21 208 206 171 648 660 AOI22_X1 $T=5750 17800 1 0 $X=5635 $Y=16285
X6679 224 411 203 8 207 206 171 650 662 AOI22_X1 $T=5750 43000 0 0 $X=5635 $Y=42885
X6680 224 17 203 13 418 206 171 635 653 AOI22_X1 $T=7460 12200 0 180 $X=6395 $Y=10685
X6681 224 28 203 33 36 206 171 636 654 AOI22_X1 $T=8790 15000 1 0 $X=8675 $Y=13485
X6682 224 480 203 20 527 206 171 640 657 AOI22_X1 $T=9930 29000 0 180 $X=8865 $Y=27485
X6683 224 34 203 30 612 206 171 642 658 AOI22_X1 $T=9360 23400 1 0 $X=9245 $Y=21885
X6684 224 35 203 31 311 206 171 650 662 AOI22_X1 $T=10310 43000 1 180 $X=9245 $Y=42885
X6685 224 14 203 18 313 206 171 643 664 AOI22_X1 $T=9740 26200 1 0 $X=9625 $Y=24685
X6686 224 23 203 27 613 206 171 635 653 AOI22_X1 $T=12020 12200 1 0 $X=11905 $Y=10685
X6687 224 46 203 49 430 206 171 650 662 AOI22_X1 $T=12400 43000 0 0 $X=12285 $Y=42885
X6688 224 41 203 44 435 206 171 635 654 AOI22_X1 $T=14490 12200 0 0 $X=14375 $Y=12085
X6689 224 66 203 62 330 206 171 638 656 AOI22_X1 $T=16010 40200 0 180 $X=14945 $Y=38685
X6690 224 73 203 64 437 206 171 636 660 AOI22_X1 $T=16010 15000 0 0 $X=15895 $Y=14885
X6691 224 85 203 87 442 206 171 640 657 AOI22_X1 $T=17340 29000 1 0 $X=17225 $Y=27485
X6692 248 89 203 86 246 249 171 635 653 AOI22_X1 $T=18670 12200 1 0 $X=18555 $Y=10685
X6693 224 100 203 96 553 206 171 648 660 AOI22_X1 $T=19430 17800 1 0 $X=19315 $Y=16285
X6694 224 80 203 82 554 206 171 641 656 AOI22_X1 $T=19430 37400 0 0 $X=19315 $Y=37285
X6695 224 108 203 113 447 206 171 640 657 AOI22_X1 $T=22470 29000 0 180 $X=21405 $Y=27485
X6696 224 102 203 105 448 206 171 641 652 AOI22_X1 $T=22470 37400 0 180 $X=21405 $Y=35885
X6697 224 356 203 107 558 206 171 636 654 AOI22_X1 $T=24370 15000 0 180 $X=23305 $Y=13485
X6698 224 145 203 141 458 206 171 634 652 AOI22_X1 $T=26650 34600 0 0 $X=26535 $Y=34485
X6699 224 140 203 142 265 206 171 645 663 AOI22_X1 $T=27980 20600 1 0 $X=27865 $Y=19085
X6700 224 370 203 143 366 206 171 636 660 AOI22_X1 $T=30450 15000 1 180 $X=29385 $Y=14885
X6706 203 501 407 298 171 639 655 XOR2_X1 $T=1000 6600 0 0 $X=885 $Y=6485
X6707 203 211 408 546 171 638 656 XOR2_X1 $T=5180 40200 0 180 $X=3925 $Y=38685
X6708 203 483 53 617 171 641 652 XOR2_X1 $T=10120 37400 1 0 $X=10005 $Y=35885
X6709 203 434 317 429 171 643 664 XOR2_X1 $T=12590 26200 0 180 $X=11335 $Y=24685
X6710 203 241 424 316 171 637 653 XOR2_X1 $T=12020 9400 0 0 $X=11905 $Y=9285
X6711 203 482 427 323 171 645 658 XOR2_X1 $T=13920 20600 1 180 $X=12665 $Y=20485
X6712 203 508 428 332 171 637 655 XOR2_X1 $T=13540 9400 1 0 $X=13425 $Y=7885
X6713 203 58 333 509 171 641 656 XOR2_X1 $T=15630 37400 0 0 $X=15515 $Y=37285
X6714 203 256 325 343 171 635 654 XOR2_X1 $T=17340 12200 0 0 $X=17225 $Y=12085
X6715 203 244 445 443 171 634 659 XOR2_X1 $T=17910 34600 1 0 $X=17795 $Y=33085
X6716 203 243 443 78 171 634 652 XOR2_X1 $T=19810 34600 1 180 $X=18555 $Y=34485
X6717 203 101 444 446 171 642 664 XOR2_X1 $T=19620 23400 0 0 $X=19505 $Y=23285
X6718 203 484 350 345 171 637 653 XOR2_X1 $T=20570 9400 0 0 $X=20455 $Y=9285
X6719 203 110 360 618 171 642 658 XOR2_X1 $T=24370 23400 1 0 $X=24255 $Y=21885
X6720 203 117 362 619 171 647 659 XOR2_X1 $T=25890 31800 0 0 $X=25775 $Y=31685
X6721 203 514 457 455 171 645 663 XOR2_X1 $T=26840 20600 1 0 $X=26725 $Y=19085
X6728 292 171 203 412 644 661 CLKBUF_X1 $T=4990 3800 1 0 $X=4875 $Y=2285
X6729 296 171 203 290 634 659 CLKBUF_X1 $T=4990 34600 1 0 $X=4875 $Y=33085
X6730 415 171 203 220 644 666 CLKBUF_X1 $T=6130 3800 0 0 $X=6015 $Y=3685
X6731 412 171 203 503 644 661 CLKBUF_X1 $T=6890 3800 0 180 $X=6205 $Y=2285
X6732 290 171 203 299 634 659 CLKBUF_X1 $T=7650 34600 0 180 $X=6965 $Y=33085
X6733 220 171 203 548 644 661 CLKBUF_X1 $T=8030 3800 0 180 $X=7345 $Y=2285
X6734 550 171 203 549 647 659 CLKBUF_X1 $T=8030 31800 1 180 $X=7345 $Y=31685
X6735 547 171 203 550 634 659 CLKBUF_X1 $T=8220 34600 0 180 $X=7535 $Y=33085
X6736 312 171 203 229 645 663 CLKBUF_X1 $T=9550 20600 1 0 $X=9435 $Y=19085
X6737 229 171 203 425 645 663 CLKBUF_X1 $T=11450 20600 0 180 $X=10765 $Y=19085
X6738 48 171 203 552 645 658 CLKBUF_X1 $T=11640 20600 0 0 $X=11525 $Y=20485
X6739 552 171 203 318 645 658 CLKBUF_X1 $T=12780 20600 1 180 $X=12095 $Y=20485
X6740 431 171 203 319 644 661 CLKBUF_X1 $T=12780 3800 1 0 $X=12665 $Y=2285
X6741 319 171 203 505 644 661 CLKBUF_X1 $T=14680 3800 0 180 $X=13995 $Y=2285
X6742 237 171 203 510 644 661 CLKBUF_X1 $T=15060 3800 1 0 $X=14945 $Y=2285
X6743 616 171 203 237 644 666 CLKBUF_X1 $T=16770 3800 1 180 $X=16085 $Y=3685
X6744 1 171 203 51 640 657 CLKBUF_X1 $T=20000 29000 1 0 $X=19885 $Y=27485
X6745 449 171 203 349 644 666 CLKBUF_X1 $T=22280 3800 0 0 $X=22165 $Y=3685
X6746 349 171 203 557 644 666 CLKBUF_X1 $T=23420 3800 1 180 $X=22735 $Y=3685
X6747 357 171 203 487 637 653 CLKBUF_X1 $T=23040 9400 0 0 $X=22925 $Y=9285
X6748 487 171 203 260 635 653 CLKBUF_X1 $T=24560 12200 1 0 $X=24445 $Y=10685
X6749 259 171 203 451 639 666 CLKBUF_X1 $T=24750 6600 1 0 $X=24635 $Y=5085
X6750 451 171 203 452 639 666 CLKBUF_X1 $T=25890 6600 0 180 $X=25205 $Y=5085
X6751 1 171 203 115 636 660 CLKBUF_X1 $T=25700 15000 0 0 $X=25585 $Y=14885
X6752 211 414 171 297 25 302 203 638 656 OAI22_X1 $T=6510 40200 1 0 $X=6395 $Y=38685
X6753 482 236 171 84 324 326 203 642 658 OAI22_X1 $T=14490 23400 1 0 $X=14375 $Y=21885
X6754 244 335 171 58 243 78 203 634 652 OAI22_X1 $T=16960 34600 1 180 $X=15895 $Y=34485
X6755 238 234 171 63 334 246 203 637 653 OAI22_X1 $T=16390 9400 0 0 $X=16275 $Y=9285
X6756 336 77 171 76 89 248 203 637 655 OAI22_X1 $T=16770 9400 1 0 $X=16655 $Y=7885
X6757 514 361 171 454 365 453 203 648 663 OAI22_X1 $T=26270 17800 1 180 $X=25205 $Y=17685
X6758 306 416 42 171 203 54 641 656 OR3_X1 $T=10120 37400 0 0 $X=10005 $Y=37285
X6759 339 68 65 171 203 329 642 664 OR3_X1 $T=15630 23400 1 180 $X=14565 $Y=23285
X6760 347 111 112 171 203 258 645 663 OR3_X1 $T=23420 20600 1 0 $X=23305 $Y=19085
X6761 213 203 19 294 171 293 637 653 NOR3_X1 $T=6890 9400 1 180 $X=6015 $Y=9285
X6762 58 203 56 54 171 230 641 656 NOR3_X1 $T=13920 37400 1 180 $X=13045 $Y=37285
X6763 69 203 327 329 171 331 643 664 NOR3_X1 $T=15630 26200 1 0 $X=15515 $Y=24685
X6764 101 203 556 258 171 255 645 658 NOR3_X1 $T=21330 20600 0 0 $X=21215 $Y=20485
.ENDS
***************************************
