/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 23:24:37 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1502180417 */

module datapath(p_0, Accumulator, Accumulator1);
   input [23:0]p_0;
   input [23:0]Accumulator;
   output [23:0]Accumulator1;

   HA_X1 i_0 (.A(p_0[0]), .B(Accumulator[0]), .CO(n_0), .S(Accumulator1[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(Accumulator[1]), .CI(n_0), .CO(n_1), .S(
      Accumulator1[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(Accumulator[2]), .CI(n_1), .CO(n_2), .S(
      Accumulator1[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(Accumulator[3]), .CI(n_2), .CO(n_3), .S(
      Accumulator1[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(Accumulator[4]), .CI(n_3), .CO(n_4), .S(
      Accumulator1[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(Accumulator[5]), .CI(n_4), .CO(n_5), .S(
      Accumulator1[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(Accumulator[6]), .CI(n_5), .CO(n_6), .S(
      Accumulator1[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(Accumulator[7]), .CI(n_6), .CO(n_7), .S(
      Accumulator1[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(Accumulator[8]), .CI(n_7), .CO(n_8), .S(
      Accumulator1[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(Accumulator[9]), .CI(n_8), .CO(n_9), .S(
      Accumulator1[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(Accumulator[10]), .CI(n_9), .CO(n_10), .S(
      Accumulator1[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(Accumulator[11]), .CI(n_10), .CO(n_11), .S(
      Accumulator1[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(Accumulator[12]), .CI(n_11), .CO(n_12), .S(
      Accumulator1[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(Accumulator[13]), .CI(n_12), .CO(n_13), .S(
      Accumulator1[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(Accumulator[14]), .CI(n_13), .CO(n_14), .S(
      Accumulator1[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(Accumulator[15]), .CI(n_14), .CO(n_15), .S(
      Accumulator1[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(Accumulator[16]), .CI(n_15), .CO(n_16), .S(
      Accumulator1[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(Accumulator[17]), .CI(n_16), .CO(n_17), .S(
      Accumulator1[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(Accumulator[18]), .CI(n_17), .CO(n_18), .S(
      Accumulator1[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(Accumulator[19]), .CI(n_18), .CO(n_19), .S(
      Accumulator1[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(Accumulator[20]), .CI(n_19), .CO(n_20), .S(
      Accumulator1[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(Accumulator[21]), .CI(n_20), .CO(n_21), .S(
      Accumulator1[21]));
   FA_X1 i_22 (.A(p_0[22]), .B(Accumulator[22]), .CI(n_21), .CO(n_22), .S(
      Accumulator1[22]));
   XOR2_X1 i_23 (.A(p_0[23]), .B(n_22), .Z(Accumulator1[23]));
endmodule

module unsigned_seq_multiplier(clk, rst, start_s, a, b, c);
   input clk;
   input rst;
   input start_s;
   input [23:0]a;
   input [23:0]b;
   output [47:0]c;

   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire [23:0]A_r;
   wire n_0_1;
   wire n_0_0;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_1_2;
   wire n_0_49;
   wire n_0_1_3;
   wire n_0_50;
   wire n_0_1_4;
   wire n_0_51;
   wire n_0_1_5;
   wire n_0_52;
   wire n_0_1_6;
   wire n_0_53;
   wire n_0_1_7;
   wire n_0_54;
   wire n_0_1_8;
   wire n_0_55;
   wire n_0_1_9;
   wire n_0_56;
   wire n_0_1_10;
   wire n_0_57;
   wire n_0_1_11;
   wire n_0_58;
   wire n_0_1_12;
   wire n_0_59;
   wire n_0_1_13;
   wire n_0_60;
   wire n_0_1_14;
   wire n_0_61;
   wire n_0_1_15;
   wire n_0_62;
   wire n_0_1_16;
   wire n_0_63;
   wire n_0_1_17;
   wire n_0_64;
   wire n_0_1_18;
   wire n_0_65;
   wire n_0_1_19;
   wire n_0_66;
   wire n_0_1_20;
   wire n_0_67;
   wire n_0_1_21;
   wire n_0_68;
   wire n_0_1_22;
   wire n_0_69;
   wire n_0_1_23;
   wire n_0_70;
   wire n_0_1_24;
   wire n_0_71;
   wire n_0_1_25;
   wire n_0_96;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_1_26;

   assign c[47] = 1'b0;

   DFFR_X1 \Accumulator_reg[22]  (.D(n_0_95), .RN(n_0_1), .CK(clk), .Q(c[46]), 
      .QN());
   DFFR_X1 \Accumulator_reg[21]  (.D(n_0_94), .RN(n_0_1), .CK(clk), .Q(c[45]), 
      .QN());
   DFFR_X1 \Accumulator_reg[20]  (.D(n_0_93), .RN(n_0_1), .CK(clk), .Q(c[44]), 
      .QN());
   DFFR_X1 \Accumulator_reg[19]  (.D(n_0_92), .RN(n_0_1), .CK(clk), .Q(c[43]), 
      .QN());
   DFFR_X1 \Accumulator_reg[18]  (.D(n_0_91), .RN(n_0_1), .CK(clk), .Q(c[42]), 
      .QN());
   DFFR_X1 \Accumulator_reg[17]  (.D(n_0_90), .RN(n_0_1), .CK(clk), .Q(c[41]), 
      .QN());
   DFFR_X1 \Accumulator_reg[16]  (.D(n_0_89), .RN(n_0_1), .CK(clk), .Q(c[40]), 
      .QN());
   DFFR_X1 \Accumulator_reg[15]  (.D(n_0_88), .RN(n_0_1), .CK(clk), .Q(c[39]), 
      .QN());
   DFFR_X1 \Accumulator_reg[14]  (.D(n_0_87), .RN(n_0_1), .CK(clk), .Q(c[38]), 
      .QN());
   DFFR_X1 \Accumulator_reg[13]  (.D(n_0_86), .RN(n_0_1), .CK(clk), .Q(c[37]), 
      .QN());
   DFFR_X1 \Accumulator_reg[12]  (.D(n_0_85), .RN(n_0_1), .CK(clk), .Q(c[36]), 
      .QN());
   DFFR_X1 \Accumulator_reg[11]  (.D(n_0_84), .RN(n_0_1), .CK(clk), .Q(c[35]), 
      .QN());
   DFFR_X1 \Accumulator_reg[10]  (.D(n_0_83), .RN(n_0_1), .CK(clk), .Q(c[34]), 
      .QN());
   DFFR_X1 \Accumulator_reg[9]  (.D(n_0_82), .RN(n_0_1), .CK(clk), .Q(c[33]), 
      .QN());
   DFFR_X1 \Accumulator_reg[8]  (.D(n_0_81), .RN(n_0_1), .CK(clk), .Q(c[32]), 
      .QN());
   DFFR_X1 \Accumulator_reg[7]  (.D(n_0_80), .RN(n_0_1), .CK(clk), .Q(c[31]), 
      .QN());
   DFFR_X1 \Accumulator_reg[6]  (.D(n_0_79), .RN(n_0_1), .CK(clk), .Q(c[30]), 
      .QN());
   DFFR_X1 \Accumulator_reg[5]  (.D(n_0_78), .RN(n_0_1), .CK(clk), .Q(c[29]), 
      .QN());
   DFFR_X1 \Accumulator_reg[4]  (.D(n_0_77), .RN(n_0_1), .CK(clk), .Q(c[28]), 
      .QN());
   DFFR_X1 \Accumulator_reg[3]  (.D(n_0_76), .RN(n_0_1), .CK(clk), .Q(c[27]), 
      .QN());
   DFFR_X1 \Accumulator_reg[2]  (.D(n_0_75), .RN(n_0_1), .CK(clk), .Q(c[26]), 
      .QN());
   DFFR_X1 \Accumulator_reg[1]  (.D(n_0_74), .RN(n_0_1), .CK(clk), .Q(c[25]), 
      .QN());
   DFFR_X1 \Accumulator_reg[0]  (.D(n_0_73), .RN(n_0_1), .CK(clk), .Q(c[24]), 
      .QN());
   datapath i_0_4 (.p_0({n_0_96, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, 
      n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, 
      n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49}), 
      .Accumulator({uc_0, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, 
      n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, 
      n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26}), .Accumulator1({
      n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, 
      n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, 
      n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72}));
   DFF_X1 \B_r_reg[23]  (.D(n_0_72), .CK(n_0_0), .Q(c[23]), .QN());
   DFF_X1 \B_r_reg[22]  (.D(n_0_119), .CK(n_0_0), .Q(c[22]), .QN());
   DFF_X1 \B_r_reg[21]  (.D(n_0_118), .CK(n_0_0), .Q(c[21]), .QN());
   DFF_X1 \B_r_reg[20]  (.D(n_0_117), .CK(n_0_0), .Q(c[20]), .QN());
   DFF_X1 \B_r_reg[19]  (.D(n_0_116), .CK(n_0_0), .Q(c[19]), .QN());
   DFF_X1 \B_r_reg[18]  (.D(n_0_115), .CK(n_0_0), .Q(c[18]), .QN());
   DFF_X1 \B_r_reg[17]  (.D(n_0_114), .CK(n_0_0), .Q(c[17]), .QN());
   DFF_X1 \B_r_reg[16]  (.D(n_0_113), .CK(n_0_0), .Q(c[16]), .QN());
   DFF_X1 \B_r_reg[15]  (.D(n_0_112), .CK(n_0_0), .Q(c[15]), .QN());
   DFF_X1 \B_r_reg[14]  (.D(n_0_111), .CK(n_0_0), .Q(c[14]), .QN());
   DFF_X1 \B_r_reg[13]  (.D(n_0_110), .CK(n_0_0), .Q(c[13]), .QN());
   DFF_X1 \B_r_reg[12]  (.D(n_0_109), .CK(n_0_0), .Q(c[12]), .QN());
   DFF_X1 \B_r_reg[11]  (.D(n_0_108), .CK(n_0_0), .Q(c[11]), .QN());
   DFF_X1 \B_r_reg[10]  (.D(n_0_107), .CK(n_0_0), .Q(c[10]), .QN());
   DFF_X1 \B_r_reg[9]  (.D(n_0_106), .CK(n_0_0), .Q(c[9]), .QN());
   DFF_X1 \B_r_reg[8]  (.D(n_0_105), .CK(n_0_0), .Q(c[8]), .QN());
   DFF_X1 \B_r_reg[7]  (.D(n_0_104), .CK(n_0_0), .Q(c[7]), .QN());
   DFF_X1 \B_r_reg[6]  (.D(n_0_103), .CK(n_0_0), .Q(c[6]), .QN());
   DFF_X1 \B_r_reg[5]  (.D(n_0_102), .CK(n_0_0), .Q(c[5]), .QN());
   DFF_X1 \B_r_reg[4]  (.D(n_0_101), .CK(n_0_0), .Q(c[4]), .QN());
   DFF_X1 \B_r_reg[3]  (.D(n_0_100), .CK(n_0_0), .Q(c[3]), .QN());
   DFF_X1 \B_r_reg[2]  (.D(n_0_99), .CK(n_0_0), .Q(c[2]), .QN());
   DFF_X1 \B_r_reg[1]  (.D(n_0_98), .CK(n_0_0), .Q(c[1]), .QN());
   DFF_X1 \B_r_reg[0]  (.D(n_0_97), .CK(n_0_0), .Q(c[0]), .QN());
   DFF_X1 \A_r_reg[23]  (.D(n_0_25), .CK(n_0_0), .Q(A_r[23]), .QN());
   DFF_X1 \A_r_reg[22]  (.D(n_0_24), .CK(n_0_0), .Q(A_r[22]), .QN());
   DFF_X1 \A_r_reg[21]  (.D(n_0_23), .CK(n_0_0), .Q(A_r[21]), .QN());
   DFF_X1 \A_r_reg[20]  (.D(n_0_22), .CK(n_0_0), .Q(A_r[20]), .QN());
   DFF_X1 \A_r_reg[19]  (.D(n_0_21), .CK(n_0_0), .Q(A_r[19]), .QN());
   DFF_X1 \A_r_reg[18]  (.D(n_0_20), .CK(n_0_0), .Q(A_r[18]), .QN());
   DFF_X1 \A_r_reg[17]  (.D(n_0_19), .CK(n_0_0), .Q(A_r[17]), .QN());
   DFF_X1 \A_r_reg[16]  (.D(n_0_18), .CK(n_0_0), .Q(A_r[16]), .QN());
   DFF_X1 \A_r_reg[15]  (.D(n_0_17), .CK(n_0_0), .Q(A_r[15]), .QN());
   DFF_X1 \A_r_reg[14]  (.D(n_0_16), .CK(n_0_0), .Q(A_r[14]), .QN());
   DFF_X1 \A_r_reg[13]  (.D(n_0_15), .CK(n_0_0), .Q(A_r[13]), .QN());
   DFF_X1 \A_r_reg[12]  (.D(n_0_14), .CK(n_0_0), .Q(A_r[12]), .QN());
   DFF_X1 \A_r_reg[11]  (.D(n_0_13), .CK(n_0_0), .Q(A_r[11]), .QN());
   DFF_X1 \A_r_reg[10]  (.D(n_0_12), .CK(n_0_0), .Q(A_r[10]), .QN());
   DFF_X1 \A_r_reg[9]  (.D(n_0_11), .CK(n_0_0), .Q(A_r[9]), .QN());
   DFF_X1 \A_r_reg[8]  (.D(n_0_10), .CK(n_0_0), .Q(A_r[8]), .QN());
   DFF_X1 \A_r_reg[7]  (.D(n_0_9), .CK(n_0_0), .Q(A_r[7]), .QN());
   DFF_X1 \A_r_reg[6]  (.D(n_0_8), .CK(n_0_0), .Q(A_r[6]), .QN());
   DFF_X1 \A_r_reg[5]  (.D(n_0_7), .CK(n_0_0), .Q(A_r[5]), .QN());
   DFF_X1 \A_r_reg[4]  (.D(n_0_6), .CK(n_0_0), .Q(A_r[4]), .QN());
   DFF_X1 \A_r_reg[3]  (.D(n_0_5), .CK(n_0_0), .Q(A_r[3]), .QN());
   DFF_X1 \A_r_reg[2]  (.D(n_0_4), .CK(n_0_0), .Q(A_r[2]), .QN());
   DFF_X1 \A_r_reg[1]  (.D(n_0_3), .CK(n_0_0), .Q(A_r[1]), .QN());
   DFF_X1 \A_r_reg[0]  (.D(n_0_2), .CK(n_0_0), .Q(A_r[0]), .QN());
   INV_X1 i_0_0_0 (.A(rst), .ZN(n_0_1));
   CLKGATETST_X1 clk_gate_B_r_reg (.CK(clk), .E(n_0_1), .SE(1'b0), .GCK(n_0_0));
   MUX2_X1 i_0_1_0 (.A(c[1]), .B(b[1]), .S(start_s), .Z(n_0_97));
   MUX2_X1 i_0_1_1 (.A(c[2]), .B(b[2]), .S(start_s), .Z(n_0_98));
   MUX2_X1 i_0_1_2 (.A(c[3]), .B(b[3]), .S(start_s), .Z(n_0_99));
   MUX2_X1 i_0_1_3 (.A(c[4]), .B(b[4]), .S(start_s), .Z(n_0_100));
   MUX2_X1 i_0_1_4 (.A(c[5]), .B(b[5]), .S(start_s), .Z(n_0_101));
   MUX2_X1 i_0_1_5 (.A(c[6]), .B(b[6]), .S(start_s), .Z(n_0_102));
   MUX2_X1 i_0_1_6 (.A(c[7]), .B(b[7]), .S(start_s), .Z(n_0_103));
   MUX2_X1 i_0_1_7 (.A(c[8]), .B(b[8]), .S(start_s), .Z(n_0_104));
   MUX2_X1 i_0_1_8 (.A(c[9]), .B(b[9]), .S(start_s), .Z(n_0_105));
   MUX2_X1 i_0_1_9 (.A(c[10]), .B(b[10]), .S(start_s), .Z(n_0_106));
   MUX2_X1 i_0_1_10 (.A(c[11]), .B(b[11]), .S(start_s), .Z(n_0_107));
   MUX2_X1 i_0_1_11 (.A(c[12]), .B(b[12]), .S(start_s), .Z(n_0_108));
   MUX2_X1 i_0_1_12 (.A(c[13]), .B(b[13]), .S(start_s), .Z(n_0_109));
   MUX2_X1 i_0_1_13 (.A(c[14]), .B(b[14]), .S(start_s), .Z(n_0_110));
   MUX2_X1 i_0_1_14 (.A(c[15]), .B(b[15]), .S(start_s), .Z(n_0_111));
   MUX2_X1 i_0_1_15 (.A(c[16]), .B(b[16]), .S(start_s), .Z(n_0_112));
   MUX2_X1 i_0_1_16 (.A(c[17]), .B(b[17]), .S(start_s), .Z(n_0_113));
   MUX2_X1 i_0_1_17 (.A(c[18]), .B(b[18]), .S(start_s), .Z(n_0_114));
   MUX2_X1 i_0_1_18 (.A(c[19]), .B(b[19]), .S(start_s), .Z(n_0_115));
   MUX2_X1 i_0_1_19 (.A(c[20]), .B(b[20]), .S(start_s), .Z(n_0_116));
   MUX2_X1 i_0_1_20 (.A(c[21]), .B(b[21]), .S(start_s), .Z(n_0_117));
   MUX2_X1 i_0_1_21 (.A(c[22]), .B(b[22]), .S(start_s), .Z(n_0_118));
   MUX2_X1 i_0_1_22 (.A(c[23]), .B(b[23]), .S(start_s), .Z(n_0_119));
   AND2_X1 i_0_1_23 (.A1(start_s), .A2(b[0]), .ZN(n_0_1_0));
   AND2_X1 i_0_1_24 (.A1(n_0_1_26), .A2(c[0]), .ZN(n_0_1_1));
   AOI22_X1 i_0_1_25 (.A1(a[0]), .A2(n_0_1_0), .B1(A_r[0]), .B2(n_0_1_1), 
      .ZN(n_0_1_2));
   INV_X1 i_0_1_26 (.A(n_0_1_2), .ZN(n_0_49));
   AOI22_X1 i_0_1_27 (.A1(a[1]), .A2(n_0_1_0), .B1(A_r[1]), .B2(n_0_1_1), 
      .ZN(n_0_1_3));
   INV_X1 i_0_1_28 (.A(n_0_1_3), .ZN(n_0_50));
   AOI22_X1 i_0_1_29 (.A1(a[2]), .A2(n_0_1_0), .B1(A_r[2]), .B2(n_0_1_1), 
      .ZN(n_0_1_4));
   INV_X1 i_0_1_30 (.A(n_0_1_4), .ZN(n_0_51));
   AOI22_X1 i_0_1_31 (.A1(a[3]), .A2(n_0_1_0), .B1(A_r[3]), .B2(n_0_1_1), 
      .ZN(n_0_1_5));
   INV_X1 i_0_1_32 (.A(n_0_1_5), .ZN(n_0_52));
   AOI22_X1 i_0_1_33 (.A1(a[4]), .A2(n_0_1_0), .B1(A_r[4]), .B2(n_0_1_1), 
      .ZN(n_0_1_6));
   INV_X1 i_0_1_34 (.A(n_0_1_6), .ZN(n_0_53));
   AOI22_X1 i_0_1_35 (.A1(a[5]), .A2(n_0_1_0), .B1(A_r[5]), .B2(n_0_1_1), 
      .ZN(n_0_1_7));
   INV_X1 i_0_1_36 (.A(n_0_1_7), .ZN(n_0_54));
   AOI22_X1 i_0_1_37 (.A1(a[6]), .A2(n_0_1_0), .B1(A_r[6]), .B2(n_0_1_1), 
      .ZN(n_0_1_8));
   INV_X1 i_0_1_38 (.A(n_0_1_8), .ZN(n_0_55));
   AOI22_X1 i_0_1_39 (.A1(a[7]), .A2(n_0_1_0), .B1(A_r[7]), .B2(n_0_1_1), 
      .ZN(n_0_1_9));
   INV_X1 i_0_1_40 (.A(n_0_1_9), .ZN(n_0_56));
   AOI22_X1 i_0_1_41 (.A1(a[8]), .A2(n_0_1_0), .B1(A_r[8]), .B2(n_0_1_1), 
      .ZN(n_0_1_10));
   INV_X1 i_0_1_42 (.A(n_0_1_10), .ZN(n_0_57));
   AOI22_X1 i_0_1_43 (.A1(a[9]), .A2(n_0_1_0), .B1(A_r[9]), .B2(n_0_1_1), 
      .ZN(n_0_1_11));
   INV_X1 i_0_1_44 (.A(n_0_1_11), .ZN(n_0_58));
   AOI22_X1 i_0_1_45 (.A1(a[10]), .A2(n_0_1_0), .B1(A_r[10]), .B2(n_0_1_1), 
      .ZN(n_0_1_12));
   INV_X1 i_0_1_46 (.A(n_0_1_12), .ZN(n_0_59));
   AOI22_X1 i_0_1_47 (.A1(a[11]), .A2(n_0_1_0), .B1(A_r[11]), .B2(n_0_1_1), 
      .ZN(n_0_1_13));
   INV_X1 i_0_1_48 (.A(n_0_1_13), .ZN(n_0_60));
   AOI22_X1 i_0_1_49 (.A1(a[12]), .A2(n_0_1_0), .B1(A_r[12]), .B2(n_0_1_1), 
      .ZN(n_0_1_14));
   INV_X1 i_0_1_50 (.A(n_0_1_14), .ZN(n_0_61));
   AOI22_X1 i_0_1_51 (.A1(a[13]), .A2(n_0_1_0), .B1(A_r[13]), .B2(n_0_1_1), 
      .ZN(n_0_1_15));
   INV_X1 i_0_1_52 (.A(n_0_1_15), .ZN(n_0_62));
   AOI22_X1 i_0_1_53 (.A1(a[14]), .A2(n_0_1_0), .B1(A_r[14]), .B2(n_0_1_1), 
      .ZN(n_0_1_16));
   INV_X1 i_0_1_54 (.A(n_0_1_16), .ZN(n_0_63));
   AOI22_X1 i_0_1_55 (.A1(a[15]), .A2(n_0_1_0), .B1(A_r[15]), .B2(n_0_1_1), 
      .ZN(n_0_1_17));
   INV_X1 i_0_1_56 (.A(n_0_1_17), .ZN(n_0_64));
   AOI22_X1 i_0_1_57 (.A1(a[16]), .A2(n_0_1_0), .B1(A_r[16]), .B2(n_0_1_1), 
      .ZN(n_0_1_18));
   INV_X1 i_0_1_58 (.A(n_0_1_18), .ZN(n_0_65));
   AOI22_X1 i_0_1_59 (.A1(a[17]), .A2(n_0_1_0), .B1(A_r[17]), .B2(n_0_1_1), 
      .ZN(n_0_1_19));
   INV_X1 i_0_1_60 (.A(n_0_1_19), .ZN(n_0_66));
   AOI22_X1 i_0_1_61 (.A1(a[18]), .A2(n_0_1_0), .B1(A_r[18]), .B2(n_0_1_1), 
      .ZN(n_0_1_20));
   INV_X1 i_0_1_62 (.A(n_0_1_20), .ZN(n_0_67));
   AOI22_X1 i_0_1_63 (.A1(a[19]), .A2(n_0_1_0), .B1(A_r[19]), .B2(n_0_1_1), 
      .ZN(n_0_1_21));
   INV_X1 i_0_1_64 (.A(n_0_1_21), .ZN(n_0_68));
   AOI22_X1 i_0_1_65 (.A1(a[20]), .A2(n_0_1_0), .B1(A_r[20]), .B2(n_0_1_1), 
      .ZN(n_0_1_22));
   INV_X1 i_0_1_66 (.A(n_0_1_22), .ZN(n_0_69));
   AOI22_X1 i_0_1_67 (.A1(a[21]), .A2(n_0_1_0), .B1(A_r[21]), .B2(n_0_1_1), 
      .ZN(n_0_1_23));
   INV_X1 i_0_1_68 (.A(n_0_1_23), .ZN(n_0_70));
   AOI22_X1 i_0_1_69 (.A1(a[22]), .A2(n_0_1_0), .B1(A_r[22]), .B2(n_0_1_1), 
      .ZN(n_0_1_24));
   INV_X1 i_0_1_70 (.A(n_0_1_24), .ZN(n_0_71));
   AOI22_X1 i_0_1_71 (.A1(a[23]), .A2(n_0_1_0), .B1(A_r[23]), .B2(n_0_1_1), 
      .ZN(n_0_1_25));
   INV_X1 i_0_1_72 (.A(n_0_1_25), .ZN(n_0_96));
   AND2_X1 i_0_1_73 (.A1(n_0_1_26), .A2(c[24]), .ZN(n_0_26));
   AND2_X1 i_0_1_74 (.A1(n_0_1_26), .A2(c[25]), .ZN(n_0_27));
   AND2_X1 i_0_1_75 (.A1(n_0_1_26), .A2(c[26]), .ZN(n_0_28));
   AND2_X1 i_0_1_76 (.A1(n_0_1_26), .A2(c[27]), .ZN(n_0_29));
   AND2_X1 i_0_1_77 (.A1(n_0_1_26), .A2(c[28]), .ZN(n_0_30));
   AND2_X1 i_0_1_78 (.A1(n_0_1_26), .A2(c[29]), .ZN(n_0_31));
   AND2_X1 i_0_1_79 (.A1(n_0_1_26), .A2(c[30]), .ZN(n_0_32));
   AND2_X1 i_0_1_80 (.A1(n_0_1_26), .A2(c[31]), .ZN(n_0_33));
   AND2_X1 i_0_1_81 (.A1(n_0_1_26), .A2(c[32]), .ZN(n_0_34));
   AND2_X1 i_0_1_82 (.A1(n_0_1_26), .A2(c[33]), .ZN(n_0_35));
   AND2_X1 i_0_1_83 (.A1(n_0_1_26), .A2(c[34]), .ZN(n_0_36));
   AND2_X1 i_0_1_84 (.A1(n_0_1_26), .A2(c[35]), .ZN(n_0_37));
   AND2_X1 i_0_1_85 (.A1(n_0_1_26), .A2(c[36]), .ZN(n_0_38));
   AND2_X1 i_0_1_86 (.A1(n_0_1_26), .A2(c[37]), .ZN(n_0_39));
   AND2_X1 i_0_1_87 (.A1(n_0_1_26), .A2(c[38]), .ZN(n_0_40));
   AND2_X1 i_0_1_88 (.A1(n_0_1_26), .A2(c[39]), .ZN(n_0_41));
   AND2_X1 i_0_1_89 (.A1(n_0_1_26), .A2(c[40]), .ZN(n_0_42));
   AND2_X1 i_0_1_90 (.A1(n_0_1_26), .A2(c[41]), .ZN(n_0_43));
   AND2_X1 i_0_1_91 (.A1(n_0_1_26), .A2(c[42]), .ZN(n_0_44));
   AND2_X1 i_0_1_92 (.A1(n_0_1_26), .A2(c[43]), .ZN(n_0_45));
   AND2_X1 i_0_1_93 (.A1(n_0_1_26), .A2(c[44]), .ZN(n_0_46));
   AND2_X1 i_0_1_94 (.A1(n_0_1_26), .A2(c[45]), .ZN(n_0_47));
   AND2_X1 i_0_1_95 (.A1(n_0_1_26), .A2(c[46]), .ZN(n_0_48));
   MUX2_X1 i_0_1_96 (.A(A_r[0]), .B(a[0]), .S(start_s), .Z(n_0_2));
   MUX2_X1 i_0_1_97 (.A(A_r[1]), .B(a[1]), .S(start_s), .Z(n_0_3));
   MUX2_X1 i_0_1_98 (.A(A_r[2]), .B(a[2]), .S(start_s), .Z(n_0_4));
   MUX2_X1 i_0_1_99 (.A(A_r[3]), .B(a[3]), .S(start_s), .Z(n_0_5));
   MUX2_X1 i_0_1_100 (.A(A_r[4]), .B(a[4]), .S(start_s), .Z(n_0_6));
   MUX2_X1 i_0_1_101 (.A(A_r[5]), .B(a[5]), .S(start_s), .Z(n_0_7));
   MUX2_X1 i_0_1_102 (.A(A_r[6]), .B(a[6]), .S(start_s), .Z(n_0_8));
   MUX2_X1 i_0_1_103 (.A(A_r[7]), .B(a[7]), .S(start_s), .Z(n_0_9));
   MUX2_X1 i_0_1_104 (.A(A_r[8]), .B(a[8]), .S(start_s), .Z(n_0_10));
   MUX2_X1 i_0_1_105 (.A(A_r[9]), .B(a[9]), .S(start_s), .Z(n_0_11));
   MUX2_X1 i_0_1_106 (.A(A_r[10]), .B(a[10]), .S(start_s), .Z(n_0_12));
   MUX2_X1 i_0_1_107 (.A(A_r[11]), .B(a[11]), .S(start_s), .Z(n_0_13));
   MUX2_X1 i_0_1_108 (.A(A_r[12]), .B(a[12]), .S(start_s), .Z(n_0_14));
   MUX2_X1 i_0_1_109 (.A(A_r[13]), .B(a[13]), .S(start_s), .Z(n_0_15));
   MUX2_X1 i_0_1_110 (.A(A_r[14]), .B(a[14]), .S(start_s), .Z(n_0_16));
   MUX2_X1 i_0_1_111 (.A(A_r[15]), .B(a[15]), .S(start_s), .Z(n_0_17));
   MUX2_X1 i_0_1_112 (.A(A_r[16]), .B(a[16]), .S(start_s), .Z(n_0_18));
   MUX2_X1 i_0_1_113 (.A(A_r[17]), .B(a[17]), .S(start_s), .Z(n_0_19));
   MUX2_X1 i_0_1_114 (.A(A_r[18]), .B(a[18]), .S(start_s), .Z(n_0_20));
   MUX2_X1 i_0_1_115 (.A(A_r[19]), .B(a[19]), .S(start_s), .Z(n_0_21));
   MUX2_X1 i_0_1_116 (.A(A_r[20]), .B(a[20]), .S(start_s), .Z(n_0_22));
   MUX2_X1 i_0_1_117 (.A(A_r[21]), .B(a[21]), .S(start_s), .Z(n_0_23));
   MUX2_X1 i_0_1_118 (.A(A_r[22]), .B(a[22]), .S(start_s), .Z(n_0_24));
   MUX2_X1 i_0_1_119 (.A(A_r[23]), .B(a[23]), .S(start_s), .Z(n_0_25));
   INV_X1 i_0_1_120 (.A(start_s), .ZN(n_0_1_26));
endmodule
