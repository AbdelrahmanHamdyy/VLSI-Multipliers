
// 	Fri Dec 23 03:48:35 2022
//	vlsi
//	localhost.localdomain

module datapath__0_72 (p_0, p_1);

output [63:0] p_0;
input [63:0] p_1;
wire n_127;
wire n_125;
wire n_126;
wire n_123;
wire n_124;
wire n_5;
wire n_122;
wire n_3;
wire n_4;
wire n_1;
wire n_2;
wire n_120;
wire n_0;
wire n_121;
wire n_11;
wire n_119;
wire n_9;
wire n_10;
wire n_7;
wire n_8;
wire n_117;
wire n_6;
wire n_118;
wire n_17;
wire n_15;
wire n_16;
wire n_13;
wire n_14;
wire n_114;
wire n_12;
wire n_115;
wire n_112;
wire n_113;
wire n_110;
wire n_108;
wire n_109;
wire n_106;
wire n_107;
wire n_104;
wire n_105;
wire n_102;
wire n_103;
wire n_100;
wire n_101;
wire n_98;
wire n_99;
wire n_96;
wire n_97;
wire n_94;
wire n_92;
wire n_93;
wire n_90;
wire n_91;
wire n_88;
wire n_89;
wire n_86;
wire n_84;
wire n_85;
wire n_82;
wire n_83;
wire n_23;
wire n_81;
wire n_21;
wire n_22;
wire n_19;
wire n_20;
wire n_31;
wire n_18;
wire n_29;
wire n_30;
wire n_27;
wire n_28;
wire n_25;
wire n_26;
wire n_77;
wire n_24;
wire n_79;
wire n_37;
wire n_76;
wire n_35;
wire n_36;
wire n_33;
wire n_34;
wire n_75;
wire n_32;
wire n_80;
wire n_73;
wire n_74;
wire n_71;
wire n_72;
wire n_69;
wire n_70;
wire n_67;
wire n_68;
wire n_43;
wire n_66;
wire n_41;
wire n_42;
wire n_39;
wire n_40;
wire n_38;
wire n_49;
wire n_128;
wire n_45;
wire n_44;
wire n_46;
wire n_129;
wire n_48;
wire n_62;
wire n_47;
wire n_63;
wire n_64;
wire n_51;
wire n_61;
wire n_50;
wire n_52;
wire n_130;
wire n_54;
wire n_60;
wire n_53;
wire n_65;
wire n_134;
wire n_132;
wire n_78;
wire n_155;
wire n_169;
wire n_58;
wire n_55;
wire n_57;
wire n_56;
wire n_59;
wire n_168;
wire n_167;
wire n_131;
wire n_157;
wire n_156;
wire n_196;
wire n_193;
wire n_192;
wire n_135;
wire n_187;
wire n_184;
wire n_181;
wire n_178;
wire n_136;
wire n_175;
wire n_163;
wire n_162;
wire n_161;
wire n_165;
wire n_173;
wire n_172;
wire n_171;
wire n_137;
wire n_145;
wire n_138;
wire n_139;
wire n_198;
wire n_197;
wire n_142;
wire n_140;
wire n_141;
wire n_146;
wire n_195;
wire n_148;
wire n_194;
wire n_191;
wire n_189;
wire n_190;
wire n_188;
wire n_186;
wire n_185;
wire n_183;
wire n_182;
wire n_180;
wire n_179;
wire n_177;
wire n_176;
wire n_153;
wire n_144;
wire n_159;
wire n_199;
wire n_147;
wire n_149;
wire n_150;
wire n_154;
wire n_158;
wire n_160;
wire n_164;
wire n_166;
wire n_170;
wire n_174;


INV_X1 i_262 (.ZN (n_199), .A (p_1[62]));
INV_X1 i_261 (.ZN (n_198), .A (p_1[61]));
INV_X1 i_260 (.ZN (n_197), .A (p_1[60]));
INV_X1 i_259 (.ZN (n_196), .A (p_1[47]));
INV_X1 i_258 (.ZN (n_195), .A (p_1[46]));
INV_X1 i_257 (.ZN (n_194), .A (p_1[45]));
INV_X1 i_256 (.ZN (n_193), .A (p_1[44]));
INV_X1 i_255 (.ZN (n_192), .A (p_1[31]));
INV_X1 i_254 (.ZN (n_191), .A (n_55));
INV_X1 i_253 (.ZN (n_190), .A (n_56));
INV_X1 i_252 (.ZN (n_189), .A (p_1[30]));
INV_X1 i_251 (.ZN (n_188), .A (p_1[29]));
INV_X1 i_250 (.ZN (n_187), .A (p_1[28]));
INV_X1 i_249 (.ZN (n_186), .A (p_1[27]));
INV_X1 i_248 (.ZN (n_185), .A (p_1[26]));
INV_X1 i_247 (.ZN (n_184), .A (p_1[25]));
INV_X1 i_246 (.ZN (n_183), .A (p_1[24]));
INV_X1 i_245 (.ZN (n_182), .A (p_1[23]));
INV_X1 i_244 (.ZN (n_181), .A (p_1[22]));
INV_X1 i_243 (.ZN (n_180), .A (p_1[21]));
INV_X1 i_242 (.ZN (n_179), .A (p_1[20]));
INV_X1 i_241 (.ZN (n_178), .A (p_1[19]));
INV_X1 i_240 (.ZN (n_177), .A (p_1[18]));
INV_X1 i_239 (.ZN (n_176), .A (p_1[17]));
INV_X1 i_238 (.ZN (n_175), .A (p_1[16]));
INV_X1 i_237 (.ZN (n_174), .A (p_1[3]));
INV_X1 i_236 (.ZN (n_173), .A (p_1[2]));
INV_X1 i_235 (.ZN (n_172), .A (p_1[1]));
INV_X1 i_234 (.ZN (n_171), .A (p_1[0]));
NAND4_X1 i_233 (.ZN (n_122), .A1 (n_174), .A2 (n_173), .A3 (n_172), .A4 (n_171));
INV_X1 i_232 (.ZN (n_123), .A (n_122));
INV_X1 i_231 (.ZN (n_170), .A (p_1[7]));
INV_X1 i_230 (.ZN (n_169), .A (p_1[6]));
INV_X1 i_229 (.ZN (n_168), .A (p_1[5]));
INV_X1 i_228 (.ZN (n_167), .A (p_1[4]));
NAND4_X1 i_227 (.ZN (n_166), .A1 (n_170), .A2 (n_169), .A3 (n_168), .A4 (n_167));
INV_X1 i_226 (.ZN (n_165), .A (n_166));
INV_X1 i_225 (.ZN (n_164), .A (p_1[11]));
INV_X1 i_224 (.ZN (n_163), .A (p_1[10]));
INV_X1 i_223 (.ZN (n_162), .A (p_1[9]));
INV_X1 i_222 (.ZN (n_161), .A (p_1[8]));
NAND4_X1 i_221 (.ZN (n_160), .A1 (n_164), .A2 (n_163), .A3 (n_162), .A4 (n_161));
INV_X1 i_220 (.ZN (n_159), .A (n_160));
INV_X1 i_219 (.ZN (n_158), .A (p_1[15]));
INV_X1 i_218 (.ZN (n_157), .A (p_1[14]));
INV_X1 i_217 (.ZN (n_156), .A (p_1[13]));
INV_X1 i_216 (.ZN (n_155), .A (p_1[12]));
NAND4_X1 i_215 (.ZN (n_154), .A1 (n_158), .A2 (n_157), .A3 (n_156), .A4 (n_155));
INV_X1 i_214 (.ZN (n_153), .A (n_154));
NAND4_X1 i_213 (.ZN (n_113), .A1 (n_123), .A2 (n_165), .A3 (n_159), .A4 (n_153));
NAND4_X1 i_211 (.ZN (n_107), .A1 (n_114), .A2 (n_177), .A3 (n_176), .A4 (n_175));
NAND4_X1 i_209 (.ZN (n_101), .A1 (n_108), .A2 (n_180), .A3 (n_179), .A4 (n_178));
INV_X1 i_208 (.ZN (n_102), .A (n_101));
NAND4_X1 i_207 (.ZN (n_150), .A1 (n_102), .A2 (n_183), .A3 (n_182), .A4 (n_181));
INV_X1 i_206 (.ZN (n_96), .A (n_150));
NAND4_X1 i_205 (.ZN (n_89), .A1 (n_96), .A2 (n_186), .A3 (n_185), .A4 (n_184));
INV_X1 i_204 (.ZN (n_90), .A (n_89));
NAND4_X1 i_203 (.ZN (n_83), .A1 (n_90), .A2 (n_189), .A3 (n_188), .A4 (n_187));
INV_X1 i_202 (.ZN (n_84), .A (n_83));
NAND4_X1 i_201 (.ZN (n_74), .A1 (n_84), .A2 (n_192), .A3 (n_191), .A4 (n_190));
INV_X1 i_200 (.ZN (n_75), .A (n_74));
NAND4_X1 i_199 (.ZN (n_68), .A1 (n_75), .A2 (n_195), .A3 (n_194), .A4 (n_193));
INV_X1 i_198 (.ZN (n_69), .A (n_68));
OR4_X1 i_197 (.ZN (n_64), .A1 (p_1[51]), .A2 (p_1[50]), .A3 (p_1[49]), .A4 (p_1[48]));
OR3_X2 i_196 (.ZN (n_63), .A1 (p_1[54]), .A2 (p_1[53]), .A3 (p_1[52]));
OR3_X2 i_195 (.ZN (n_149), .A1 (n_64), .A2 (n_63), .A3 (p_1[55]));
INV_X2 i_194 (.ZN (n_148), .A (n_149));
OR4_X1 i_190 (.ZN (n_147), .A1 (p_1[59]), .A2 (p_1[58]), .A3 (p_1[57]), .A4 (p_1[56]));
INV_X1 i_189 (.ZN (n_146), .A (n_147));
NAND4_X1 i_188 (.ZN (n_145), .A1 (n_69), .A2 (n_196), .A3 (n_148), .A4 (n_146));
INV_X1 i_187 (.ZN (n_60), .A (n_145));
NAND4_X1 i_186 (.ZN (p_0[63]), .A1 (n_60), .A2 (n_199), .A3 (n_198), .A4 (n_197));
NAND3_X1 i_185 (.ZN (n_144), .A1 (n_123), .A2 (n_165), .A3 (n_159));
INV_X1 i_184 (.ZN (n_117), .A (n_144));
NAND4_X1 i_183 (.ZN (n_109), .A1 (n_117), .A2 (n_176), .A3 (n_175), .A4 (n_153));
INV_X1 i_182 (.ZN (n_110), .A (n_109));
NAND4_X1 i_181 (.ZN (n_103), .A1 (n_110), .A2 (n_179), .A3 (n_178), .A4 (n_177));
INV_X1 i_180 (.ZN (n_104), .A (n_103));
NAND4_X1 i_179 (.ZN (n_97), .A1 (n_104), .A2 (n_182), .A3 (n_181), .A4 (n_180));
INV_X1 i_178 (.ZN (n_98), .A (n_97));
NAND4_X1 i_177 (.ZN (n_91), .A1 (n_98), .A2 (n_185), .A3 (n_184), .A4 (n_183));
NAND4_X1 i_175 (.ZN (n_85), .A1 (n_92), .A2 (n_188), .A3 (n_187), .A4 (n_186));
INV_X1 i_174 (.ZN (n_86), .A (n_85));
NAND4_X1 i_173 (.ZN (n_76), .A1 (n_86), .A2 (n_192), .A3 (n_189), .A4 (n_190));
INV_X1 i_172 (.ZN (n_77), .A (n_76));
NAND4_X1 i_171 (.ZN (n_70), .A1 (n_77), .A2 (n_194), .A3 (n_193), .A4 (n_191));
INV_X1 i_170 (.ZN (n_71), .A (n_70));
NAND4_X2 i_169 (.ZN (n_61), .A1 (n_71), .A2 (n_196), .A3 (n_195), .A4 (n_148));
INV_X1 i_168 (.ZN (n_62), .A (n_61));
NAND4_X1 i_167 (.ZN (n_142), .A1 (n_62), .A2 (n_198), .A3 (n_197), .A4 (n_146));
NAND2_X1 i_166 (.ZN (n_141), .A1 (n_142), .A2 (p_1[62]));
NAND2_X1 i_165 (.ZN (n_140), .A1 (n_141), .A2 (p_0[63]));
INV_X1 i_164 (.ZN (p_0[62]), .A (n_140));
INV_X1 i_163 (.ZN (n_139), .A (n_142));
AOI21_X1 i_162 (.ZN (n_138), .A (n_198), .B1 (n_60), .B2 (n_197));
NOR2_X1 i_161 (.ZN (p_0[61]), .A1 (n_138), .A2 (n_139));
XNOR2_X1 i_160 (.ZN (n_137), .A (n_145), .B (p_1[60]));
INV_X1 i_159 (.ZN (p_0[60]), .A (n_137));
NAND2_X1 i_158 (.ZN (n_126), .A1 (n_172), .A2 (n_171));
INV_X1 i_157 (.ZN (n_127), .A (n_126));
NAND2_X1 i_156 (.ZN (n_124), .A1 (n_127), .A2 (n_173));
INV_X1 i_155 (.ZN (n_125), .A (n_124));
NAND2_X1 i_154 (.ZN (n_119), .A1 (n_123), .A2 (n_165));
NAND3_X1 i_153 (.ZN (n_118), .A1 (n_163), .A2 (n_162), .A3 (n_161));
NAND2_X1 i_152 (.ZN (n_136), .A1 (n_114), .A2 (n_175));
INV_X1 i_151 (.ZN (n_112), .A (n_136));
NAND2_X1 i_150 (.ZN (n_105), .A1 (n_108), .A2 (n_178));
INV_X1 i_149 (.ZN (n_106), .A (n_105));
NAND2_X1 i_148 (.ZN (n_99), .A1 (n_102), .A2 (n_181));
INV_X1 i_147 (.ZN (n_100), .A (n_99));
NAND2_X1 i_146 (.ZN (n_93), .A1 (n_96), .A2 (n_184));
INV_X1 i_145 (.ZN (n_94), .A (n_93));
NAND2_X1 i_144 (.ZN (n_135), .A1 (n_90), .A2 (n_187));
INV_X1 i_143 (.ZN (n_88), .A (n_135));
NAND2_X1 i_142 (.ZN (n_81), .A1 (n_84), .A2 (n_192));
INV_X1 i_141 (.ZN (n_82), .A (n_81));
NAND2_X1 i_140 (.ZN (n_72), .A1 (n_75), .A2 (n_193));
INV_X1 i_139 (.ZN (n_73), .A (n_72));
NAND2_X1 i_138 (.ZN (n_66), .A1 (n_69), .A2 (n_196));
INV_X1 i_137 (.ZN (n_134), .A (p_1[58]));
INV_X1 i_135 (.ZN (n_132), .A (p_1[56]));
NAND2_X1 i_134 (.ZN (n_131), .A1 (n_157), .A2 (n_156));
INV_X1 i_133 (.ZN (n_78), .A (n_131));
NAND2_X1 i_132 (.ZN (n_59), .A1 (n_168), .A2 (n_167));
INV_X1 i_131 (.ZN (n_58), .A (n_59));
OR4_X1 i_130 (.ZN (n_79), .A1 (p_1[35]), .A2 (p_1[34]), .A3 (p_1[33]), .A4 (p_1[32]));
OR2_X1 i_129 (.ZN (n_57), .A1 (n_79), .A2 (p_1[36]));
OR4_X1 i_128 (.ZN (n_56), .A1 (p_1[39]), .A2 (n_57), .A3 (p_1[38]), .A4 (p_1[37]));
OR3_X1 i_127 (.ZN (n_80), .A1 (p_1[42]), .A2 (p_1[41]), .A3 (p_1[40]));
OR2_X1 i_126 (.ZN (n_55), .A1 (n_80), .A2 (p_1[43]));
INV_X1 i_125 (.ZN (n_120), .A (n_119));
NAND2_X1 i_124 (.ZN (n_121), .A1 (n_169), .A2 (n_58));
INV_X1 i_122 (.ZN (n_114), .A (n_113));
NAND2_X1 i_121 (.ZN (n_115), .A1 (n_78), .A2 (n_155));
INV_X1 i_119 (.ZN (n_108), .A (n_107));
INV_X1 i_117 (.ZN (n_92), .A (n_91));
INV_X1 i_115 (.ZN (n_67), .A (n_66));
NAND3_X1 i_114 (.ZN (n_65), .A1 (n_134), .A2 (n_130), .A3 (n_132));
INV_X1 i_193 (.ZN (n_130), .A (p_1[57]));
INV_X1 i_192 (.ZN (n_129), .A (p_1[53]));
INV_X1 i_191 (.ZN (n_128), .A (p_1[51]));
NOR2_X1 i_113 (.ZN (n_54), .A1 (n_65), .A2 (n_61));
INV_X1 i_112 (.ZN (n_53), .A (n_54));
AOI21_X1 i_111 (.ZN (p_0[59]), .A (n_60), .B1 (p_1[59]), .B2 (n_53));
OR3_X1 i_110 (.ZN (n_52), .A1 (p_1[57]), .A2 (p_1[56]), .A3 (n_61));
AOI21_X1 i_109 (.ZN (p_0[58]), .A (n_54), .B1 (p_1[58]), .B2 (n_52));
NOR2_X1 i_108 (.ZN (n_51), .A1 (p_1[56]), .A2 (n_61));
OAI21_X1 i_107 (.ZN (n_50), .A (n_52), .B1 (n_130), .B2 (n_51));
INV_X1 i_106 (.ZN (p_0[57]), .A (n_50));
AOI21_X1 i_105 (.ZN (p_0[56]), .A (n_51), .B1 (p_1[56]), .B2 (n_61));
OR2_X1 i_104 (.ZN (n_49), .A1 (n_66), .A2 (n_64));
NOR2_X1 i_103 (.ZN (n_48), .A1 (n_63), .A2 (n_49));
INV_X1 i_102 (.ZN (n_47), .A (n_48));
AOI21_X1 i_101 (.ZN (p_0[55]), .A (n_62), .B1 (p_1[55]), .B2 (n_47));
OR3_X1 i_100 (.ZN (n_46), .A1 (p_1[53]), .A2 (p_1[52]), .A3 (n_49));
AOI21_X1 i_99 (.ZN (p_0[54]), .A (n_48), .B1 (p_1[54]), .B2 (n_46));
NOR2_X1 i_98 (.ZN (n_45), .A1 (p_1[52]), .A2 (n_49));
OAI21_X1 i_97 (.ZN (n_44), .A (n_46), .B1 (n_129), .B2 (n_45));
INV_X1 i_96 (.ZN (p_0[53]), .A (n_44));
AOI21_X1 i_95 (.ZN (p_0[52]), .A (n_45), .B1 (p_1[52]), .B2 (n_49));
NOR2_X1 i_94 (.ZN (n_43), .A1 (p_1[48]), .A2 (n_66));
INV_X1 i_93 (.ZN (n_42), .A (n_43));
NOR2_X1 i_92 (.ZN (n_41), .A1 (p_1[49]), .A2 (n_42));
INV_X1 i_91 (.ZN (n_40), .A (n_41));
NOR2_X1 i_90 (.ZN (n_39), .A1 (p_1[50]), .A2 (n_40));
OAI21_X1 i_89 (.ZN (n_38), .A (n_49), .B1 (n_128), .B2 (n_39));
INV_X1 i_88 (.ZN (p_0[51]), .A (n_38));
AOI21_X1 i_87 (.ZN (p_0[50]), .A (n_39), .B1 (p_1[50]), .B2 (n_40));
AOI21_X1 i_86 (.ZN (p_0[49]), .A (n_41), .B1 (p_1[49]), .B2 (n_42));
AOI21_X1 i_85 (.ZN (p_0[48]), .A (n_43), .B1 (p_1[48]), .B2 (n_66));
AOI21_X1 i_84 (.ZN (p_0[47]), .A (n_67), .B1 (p_1[47]), .B2 (n_68));
AOI21_X1 i_83 (.ZN (p_0[46]), .A (n_69), .B1 (p_1[46]), .B2 (n_70));
AOI21_X1 i_82 (.ZN (p_0[45]), .A (n_71), .B1 (p_1[45]), .B2 (n_72));
AOI21_X1 i_81 (.ZN (p_0[44]), .A (n_73), .B1 (p_1[44]), .B2 (n_74));
NOR2_X1 i_80 (.ZN (n_37), .A1 (p_1[40]), .A2 (n_76));
INV_X1 i_79 (.ZN (n_36), .A (n_37));
NOR2_X1 i_78 (.ZN (n_35), .A1 (p_1[41]), .A2 (n_36));
INV_X1 i_77 (.ZN (n_34), .A (n_35));
NOR2_X1 i_76 (.ZN (n_33), .A1 (n_80), .A2 (n_76));
INV_X1 i_75 (.ZN (n_32), .A (n_33));
AOI21_X1 i_74 (.ZN (p_0[43]), .A (n_75), .B1 (p_1[43]), .B2 (n_32));
AOI21_X1 i_73 (.ZN (p_0[42]), .A (n_33), .B1 (p_1[42]), .B2 (n_34));
AOI21_X1 i_72 (.ZN (p_0[41]), .A (n_35), .B1 (p_1[41]), .B2 (n_36));
AOI21_X1 i_71 (.ZN (p_0[40]), .A (n_37), .B1 (p_1[40]), .B2 (n_76));
NOR2_X1 i_70 (.ZN (n_31), .A1 (n_81), .A2 (n_79));
INV_X1 i_69 (.ZN (n_30), .A (n_31));
NOR2_X1 i_68 (.ZN (n_29), .A1 (p_1[36]), .A2 (n_30));
INV_X1 i_67 (.ZN (n_28), .A (n_29));
NOR2_X1 i_66 (.ZN (n_27), .A1 (p_1[37]), .A2 (n_28));
INV_X1 i_65 (.ZN (n_26), .A (n_27));
NOR2_X1 i_64 (.ZN (n_25), .A1 (p_1[38]), .A2 (n_26));
INV_X1 i_63 (.ZN (n_24), .A (n_25));
AOI21_X1 i_62 (.ZN (p_0[39]), .A (n_77), .B1 (p_1[39]), .B2 (n_24));
AOI21_X1 i_61 (.ZN (p_0[38]), .A (n_25), .B1 (p_1[38]), .B2 (n_26));
AOI21_X1 i_60 (.ZN (p_0[37]), .A (n_27), .B1 (p_1[37]), .B2 (n_28));
AOI21_X1 i_59 (.ZN (p_0[36]), .A (n_29), .B1 (p_1[36]), .B2 (n_30));
NOR2_X1 i_58 (.ZN (n_23), .A1 (p_1[32]), .A2 (n_81));
INV_X1 i_57 (.ZN (n_22), .A (n_23));
NOR2_X1 i_56 (.ZN (n_21), .A1 (p_1[33]), .A2 (n_22));
INV_X1 i_55 (.ZN (n_20), .A (n_21));
NOR2_X1 i_54 (.ZN (n_19), .A1 (p_1[34]), .A2 (n_20));
INV_X1 i_53 (.ZN (n_18), .A (n_19));
AOI21_X1 i_52 (.ZN (p_0[35]), .A (n_31), .B1 (p_1[35]), .B2 (n_18));
AOI21_X1 i_51 (.ZN (p_0[34]), .A (n_19), .B1 (p_1[34]), .B2 (n_20));
AOI21_X1 i_50 (.ZN (p_0[33]), .A (n_21), .B1 (p_1[33]), .B2 (n_22));
AOI21_X1 i_49 (.ZN (p_0[32]), .A (n_23), .B1 (p_1[32]), .B2 (n_81));
AOI21_X1 i_48 (.ZN (p_0[31]), .A (n_82), .B1 (p_1[31]), .B2 (n_83));
AOI21_X1 i_47 (.ZN (p_0[30]), .A (n_84), .B1 (p_1[30]), .B2 (n_85));
AOI21_X1 i_46 (.ZN (p_0[29]), .A (n_86), .B1 (p_1[29]), .B2 (n_135));
AOI21_X1 i_45 (.ZN (p_0[28]), .A (n_88), .B1 (p_1[28]), .B2 (n_89));
AOI21_X1 i_44 (.ZN (p_0[27]), .A (n_90), .B1 (p_1[27]), .B2 (n_91));
AOI21_X1 i_43 (.ZN (p_0[26]), .A (n_92), .B1 (p_1[26]), .B2 (n_93));
AOI21_X1 i_42 (.ZN (p_0[25]), .A (n_94), .B1 (p_1[25]), .B2 (n_150));
AOI21_X1 i_41 (.ZN (p_0[24]), .A (n_96), .B1 (p_1[24]), .B2 (n_97));
AOI21_X1 i_40 (.ZN (p_0[23]), .A (n_98), .B1 (p_1[23]), .B2 (n_99));
AOI21_X1 i_39 (.ZN (p_0[22]), .A (n_100), .B1 (p_1[22]), .B2 (n_101));
AOI21_X1 i_38 (.ZN (p_0[21]), .A (n_102), .B1 (p_1[21]), .B2 (n_103));
AOI21_X1 i_37 (.ZN (p_0[20]), .A (n_104), .B1 (p_1[20]), .B2 (n_105));
AOI21_X1 i_36 (.ZN (p_0[19]), .A (n_106), .B1 (p_1[19]), .B2 (n_107));
AOI21_X1 i_35 (.ZN (p_0[18]), .A (n_108), .B1 (p_1[18]), .B2 (n_109));
AOI21_X1 i_34 (.ZN (p_0[17]), .A (n_110), .B1 (p_1[17]), .B2 (n_136));
AOI21_X1 i_33 (.ZN (p_0[16]), .A (n_112), .B1 (p_1[16]), .B2 (n_113));
NOR2_X1 i_32 (.ZN (n_17), .A1 (p_1[12]), .A2 (n_144));
INV_X1 i_31 (.ZN (n_16), .A (n_17));
NOR2_X1 i_30 (.ZN (n_15), .A1 (p_1[13]), .A2 (n_16));
INV_X1 i_29 (.ZN (n_14), .A (n_15));
NOR2_X1 i_28 (.ZN (n_13), .A1 (n_144), .A2 (n_115));
INV_X1 i_27 (.ZN (n_12), .A (n_13));
AOI21_X1 i_26 (.ZN (p_0[15]), .A (n_114), .B1 (p_1[15]), .B2 (n_12));
AOI21_X1 i_25 (.ZN (p_0[14]), .A (n_13), .B1 (p_1[14]), .B2 (n_14));
AOI21_X1 i_24 (.ZN (p_0[13]), .A (n_15), .B1 (p_1[13]), .B2 (n_16));
AOI21_X1 i_23 (.ZN (p_0[12]), .A (n_17), .B1 (p_1[12]), .B2 (n_144));
NOR2_X1 i_22 (.ZN (n_11), .A1 (p_1[8]), .A2 (n_119));
INV_X1 i_21 (.ZN (n_10), .A (n_11));
NOR2_X1 i_20 (.ZN (n_9), .A1 (p_1[9]), .A2 (n_10));
INV_X1 i_19 (.ZN (n_8), .A (n_9));
NOR2_X1 i_18 (.ZN (n_7), .A1 (n_119), .A2 (n_118));
INV_X1 i_17 (.ZN (n_6), .A (n_7));
AOI21_X1 i_16 (.ZN (p_0[11]), .A (n_117), .B1 (p_1[11]), .B2 (n_6));
AOI21_X1 i_15 (.ZN (p_0[10]), .A (n_7), .B1 (p_1[10]), .B2 (n_8));
AOI21_X1 i_14 (.ZN (p_0[9]), .A (n_9), .B1 (p_1[9]), .B2 (n_10));
AOI21_X1 i_13 (.ZN (p_0[8]), .A (n_11), .B1 (p_1[8]), .B2 (n_119));
NOR2_X1 i_12 (.ZN (n_5), .A1 (p_1[4]), .A2 (n_122));
INV_X1 i_11 (.ZN (n_4), .A (n_5));
NOR2_X1 i_10 (.ZN (n_3), .A1 (p_1[5]), .A2 (n_4));
INV_X1 i_9 (.ZN (n_2), .A (n_3));
NOR2_X1 i_8 (.ZN (n_1), .A1 (n_122), .A2 (n_121));
INV_X1 i_7 (.ZN (n_0), .A (n_1));
AOI21_X1 i_6 (.ZN (p_0[7]), .A (n_120), .B1 (p_1[7]), .B2 (n_0));
AOI21_X1 i_5 (.ZN (p_0[6]), .A (n_1), .B1 (p_1[6]), .B2 (n_2));
AOI21_X1 i_4 (.ZN (p_0[5]), .A (n_3), .B1 (p_1[5]), .B2 (n_4));
AOI21_X1 i_3 (.ZN (p_0[4]), .A (n_5), .B1 (p_1[4]), .B2 (n_122));
AOI21_X1 i_2 (.ZN (p_0[3]), .A (n_123), .B1 (p_1[3]), .B2 (n_124));
AOI21_X1 i_1 (.ZN (p_0[2]), .A (n_125), .B1 (p_1[2]), .B2 (n_126));
AOI21_X1 i_0 (.ZN (p_0[1]), .A (n_127), .B1 (p_1[1]), .B2 (p_1[0]));

endmodule //datapath__0_72

module datapath__0_67 (p_0, b);

output [31:0] p_0;
input [31:0] b;
wire n_62;
wire n_60;
wire n_61;
wire n_58;
wire n_59;
wire n_5;
wire n_57;
wire n_1;
wire n_56;
wire n_7;
wire n_54;
wire n_53;
wire n_13;
wire n_51;
wire n_50;
wire n_21;
wire n_19;
wire n_20;
wire n_45;
wire n_18;
wire n_48;
wire n_46;
wire n_25;
wire n_44;
wire n_27;
wire n_24;
wire n_43;
wire n_26;
wire n_41;
wire n_42;
wire n_29;
wire n_40;
wire n_28;
wire n_30;
wire n_63;
wire n_32;
wire n_39;
wire n_31;
wire n_47;
wire n_34;
wire n_38;
wire n_36;
wire n_33;
wire n_37;
wire n_35;
wire n_0;
wire n_68;
wire n_49;
wire n_4;
wire n_11;
wire n_6;
wire n_10;
wire n_79;
wire n_12;
wire n_52;
wire n_16;
wire n_17;
wire n_55;
wire n_76;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_70;
wire n_69;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_77;
wire n_78;
wire n_80;
wire n_81;
wire n_85;
wire n_84;
wire n_83;
wire n_82;


INV_X1 i_116 (.ZN (n_85), .A (b[3]));
INV_X1 i_115 (.ZN (n_84), .A (b[2]));
INV_X1 i_114 (.ZN (n_83), .A (b[1]));
INV_X1 i_113 (.ZN (n_82), .A (b[0]));
NAND2_X1 i_112 (.ZN (n_61), .A1 (n_83), .A2 (n_82));
INV_X1 i_111 (.ZN (n_62), .A (n_61));
NAND2_X1 i_110 (.ZN (n_59), .A1 (n_62), .A2 (n_84));
INV_X1 i_109 (.ZN (n_60), .A (n_59));
NAND2_X1 i_108 (.ZN (n_57), .A1 (n_60), .A2 (n_85));
INV_X1 i_107 (.ZN (n_58), .A (n_57));
OR3_X1 i_106 (.ZN (n_56), .A1 (b[6]), .A2 (b[5]), .A3 (b[4]));
OR2_X1 i_105 (.ZN (n_81), .A1 (n_56), .A2 (b[7]));
INV_X1 i_104 (.ZN (n_80), .A (n_81));
NAND2_X1 i_103 (.ZN (n_54), .A1 (n_80), .A2 (n_58));
INV_X1 i_102 (.ZN (n_79), .A (n_54));
OR3_X1 i_101 (.ZN (n_53), .A1 (b[10]), .A2 (b[9]), .A3 (b[8]));
OR2_X1 i_100 (.ZN (n_78), .A1 (n_53), .A2 (b[11]));
INV_X1 i_99 (.ZN (n_77), .A (n_78));
NAND2_X1 i_98 (.ZN (n_51), .A1 (n_79), .A2 (n_77));
INV_X1 i_97 (.ZN (n_76), .A (n_51));
OR3_X1 i_96 (.ZN (n_50), .A1 (b[14]), .A2 (b[13]), .A3 (b[12]));
OR2_X1 i_95 (.ZN (n_75), .A1 (n_50), .A2 (b[15]));
INV_X1 i_93 (.ZN (n_74), .A (n_75));
NAND2_X1 i_92 (.ZN (n_48), .A1 (n_76), .A2 (n_74));
XNOR2_X1 i_91 (.ZN (n_73), .A (n_48), .B (b[16]));
INV_X1 i_90 (.ZN (p_0[16]), .A (n_73));
INV_X1 i_89 (.ZN (n_72), .A (n_13));
INV_X1 i_88 (.ZN (n_71), .A (n_48));
AOI21_X1 i_87 (.ZN (p_0[15]), .A (n_71), .B1 (n_72), .B2 (b[15]));
INV_X1 i_86 (.ZN (n_70), .A (b[13]));
INV_X1 i_85 (.ZN (n_69), .A (b[12]));
NAND3_X1 i_84 (.ZN (n_68), .A1 (n_76), .A2 (n_70), .A3 (n_69));
OAI21_X1 i_83 (.ZN (n_67), .A (b[13]), .B1 (n_51), .B2 (b[12]));
NAND2_X1 i_82 (.ZN (n_66), .A1 (n_67), .A2 (n_68));
INV_X1 i_81 (.ZN (p_0[13]), .A (n_66));
XNOR2_X1 i_80 (.ZN (n_65), .A (n_51), .B (b[12]));
INV_X1 i_79 (.ZN (p_0[12]), .A (n_65));
INV_X1 i_42 (.ZN (n_64), .A (n_7));
AOI21_X1 i_33 (.ZN (p_0[11]), .A (n_76), .B1 (n_64), .B2 (b[11]));
INV_X1 i_32 (.ZN (n_55), .A (b[9]));
INV_X1 i_31 (.ZN (n_52), .A (b[8]));
NAND3_X1 i_30 (.ZN (n_49), .A1 (n_79), .A2 (n_55), .A3 (n_52));
OAI21_X1 i_27 (.ZN (n_17), .A (b[9]), .B1 (n_54), .B2 (b[8]));
NAND2_X1 i_26 (.ZN (n_16), .A1 (n_17), .A2 (n_49));
INV_X1 i_24 (.ZN (p_0[9]), .A (n_16));
XNOR2_X1 i_23 (.ZN (p_0[8]), .A (n_54), .B (n_52));
INV_X1 i_22 (.ZN (n_12), .A (n_1));
AOI21_X1 i_21 (.ZN (p_0[7]), .A (n_79), .B1 (n_12), .B2 (b[7]));
INV_X1 i_20 (.ZN (n_11), .A (b[5]));
INV_X1 i_17 (.ZN (n_10), .A (b[4]));
NAND2_X1 i_16 (.ZN (n_6), .A1 (n_58), .A2 (n_10));
XNOR2_X1 i_14 (.ZN (p_0[5]), .A (n_6), .B (n_11));
INV_X1 i_13 (.ZN (n_5), .A (n_6));
NAND2_X1 i_12 (.ZN (n_4), .A1 (n_5), .A2 (n_11));
OR2_X1 i_6 (.ZN (n_0), .A1 (n_48), .A2 (b[16]));
INV_X1 i_94 (.ZN (n_63), .A (b[25]));
OR3_X1 i_78 (.ZN (n_47), .A1 (b[26]), .A2 (b[25]), .A3 (b[24]));
OR3_X1 i_77 (.ZN (n_46), .A1 (b[18]), .A2 (b[16]), .A3 (b[17]));
NOR3_X1 i_76 (.ZN (n_45), .A1 (b[19]), .A2 (n_46), .A3 (n_48));
INV_X1 i_75 (.ZN (n_44), .A (n_45));
NOR4_X1 i_74 (.ZN (n_43), .A1 (b[22]), .A2 (b[21]), .A3 (b[20]), .A4 (n_44));
INV_X1 i_73 (.ZN (n_42), .A (n_43));
NOR2_X1 i_72 (.ZN (n_41), .A1 (b[23]), .A2 (n_42));
INV_X1 i_71 (.ZN (n_40), .A (n_41));
NOR3_X1 i_70 (.ZN (n_39), .A1 (b[27]), .A2 (n_47), .A3 (n_40));
INV_X1 i_69 (.ZN (n_38), .A (n_39));
NOR4_X1 i_68 (.ZN (n_37), .A1 (b[29]), .A2 (b[28]), .A3 (b[30]), .A4 (n_38));
XNOR2_X1 i_67 (.ZN (p_0[31]), .A (b[31]), .B (n_37));
NOR3_X1 i_66 (.ZN (n_36), .A1 (b[29]), .A2 (b[28]), .A3 (n_38));
INV_X1 i_65 (.ZN (n_35), .A (n_36));
AOI21_X1 i_64 (.ZN (p_0[30]), .A (n_37), .B1 (b[30]), .B2 (n_35));
NOR2_X1 i_63 (.ZN (n_34), .A1 (b[28]), .A2 (n_38));
INV_X1 i_62 (.ZN (n_33), .A (n_34));
AOI21_X1 i_61 (.ZN (p_0[29]), .A (n_36), .B1 (b[29]), .B2 (n_33));
AOI21_X1 i_60 (.ZN (p_0[28]), .A (n_34), .B1 (b[28]), .B2 (n_38));
NOR2_X1 i_59 (.ZN (n_32), .A1 (n_47), .A2 (n_40));
INV_X1 i_58 (.ZN (n_31), .A (n_32));
AOI21_X1 i_57 (.ZN (p_0[27]), .A (n_39), .B1 (b[27]), .B2 (n_31));
OR3_X1 i_56 (.ZN (n_30), .A1 (b[25]), .A2 (b[24]), .A3 (n_40));
AOI21_X1 i_55 (.ZN (p_0[26]), .A (n_32), .B1 (b[26]), .B2 (n_30));
NOR2_X1 i_54 (.ZN (n_29), .A1 (b[24]), .A2 (n_40));
OAI21_X1 i_53 (.ZN (n_28), .A (n_30), .B1 (n_63), .B2 (n_29));
INV_X1 i_52 (.ZN (p_0[25]), .A (n_28));
AOI21_X1 i_51 (.ZN (p_0[24]), .A (n_29), .B1 (b[24]), .B2 (n_40));
AOI21_X1 i_50 (.ZN (p_0[23]), .A (n_41), .B1 (b[23]), .B2 (n_42));
NOR3_X1 i_49 (.ZN (n_27), .A1 (b[21]), .A2 (b[20]), .A3 (n_44));
INV_X1 i_48 (.ZN (n_26), .A (n_27));
AOI21_X1 i_47 (.ZN (p_0[22]), .A (n_43), .B1 (b[22]), .B2 (n_26));
NOR2_X1 i_46 (.ZN (n_25), .A1 (b[20]), .A2 (n_44));
INV_X1 i_45 (.ZN (n_24), .A (n_25));
AOI21_X1 i_44 (.ZN (p_0[21]), .A (n_27), .B1 (b[21]), .B2 (n_24));
AOI21_X1 i_43 (.ZN (p_0[20]), .A (n_25), .B1 (b[20]), .B2 (n_44));
NOR2_X1 i_40 (.ZN (n_21), .A1 (b[17]), .A2 (n_0));
INV_X1 i_39 (.ZN (n_20), .A (n_21));
NOR2_X1 i_38 (.ZN (n_19), .A1 (n_48), .A2 (n_46));
INV_X1 i_37 (.ZN (n_18), .A (n_19));
AOI21_X1 i_36 (.ZN (p_0[19]), .A (n_45), .B1 (b[19]), .B2 (n_18));
AOI21_X1 i_35 (.ZN (p_0[18]), .A (n_19), .B1 (b[18]), .B2 (n_20));
AOI21_X1 i_34 (.ZN (p_0[17]), .A (n_21), .B1 (b[17]), .B2 (n_0));
NOR2_X1 i_28 (.ZN (n_13), .A1 (n_51), .A2 (n_50));
AOI21_X1 i_25 (.ZN (p_0[14]), .A (n_13), .B1 (b[14]), .B2 (n_68));
NOR2_X1 i_18 (.ZN (n_7), .A1 (n_54), .A2 (n_53));
AOI21_X1 i_15 (.ZN (p_0[10]), .A (n_7), .B1 (b[10]), .B2 (n_49));
NOR2_X1 i_8 (.ZN (n_1), .A1 (n_57), .A2 (n_56));
AOI21_X1 i_5 (.ZN (p_0[6]), .A (n_1), .B1 (b[6]), .B2 (n_4));
AOI21_X1 i_3 (.ZN (p_0[4]), .A (n_5), .B1 (b[4]), .B2 (n_57));
AOI21_X1 i_2 (.ZN (p_0[3]), .A (n_58), .B1 (b[3]), .B2 (n_59));
AOI21_X1 i_1 (.ZN (p_0[2]), .A (n_60), .B1 (b[2]), .B2 (n_61));
AOI21_X1 i_0 (.ZN (p_0[1]), .A (n_62), .B1 (b[1]), .B2 (b[0]));

endmodule //datapath__0_67

module datapath__0_66 (multiplicand, A, p_0);

output [31:0] p_0;
input [31:0] A;
input [31:0] multiplicand;
wire n_0;
wire n_154;
wire n_1;
wire n_153;
wire n_152;
wire n_2;
wire n_157;
wire n_151;
wire n_3;
wire n_158;
wire n_164;
wire n_161;
wire n_149;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_146;
wire n_137;
wire n_11;
wire n_5;
wire n_147;
wire n_141;
wire n_8;
wire n_144;
wire n_142;
wire n_148;
wire n_139;
wire n_135;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_132;
wire n_123;
wire n_19;
wire n_13;
wire n_133;
wire n_127;
wire n_16;
wire n_130;
wire n_128;
wire n_134;
wire n_125;
wire n_121;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_118;
wire n_109;
wire n_27;
wire n_21;
wire n_119;
wire n_113;
wire n_24;
wire n_116;
wire n_114;
wire n_120;
wire n_111;
wire n_107;
wire n_34;
wire n_33;
wire n_30;
wire n_31;
wire n_28;
wire n_104;
wire n_95;
wire n_35;
wire n_29;
wire n_105;
wire n_99;
wire n_32;
wire n_102;
wire n_100;
wire n_106;
wire n_97;
wire n_93;
wire n_42;
wire n_41;
wire n_38;
wire n_39;
wire n_36;
wire n_82;
wire n_72;
wire n_43;
wire n_37;
wire n_81;
wire n_84;
wire n_74;
wire n_40;
wire n_83;
wire n_79;
wire n_76;
wire n_86;
wire n_51;
wire n_50;
wire n_69;
wire n_64;
wire n_63;
wire n_62;
wire n_58;
wire n_55;
wire n_54;
wire n_160;
wire n_166;
wire n_163;
wire n_61;
wire n_60;
wire n_57;
wire n_56;
wire n_59;
wire n_159;
wire n_67;
wire n_65;
wire n_70;
wire n_77;
wire n_165;
wire n_162;
wire n_92;
wire n_66;
wire n_89;
wire n_68;
wire n_87;
wire n_71;
wire n_75;
wire n_78;
wire n_88;
wire n_90;
wire n_96;
wire n_94;
wire n_103;
wire n_98;
wire n_101;
wire n_108;
wire n_112;
wire n_115;
wire n_110;
wire n_117;
wire n_122;
wire n_126;
wire n_129;
wire n_124;
wire n_131;
wire n_136;
wire n_140;
wire n_143;
wire n_138;
wire n_145;
wire n_150;
wire n_156;
wire n_155;
wire n_179;
wire n_184;
wire n_169;
wire n_171;
wire n_44;
wire n_45;
wire n_53;
wire n_183;
wire n_168;
wire n_46;
wire n_48;
wire n_47;
wire n_167;
wire n_49;
wire n_52;
wire n_185;
wire n_187;
wire n_186;
wire n_73;
wire n_85;
wire n_80;
wire n_189;
wire n_91;
wire n_188;
wire n_182;
wire n_175;
wire n_170;
wire n_173;
wire n_172;
wire n_176;
wire n_174;
wire n_178;
wire n_177;
wire n_181;
wire n_180;


OAI22_X1 i_221 (.ZN (n_189), .A1 (n_165), .A2 (n_162), .B1 (multiplicand[27]), .B2 (A[27]));
INV_X1 i_220 (.ZN (n_188), .A (n_189));
NAND2_X1 i_219 (.ZN (n_66), .A1 (multiplicand[26]), .A2 (A[26]));
INV_X1 i_218 (.ZN (n_187), .A (multiplicand[25]));
INV_X1 i_217 (.ZN (n_186), .A (A[25]));
NOR2_X1 i_216 (.ZN (n_185), .A1 (multiplicand[26]), .A2 (A[26]));
AOI21_X1 i_215 (.ZN (n_184), .A (n_185), .B1 (n_187), .B2 (n_186));
NAND2_X1 i_214 (.ZN (n_183), .A1 (multiplicand[25]), .A2 (A[25]));
NAND2_X1 i_213 (.ZN (n_69), .A1 (multiplicand[24]), .A2 (A[24]));
INV_X1 i_212 (.ZN (n_182), .A (n_69));
INV_X1 i_211 (.ZN (n_181), .A (multiplicand[24]));
INV_X1 i_210 (.ZN (n_180), .A (A[24]));
NAND2_X1 i_209 (.ZN (n_179), .A1 (n_181), .A2 (n_180));
INV_X1 i_208 (.ZN (n_178), .A (n_79));
INV_X1 i_207 (.ZN (n_83), .A (n_84));
NOR2_X1 i_206 (.ZN (n_82), .A1 (multiplicand[22]), .A2 (A[22]));
INV_X1 i_205 (.ZN (n_81), .A (n_82));
NAND2_X1 i_204 (.ZN (n_177), .A1 (n_81), .A2 (n_83));
INV_X1 i_203 (.ZN (n_176), .A (n_177));
OAI211_X1 i_202 (.ZN (n_78), .A (n_178), .B (n_176), .C1 (multiplicand[23]), .C2 (A[23]));
NOR4_X1 i_201 (.ZN (n_93), .A1 (n_101), .A2 (n_98), .A3 (n_97), .A4 (n_94));
OR2_X1 i_200 (.ZN (n_175), .A1 (n_78), .A2 (n_93));
NOR2_X1 i_199 (.ZN (n_86), .A1 (multiplicand[23]), .A2 (A[23]));
NAND2_X1 i_125 (.ZN (n_76), .A1 (multiplicand[20]), .A2 (A[20]));
NAND2_X1 i_123 (.ZN (n_75), .A1 (multiplicand[21]), .A2 (A[21]));
NAND2_X1 i_122 (.ZN (n_174), .A1 (n_75), .A2 (n_76));
OAI211_X1 i_120 (.ZN (n_173), .A (n_176), .B (n_174), .C1 (multiplicand[23]), .C2 (A[23]));
NAND2_X1 i_118 (.ZN (n_172), .A1 (multiplicand[23]), .A2 (A[23]));
NAND2_X1 i_117 (.ZN (n_171), .A1 (multiplicand[22]), .A2 (A[22]));
OAI211_X1 i_115 (.ZN (n_170), .A (n_173), .B (n_172), .C1 (n_86), .C2 (n_171));
INV_X1 i_114 (.ZN (n_71), .A (n_170));
NAND2_X1 i_113 (.ZN (n_169), .A1 (n_71), .A2 (n_175));
AOI21_X1 i_112 (.ZN (n_168), .A (n_182), .B1 (n_169), .B2 (n_179));
NAND2_X1 i_110 (.ZN (n_167), .A1 (n_183), .A2 (n_168));
NAND2_X1 i_108 (.ZN (n_91), .A1 (n_184), .A2 (n_167));
NAND3_X1 i_107 (.ZN (n_85), .A1 (n_91), .A2 (n_188), .A3 (n_66));
NAND2_X1 i_105 (.ZN (n_80), .A1 (n_91), .A2 (n_66));
NAND2_X1 i_104 (.ZN (n_73), .A1 (n_80), .A2 (n_189));
NAND2_X1 i_103 (.ZN (p_0[27]), .A1 (n_73), .A2 (n_85));
NAND2_X1 i_101 (.ZN (n_53), .A1 (n_187), .A2 (n_186));
INV_X1 i_98 (.ZN (n_52), .A (n_185));
NAND2_X1 i_81 (.ZN (n_49), .A1 (n_52), .A2 (n_66));
AOI21_X1 i_80 (.ZN (n_48), .A (n_49), .B1 (n_167), .B2 (n_53));
NAND3_X1 i_79 (.ZN (n_47), .A1 (n_167), .A2 (n_53), .A3 (n_49));
INV_X1 i_77 (.ZN (n_46), .A (n_47));
OR2_X1 i_76 (.ZN (p_0[26]), .A1 (n_46), .A2 (n_48));
INV_X1 i_75 (.ZN (n_45), .A (n_168));
NAND2_X1 i_74 (.ZN (n_44), .A1 (n_53), .A2 (n_183));
XNOR2_X1 i_73 (.ZN (p_0[25]), .A (n_44), .B (n_45));
INV_X1 i_72 (.ZN (n_72), .A (n_171));
INV_X1 i_71 (.ZN (n_51), .A (n_169));
INV_X1 i_70 (.ZN (n_90), .A (n_184));
INV_X1 i_69 (.ZN (n_88), .A (n_179));
INV_X1 i_198 (.ZN (n_166), .A (multiplicand[30]));
INV_X1 i_197 (.ZN (n_165), .A (multiplicand[27]));
INV_X1 i_196 (.ZN (n_164), .A (multiplicand[3]));
INV_X1 i_195 (.ZN (n_163), .A (A[31]));
INV_X1 i_194 (.ZN (n_162), .A (A[27]));
INV_X1 i_193 (.ZN (n_161), .A (A[3]));
NAND2_X1 i_192 (.ZN (n_160), .A1 (n_166), .A2 (n_163));
NOR2_X1 i_191 (.ZN (n_159), .A1 (multiplicand[28]), .A2 (A[28]));
NAND2_X1 i_190 (.ZN (n_158), .A1 (n_164), .A2 (n_161));
NAND2_X1 i_189 (.ZN (n_157), .A1 (multiplicand[2]), .A2 (A[2]));
INV_X1 i_188 (.ZN (n_156), .A (n_157));
NOR2_X1 i_187 (.ZN (n_155), .A1 (multiplicand[1]), .A2 (A[1]));
NAND2_X1 i_186 (.ZN (n_154), .A1 (multiplicand[0]), .A2 (A[0]));
NAND2_X1 i_185 (.ZN (n_153), .A1 (multiplicand[1]), .A2 (A[1]));
AOI21_X1 i_184 (.ZN (n_152), .A (n_155), .B1 (n_154), .B2 (n_153));
OAI22_X1 i_183 (.ZN (n_151), .A1 (multiplicand[2]), .A2 (A[2]), .B1 (n_156), .B2 (n_152));
OAI21_X1 i_182 (.ZN (n_150), .A (n_151), .B1 (n_164), .B2 (n_161));
NAND2_X1 i_181 (.ZN (n_149), .A1 (n_158), .A2 (n_150));
NOR2_X1 i_180 (.ZN (n_148), .A1 (multiplicand[7]), .A2 (A[7]));
NOR2_X1 i_179 (.ZN (n_147), .A1 (multiplicand[5]), .A2 (A[5]));
NOR2_X1 i_178 (.ZN (n_146), .A1 (multiplicand[6]), .A2 (A[6]));
OR3_X1 i_177 (.ZN (n_145), .A1 (n_148), .A2 (n_146), .A3 (n_147));
NOR2_X1 i_176 (.ZN (n_144), .A1 (multiplicand[4]), .A2 (A[4]));
NOR3_X1 i_175 (.ZN (n_143), .A1 (n_145), .A2 (n_144), .A3 (n_149));
NAND2_X1 i_174 (.ZN (n_142), .A1 (multiplicand[4]), .A2 (A[4]));
NAND2_X1 i_173 (.ZN (n_141), .A1 (multiplicand[5]), .A2 (A[5]));
AOI21_X1 i_172 (.ZN (n_140), .A (n_145), .B1 (n_142), .B2 (n_141));
AND2_X1 i_171 (.ZN (n_139), .A1 (multiplicand[7]), .A2 (A[7]));
NAND2_X1 i_170 (.ZN (n_138), .A1 (multiplicand[6]), .A2 (A[6]));
INV_X1 i_169 (.ZN (n_137), .A (n_138));
NOR2_X1 i_168 (.ZN (n_136), .A1 (n_148), .A2 (n_138));
NOR4_X1 i_167 (.ZN (n_135), .A1 (n_139), .A2 (n_136), .A3 (n_140), .A4 (n_143));
NOR2_X1 i_166 (.ZN (n_134), .A1 (multiplicand[11]), .A2 (A[11]));
NOR2_X1 i_165 (.ZN (n_133), .A1 (multiplicand[9]), .A2 (A[9]));
NOR2_X1 i_164 (.ZN (n_132), .A1 (multiplicand[10]), .A2 (A[10]));
OR3_X1 i_163 (.ZN (n_131), .A1 (n_134), .A2 (n_132), .A3 (n_133));
NOR2_X1 i_162 (.ZN (n_130), .A1 (multiplicand[8]), .A2 (A[8]));
NOR3_X1 i_161 (.ZN (n_129), .A1 (n_131), .A2 (n_130), .A3 (n_135));
NAND2_X1 i_160 (.ZN (n_128), .A1 (multiplicand[8]), .A2 (A[8]));
NAND2_X1 i_159 (.ZN (n_127), .A1 (multiplicand[9]), .A2 (A[9]));
AOI21_X1 i_158 (.ZN (n_126), .A (n_131), .B1 (n_128), .B2 (n_127));
AND2_X1 i_157 (.ZN (n_125), .A1 (multiplicand[11]), .A2 (A[11]));
NAND2_X1 i_156 (.ZN (n_124), .A1 (multiplicand[10]), .A2 (A[10]));
INV_X1 i_155 (.ZN (n_123), .A (n_124));
NOR2_X1 i_154 (.ZN (n_122), .A1 (n_134), .A2 (n_124));
NOR4_X1 i_153 (.ZN (n_121), .A1 (n_125), .A2 (n_122), .A3 (n_126), .A4 (n_129));
NOR2_X1 i_152 (.ZN (n_120), .A1 (multiplicand[15]), .A2 (A[15]));
NOR2_X1 i_151 (.ZN (n_119), .A1 (multiplicand[13]), .A2 (A[13]));
NOR2_X1 i_150 (.ZN (n_118), .A1 (multiplicand[14]), .A2 (A[14]));
OR3_X1 i_149 (.ZN (n_117), .A1 (n_120), .A2 (n_118), .A3 (n_119));
NOR2_X1 i_148 (.ZN (n_116), .A1 (multiplicand[12]), .A2 (A[12]));
NOR3_X2 i_147 (.ZN (n_115), .A1 (n_117), .A2 (n_116), .A3 (n_121));
NAND2_X1 i_146 (.ZN (n_114), .A1 (multiplicand[12]), .A2 (A[12]));
NAND2_X1 i_145 (.ZN (n_113), .A1 (multiplicand[13]), .A2 (A[13]));
AOI21_X1 i_144 (.ZN (n_112), .A (n_117), .B1 (n_114), .B2 (n_113));
AND2_X1 i_143 (.ZN (n_111), .A1 (multiplicand[15]), .A2 (A[15]));
NAND2_X1 i_142 (.ZN (n_110), .A1 (multiplicand[14]), .A2 (A[14]));
INV_X1 i_141 (.ZN (n_109), .A (n_110));
NOR2_X1 i_140 (.ZN (n_108), .A1 (n_120), .A2 (n_110));
NOR4_X1 i_139 (.ZN (n_107), .A1 (n_111), .A2 (n_108), .A3 (n_112), .A4 (n_115));
NOR2_X1 i_138 (.ZN (n_106), .A1 (multiplicand[19]), .A2 (A[19]));
NOR2_X1 i_137 (.ZN (n_105), .A1 (multiplicand[17]), .A2 (A[17]));
NOR2_X1 i_136 (.ZN (n_104), .A1 (multiplicand[18]), .A2 (A[18]));
OR3_X1 i_135 (.ZN (n_103), .A1 (n_106), .A2 (n_104), .A3 (n_105));
NOR2_X1 i_134 (.ZN (n_102), .A1 (multiplicand[16]), .A2 (A[16]));
NOR3_X1 i_133 (.ZN (n_101), .A1 (n_103), .A2 (n_102), .A3 (n_107));
NAND2_X1 i_132 (.ZN (n_100), .A1 (multiplicand[16]), .A2 (A[16]));
NAND2_X1 i_131 (.ZN (n_99), .A1 (multiplicand[17]), .A2 (A[17]));
AOI21_X1 i_130 (.ZN (n_98), .A (n_103), .B1 (n_100), .B2 (n_99));
AND2_X1 i_129 (.ZN (n_97), .A1 (multiplicand[19]), .A2 (A[19]));
NAND2_X1 i_128 (.ZN (n_96), .A1 (multiplicand[18]), .A2 (A[18]));
INV_X1 i_127 (.ZN (n_95), .A (n_96));
NOR2_X1 i_126 (.ZN (n_94), .A1 (n_106), .A2 (n_96));
NOR2_X1 i_124 (.ZN (n_92), .A1 (multiplicand[27]), .A2 (A[27]));
OR2_X1 i_121 (.ZN (n_89), .A1 (n_92), .A2 (n_90));
OR2_X1 i_119 (.ZN (n_87), .A1 (n_89), .A2 (n_88));
NOR2_X1 i_116 (.ZN (n_84), .A1 (multiplicand[21]), .A2 (A[21]));
NOR2_X1 i_111 (.ZN (n_79), .A1 (multiplicand[20]), .A2 (A[20]));
NOR3_X1 i_109 (.ZN (n_77), .A1 (n_87), .A2 (n_78), .A3 (n_93));
INV_X1 i_106 (.ZN (n_74), .A (n_75));
NOR2_X1 i_102 (.ZN (n_70), .A1 (n_87), .A2 (n_71));
NAND2_X1 i_100 (.ZN (n_68), .A1 (multiplicand[25]), .A2 (A[25]));
AOI21_X1 i_99 (.ZN (n_67), .A (n_89), .B1 (n_69), .B2 (n_68));
OAI22_X1 i_97 (.ZN (n_65), .A1 (n_165), .A2 (n_162), .B1 (n_92), .B2 (n_66));
NOR4_X1 i_96 (.ZN (n_64), .A1 (n_67), .A2 (n_65), .A3 (n_70), .A4 (n_77));
AOI21_X1 i_95 (.ZN (n_63), .A (n_159), .B1 (multiplicand[28]), .B2 (A[28]));
AOI21_X1 i_94 (.ZN (n_62), .A (n_159), .B1 (n_64), .B2 (n_63));
AOI21_X1 i_93 (.ZN (n_61), .A (n_62), .B1 (multiplicand[29]), .B2 (A[29]));
NOR2_X1 i_92 (.ZN (n_60), .A1 (multiplicand[29]), .A2 (A[29]));
OAI22_X1 i_91 (.ZN (n_59), .A1 (n_166), .A2 (n_163), .B1 (multiplicand[29]), .B2 (A[29]));
AOI21_X1 i_90 (.ZN (n_58), .A (n_60), .B1 (multiplicand[29]), .B2 (A[29]));
OAI21_X1 i_89 (.ZN (n_57), .A (n_160), .B1 (n_61), .B2 (n_59));
XNOR2_X1 i_88 (.ZN (n_56), .A (multiplicand[31]), .B (multiplicand[30]));
XOR2_X1 i_87 (.Z (p_0[31]), .A (n_57), .B (n_56));
NOR2_X1 i_86 (.ZN (n_55), .A1 (n_61), .A2 (n_60));
OAI21_X1 i_85 (.ZN (n_54), .A (n_160), .B1 (n_166), .B2 (n_163));
XNOR2_X1 i_84 (.ZN (p_0[30]), .A (n_55), .B (n_54));
XOR2_X1 i_83 (.Z (p_0[29]), .A (n_62), .B (n_58));
XNOR2_X1 i_82 (.ZN (p_0[28]), .A (n_64), .B (n_63));
OAI21_X1 i_78 (.ZN (n_50), .A (n_69), .B1 (multiplicand[24]), .B2 (A[24]));
XOR2_X1 i_68 (.Z (p_0[24]), .A (n_51), .B (n_50));
AOI21_X1 i_67 (.ZN (n_43), .A (n_86), .B1 (multiplicand[23]), .B2 (A[23]));
OAI21_X1 i_66 (.ZN (n_42), .A (n_76), .B1 (multiplicand[20]), .B2 (A[20]));
AOI21_X1 i_65 (.ZN (n_41), .A (n_79), .B1 (n_93), .B2 (n_76));
OAI21_X1 i_64 (.ZN (n_40), .A (n_83), .B1 (n_74), .B2 (n_41));
INV_X1 i_63 (.ZN (n_39), .A (n_40));
NOR2_X1 i_62 (.ZN (n_38), .A1 (n_84), .A2 (n_74));
OAI21_X1 i_61 (.ZN (n_37), .A (n_81), .B1 (n_72), .B2 (n_39));
XNOR2_X1 i_60 (.ZN (p_0[23]), .A (n_43), .B (n_37));
NOR2_X1 i_59 (.ZN (n_36), .A1 (n_82), .A2 (n_72));
XOR2_X1 i_58 (.Z (p_0[22]), .A (n_39), .B (n_36));
XOR2_X1 i_57 (.Z (p_0[21]), .A (n_41), .B (n_38));
XOR2_X1 i_56 (.Z (p_0[20]), .A (n_93), .B (n_42));
NOR2_X1 i_55 (.ZN (n_35), .A1 (n_106), .A2 (n_97));
OAI21_X1 i_54 (.ZN (n_34), .A (n_100), .B1 (multiplicand[16]), .B2 (A[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_102), .B1 (n_107), .B2 (n_100));
INV_X1 i_52 (.ZN (n_32), .A (n_33));
AOI21_X1 i_51 (.ZN (n_31), .A (n_105), .B1 (n_99), .B2 (n_32));
AOI21_X1 i_50 (.ZN (n_30), .A (n_105), .B1 (multiplicand[17]), .B2 (A[17]));
OAI22_X1 i_49 (.ZN (n_29), .A1 (multiplicand[18]), .A2 (A[18]), .B1 (n_95), .B2 (n_31));
XNOR2_X1 i_48 (.ZN (p_0[19]), .A (n_35), .B (n_29));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_104), .A2 (n_95));
XOR2_X1 i_46 (.Z (p_0[18]), .A (n_31), .B (n_28));
XOR2_X1 i_45 (.Z (p_0[17]), .A (n_33), .B (n_30));
XOR2_X1 i_44 (.Z (p_0[16]), .A (n_107), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_120), .A2 (n_111));
OAI21_X1 i_42 (.ZN (n_26), .A (n_114), .B1 (multiplicand[12]), .B2 (A[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_116), .B1 (n_121), .B2 (n_114));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_119), .B1 (n_113), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_119), .B1 (multiplicand[13]), .B2 (A[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (multiplicand[14]), .A2 (A[14]), .B1 (n_109), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (p_0[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_118), .A2 (n_109));
XOR2_X1 i_34 (.Z (p_0[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (p_0[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (p_0[12]), .A (n_121), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_134), .A2 (n_125));
AOI21_X1 i_30 (.ZN (n_18), .A (n_130), .B1 (multiplicand[8]), .B2 (A[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_130), .B1 (n_135), .B2 (n_128));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_133), .B1 (n_127), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_133), .B1 (multiplicand[9]), .B2 (A[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (multiplicand[10]), .A2 (A[10]), .B1 (n_123), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (p_0[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_132), .A2 (n_123));
XOR2_X1 i_22 (.Z (p_0[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (p_0[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (p_0[8]), .A (n_135), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_148), .A2 (n_139));
OAI21_X1 i_18 (.ZN (n_10), .A (n_142), .B1 (multiplicand[4]), .B2 (A[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_144), .B1 (n_149), .B2 (n_142));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_147), .B1 (n_141), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_147), .B1 (multiplicand[5]), .B2 (A[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (multiplicand[6]), .A2 (A[6]), .B1 (n_137), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (p_0[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_146), .A2 (n_137));
XOR2_X1 i_10 (.Z (p_0[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (p_0[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (p_0[4]), .A (n_149), .B (n_10));
OAI21_X1 i_7 (.ZN (n_3), .A (n_158), .B1 (n_164), .B2 (n_161));
XOR2_X1 i_6 (.Z (p_0[3]), .A (n_151), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_157), .B1 (multiplicand[2]), .B2 (A[2]));
XNOR2_X1 i_4 (.ZN (p_0[2]), .A (n_152), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_153), .B1 (multiplicand[1]), .B2 (A[1]));
XOR2_X1 i_2 (.Z (p_0[1]), .A (n_154), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_154), .B1 (multiplicand[0]), .B2 (A[0]));
INV_X1 i_0 (.ZN (p_0[0]), .A (n_0));

endmodule //datapath__0_66

module datapath__0_65 (A, p_0, multiplicand);

output [31:0] p_0;
input [31:0] A;
input [31:0] multiplicand;
wire n_102;
wire n_123;
wire n_101;
wire n_0;
wire n_111;
wire n_104;
wire n_3;
wire n_1;
wire n_109;
wire n_100;
wire n_4;
wire n_2;
wire n_110;
wire n_124;
wire n_108;
wire n_126;
wire n_97;
wire n_5;
wire n_112;
wire n_96;
wire n_11;
wire n_6;
wire n_115;
wire n_128;
wire n_9;
wire n_7;
wire n_116;
wire n_129;
wire n_12;
wire n_8;
wire n_93;
wire n_10;
wire n_95;
wire n_127;
wire n_114;
wire n_130;
wire n_28;
wire n_13;
wire n_118;
wire n_229;
wire n_18;
wire n_14;
wire n_161;
wire n_227;
wire n_17;
wire n_15;
wire n_224;
wire n_218;
wire n_19;
wire n_16;
wire n_160;
wire n_223;
wire n_131;
wire n_222;
wire n_230;
wire n_27;
wire n_20;
wire n_213;
wire n_132;
wire n_26;
wire n_21;
wire n_159;
wire n_202;
wire n_24;
wire n_22;
wire n_158;
wire n_200;
wire n_29;
wire n_23;
wire n_157;
wire n_209;
wire n_25;
wire n_203;
wire n_215;
wire n_117;
wire n_234;
wire n_233;
wire n_207;
wire n_208;
wire n_156;
wire n_30;
wire n_155;
wire n_88;
wire n_31;
wire n_35;
wire n_37;
wire n_36;
wire n_33;
wire n_32;
wire n_91;
wire n_87;
wire n_89;
wire n_85;
wire n_38;
wire n_34;
wire n_84;
wire n_154;
wire n_90;
wire n_133;
wire n_240;
wire n_153;
wire n_152;
wire n_39;
wire n_120;
wire n_137;
wire n_40;
wire n_44;
wire n_46;
wire n_45;
wire n_42;
wire n_41;
wire n_83;
wire n_80;
wire n_81;
wire n_78;
wire n_47;
wire n_43;
wire n_77;
wire n_185;
wire n_82;
wire n_151;
wire n_150;
wire n_149;
wire n_148;
wire n_48;
wire n_121;
wire n_141;
wire n_49;
wire n_53;
wire n_55;
wire n_54;
wire n_51;
wire n_50;
wire n_76;
wire n_73;
wire n_74;
wire n_71;
wire n_56;
wire n_52;
wire n_70;
wire n_172;
wire n_75;
wire n_179;
wire n_147;
wire n_146;
wire n_68;
wire n_63;
wire n_58;
wire n_57;
wire n_145;
wire n_64;
wire n_67;
wire n_122;
wire n_60;
wire n_59;
wire n_61;
wire n_66;
wire n_65;
wire n_62;
wire n_69;
wire n_164;
wire n_163;
wire n_143;
wire n_72;
wire n_142;
wire n_139;
wire n_79;
wire n_138;
wire n_135;
wire n_86;
wire n_134;
wire n_92;
wire n_94;
wire n_98;
wire n_106;
wire n_103;
wire n_107;
wire n_99;
wire n_125;
wire n_105;
wire n_113;
wire n_220;
wire n_119;
wire n_136;
wire n_140;
wire n_144;
wire n_176;
wire n_180;
wire n_190;
wire n_235;
wire n_191;
wire n_239;
wire n_195;
wire n_196;
wire n_211;
wire n_165;
wire n_162;
wire n_167;
wire n_173;
wire n_169;
wire n_243;
wire n_166;
wire n_168;
wire n_242;
wire n_171;
wire n_170;
wire n_178;
wire n_174;
wire n_175;
wire n_186;
wire n_181;
wire n_183;
wire n_182;
wire n_184;
wire n_189;
wire n_187;
wire n_188;
wire n_192;
wire n_193;
wire n_194;
wire n_241;
wire n_204;
wire n_197;
wire n_198;
wire n_201;
wire n_199;
wire n_212;
wire n_205;
wire n_210;
wire n_214;
wire n_206;
wire n_231;
wire n_216;
wire n_219;
wire n_217;
wire n_226;
wire n_221;
wire n_228;
wire n_225;
wire n_232;
wire n_236;
wire n_237;


INV_X1 i_275 (.ZN (n_243), .A (multiplicand[28]));
INV_X1 i_274 (.ZN (n_242), .A (A[28]));
NAND2_X1 i_273 (.ZN (n_241), .A1 (multiplicand[19]), .A2 (n_136));
INV_X1 i_272 (.ZN (n_240), .A (n_241));
INV_X1 i_271 (.ZN (n_239), .A (n_89));
INV_X1 i_269 (.ZN (n_237), .A (n_86));
NAND3_X1 i_268 (.ZN (n_236), .A1 (n_237), .A2 (n_239), .A3 (n_91));
AOI21_X1 i_267 (.ZN (n_235), .A (n_240), .B1 (n_236), .B2 (n_84));
NOR3_X1 i_266 (.ZN (n_234), .A1 (n_97), .A2 (n_112), .A3 (n_113));
OAI221_X1 i_265 (.ZN (n_233), .A (n_92), .B1 (multiplicand[7]), .B2 (n_130), .C1 (n_113), .C2 (n_94));
OR2_X1 i_264 (.ZN (n_232), .A1 (n_233), .A2 (n_234));
INV_X1 i_263 (.ZN (n_231), .A (n_232));
INV_X1 i_262 (.ZN (n_230), .A (A[11]));
NOR2_X1 i_261 (.ZN (n_229), .A1 (multiplicand[8]), .A2 (n_131));
INV_X1 i_260 (.ZN (n_228), .A (A[9]));
NOR2_X1 i_259 (.ZN (n_227), .A1 (multiplicand[9]), .A2 (n_228));
INV_X1 i_258 (.ZN (n_226), .A (A[10]));
NAND2_X1 i_257 (.ZN (n_225), .A1 (multiplicand[10]), .A2 (n_226));
INV_X1 i_256 (.ZN (n_224), .A (n_225));
NAND2_X1 i_255 (.ZN (n_223), .A1 (multiplicand[9]), .A2 (n_228));
NAND2_X1 i_254 (.ZN (n_222), .A1 (multiplicand[11]), .A2 (n_230));
NAND2_X1 i_253 (.ZN (n_221), .A1 (n_223), .A2 (n_222));
NOR2_X1 i_252 (.ZN (n_220), .A1 (n_224), .A2 (n_221));
OAI21_X1 i_251 (.ZN (n_219), .A (n_220), .B1 (n_229), .B2 (n_227));
NOR2_X1 i_250 (.ZN (n_218), .A1 (multiplicand[10]), .A2 (n_226));
NAND2_X1 i_249 (.ZN (n_217), .A1 (n_218), .A2 (n_222));
OAI211_X1 i_248 (.ZN (n_216), .A (n_219), .B (n_217), .C1 (n_230), .C2 (multiplicand[11]));
INV_X1 i_247 (.ZN (n_215), .A (n_216));
OAI21_X1 i_246 (.ZN (n_214), .A (n_215), .B1 (n_117), .B2 (n_231));
NAND2_X1 i_245 (.ZN (n_213), .A1 (multiplicand[12]), .A2 (n_132));
INV_X1 i_244 (.ZN (n_212), .A (A[14]));
NAND2_X1 i_243 (.ZN (n_211), .A1 (multiplicand[14]), .A2 (n_212));
INV_X1 i_242 (.ZN (n_210), .A (A[13]));
NAND2_X1 i_241 (.ZN (n_209), .A1 (multiplicand[13]), .A2 (n_210));
INV_X1 i_240 (.ZN (n_208), .A (A[15]));
NAND2_X1 i_239 (.ZN (n_207), .A1 (multiplicand[15]), .A2 (n_208));
NAND2_X1 i_238 (.ZN (n_206), .A1 (n_209), .A2 (n_207));
INV_X1 i_237 (.ZN (n_205), .A (n_206));
NAND4_X1 i_236 (.ZN (n_204), .A1 (n_214), .A2 (n_213), .A3 (n_211), .A4 (n_205));
NOR2_X1 i_235 (.ZN (n_203), .A1 (multiplicand[12]), .A2 (n_132));
NOR2_X1 i_234 (.ZN (n_202), .A1 (multiplicand[13]), .A2 (n_210));
OAI211_X1 i_233 (.ZN (n_201), .A (n_211), .B (n_205), .C1 (n_203), .C2 (n_202));
NOR2_X1 i_232 (.ZN (n_200), .A1 (multiplicand[14]), .A2 (n_212));
NAND2_X1 i_231 (.ZN (n_199), .A1 (n_200), .A2 (n_207));
OAI211_X1 i_230 (.ZN (n_198), .A (n_201), .B (n_199), .C1 (n_208), .C2 (multiplicand[15]));
INV_X1 i_229 (.ZN (n_197), .A (n_198));
NAND2_X1 i_228 (.ZN (n_196), .A1 (n_204), .A2 (n_197));
NAND2_X1 i_227 (.ZN (n_195), .A1 (multiplicand[16]), .A2 (n_133));
NAND3_X1 i_226 (.ZN (n_194), .A1 (n_196), .A2 (n_241), .A3 (n_195));
INV_X1 i_225 (.ZN (n_193), .A (n_194));
NAND3_X1 i_224 (.ZN (n_192), .A1 (n_91), .A2 (n_193), .A3 (n_239));
OAI21_X1 i_223 (.ZN (n_191), .A (n_192), .B1 (multiplicand[19]), .B2 (n_136));
NAND2_X1 i_222 (.ZN (n_190), .A1 (multiplicand[23]), .A2 (n_140));
NOR2_X1 i_221 (.ZN (n_189), .A1 (n_82), .A2 (n_81));
OAI211_X1 i_220 (.ZN (n_188), .A (n_190), .B (n_189), .C1 (A[20]), .C2 (n_120));
INV_X1 i_219 (.ZN (n_187), .A (n_188));
OAI21_X1 i_218 (.ZN (n_186), .A (n_187), .B1 (n_235), .B2 (n_191));
INV_X1 i_217 (.ZN (n_185), .A (n_189));
OR2_X1 i_216 (.ZN (n_184), .A1 (n_185), .A2 (n_79));
INV_X1 i_215 (.ZN (n_183), .A (n_184));
OAI21_X1 i_214 (.ZN (n_182), .A (n_77), .B1 (multiplicand[23]), .B2 (n_140));
OAI21_X1 i_213 (.ZN (n_181), .A (n_190), .B1 (n_183), .B2 (n_182));
NAND2_X1 i_212 (.ZN (n_180), .A1 (n_186), .A2 (n_181));
NOR2_X1 i_211 (.ZN (n_179), .A1 (n_121), .A2 (A[24]));
INV_X1 i_210 (.ZN (n_178), .A (n_74));
NAND2_X1 i_208 (.ZN (n_176), .A1 (multiplicand[27]), .A2 (n_144));
NAND3_X1 i_207 (.ZN (n_175), .A1 (n_76), .A2 (n_178), .A3 (n_176));
NOR2_X1 i_206 (.ZN (n_174), .A1 (n_175), .A2 (n_179));
NAND2_X1 i_205 (.ZN (n_173), .A1 (n_180), .A2 (n_174));
NAND2_X1 i_204 (.ZN (n_172), .A1 (n_76), .A2 (n_178));
NOR2_X1 i_203 (.ZN (n_171), .A1 (n_172), .A2 (n_72));
OAI21_X1 i_202 (.ZN (n_170), .A (n_70), .B1 (multiplicand[27]), .B2 (n_144));
OAI21_X1 i_201 (.ZN (n_169), .A (n_176), .B1 (n_171), .B2 (n_170));
AOI21_X1 i_200 (.ZN (n_168), .A (n_242), .B1 (n_173), .B2 (n_169));
NAND3_X1 i_199 (.ZN (n_167), .A1 (n_173), .A2 (n_242), .A3 (n_169));
INV_X1 i_198 (.ZN (n_166), .A (n_167));
OAI21_X1 i_197 (.ZN (n_165), .A (n_243), .B1 (n_166), .B2 (n_168));
NAND2_X1 i_196 (.ZN (n_164), .A1 (n_173), .A2 (n_169));
NAND2_X1 i_195 (.ZN (n_163), .A1 (n_164), .A2 (A[28]));
NAND3_X1 i_194 (.ZN (n_162), .A1 (n_163), .A2 (multiplicand[28]), .A3 (n_167));
NAND2_X1 i_193 (.ZN (p_0[28]), .A1 (n_165), .A2 (n_162));
INV_X1 i_192 (.ZN (n_161), .A (n_223));
INV_X1 i_191 (.ZN (n_160), .A (n_218));
INV_X1 i_190 (.ZN (n_159), .A (n_209));
INV_X1 i_189 (.ZN (n_158), .A (n_211));
INV_X1 i_188 (.ZN (n_157), .A (n_200));
INV_X1 i_187 (.ZN (n_156), .A (n_196));
INV_X1 i_186 (.ZN (n_155), .A (n_195));
NAND2_X1 i_185 (.ZN (n_154), .A1 (n_91), .A2 (n_239));
NOR2_X1 i_184 (.ZN (n_153), .A1 (multiplicand[19]), .A2 (n_136));
NOR2_X1 i_183 (.ZN (n_152), .A1 (n_235), .A2 (n_191));
NOR2_X1 i_182 (.ZN (n_151), .A1 (n_120), .A2 (A[20]));
INV_X1 i_181 (.ZN (n_150), .A (n_190));
NOR2_X1 i_180 (.ZN (n_149), .A1 (multiplicand[23]), .A2 (n_140));
INV_X1 i_179 (.ZN (n_148), .A (n_180));
INV_X1 i_178 (.ZN (n_147), .A (n_176));
NOR2_X1 i_177 (.ZN (n_146), .A1 (multiplicand[27]), .A2 (n_144));
INV_X1 i_176 (.ZN (n_145), .A (A[29]));
INV_X1 i_175 (.ZN (n_144), .A (A[27]));
INV_X1 i_174 (.ZN (n_143), .A (A[26]));
INV_X1 i_173 (.ZN (n_142), .A (A[25]));
INV_X1 i_172 (.ZN (n_141), .A (A[24]));
INV_X1 i_171 (.ZN (n_140), .A (A[23]));
INV_X1 i_170 (.ZN (n_139), .A (A[22]));
INV_X1 i_169 (.ZN (n_138), .A (A[21]));
INV_X1 i_168 (.ZN (n_137), .A (A[20]));
INV_X1 i_167 (.ZN (n_136), .A (A[19]));
INV_X1 i_166 (.ZN (n_135), .A (A[18]));
INV_X1 i_165 (.ZN (n_134), .A (A[17]));
INV_X1 i_164 (.ZN (n_133), .A (A[16]));
INV_X1 i_163 (.ZN (n_132), .A (A[12]));
INV_X1 i_162 (.ZN (n_131), .A (A[8]));
INV_X1 i_161 (.ZN (n_130), .A (A[7]));
INV_X1 i_160 (.ZN (n_129), .A (A[6]));
INV_X1 i_159 (.ZN (n_128), .A (A[5]));
INV_X1 i_158 (.ZN (n_127), .A (A[4]));
INV_X1 i_157 (.ZN (n_126), .A (A[3]));
INV_X1 i_156 (.ZN (n_125), .A (A[2]));
INV_X1 i_155 (.ZN (n_124), .A (A[1]));
INV_X1 i_154 (.ZN (n_123), .A (A[0]));
INV_X1 i_153 (.ZN (n_122), .A (multiplicand[30]));
INV_X1 i_152 (.ZN (n_121), .A (multiplicand[24]));
INV_X1 i_151 (.ZN (n_120), .A (multiplicand[20]));
NAND2_X1 i_150 (.ZN (n_119), .A1 (n_131), .A2 (multiplicand[8]));
INV_X1 i_149 (.ZN (n_118), .A (n_119));
NAND2_X1 i_148 (.ZN (n_117), .A1 (n_220), .A2 (n_119));
NAND2_X1 i_147 (.ZN (n_116), .A1 (n_129), .A2 (multiplicand[6]));
NAND2_X1 i_146 (.ZN (n_115), .A1 (n_128), .A2 (multiplicand[5]));
NAND2_X1 i_145 (.ZN (n_114), .A1 (n_130), .A2 (multiplicand[7]));
NAND3_X1 i_144 (.ZN (n_113), .A1 (n_116), .A2 (n_114), .A3 (n_115));
AND2_X1 i_143 (.ZN (n_112), .A1 (n_127), .A2 (multiplicand[4]));
AND2_X1 i_142 (.ZN (n_111), .A1 (n_124), .A2 (multiplicand[1]));
NAND2_X1 i_141 (.ZN (n_110), .A1 (n_125), .A2 (multiplicand[2]));
INV_X1 i_140 (.ZN (n_109), .A (n_110));
NAND2_X1 i_139 (.ZN (n_108), .A1 (n_126), .A2 (multiplicand[3]));
INV_X1 i_138 (.ZN (n_107), .A (n_108));
NOR3_X1 i_137 (.ZN (n_106), .A1 (n_111), .A2 (n_107), .A3 (n_109));
NOR2_X1 i_136 (.ZN (n_105), .A1 (n_123), .A2 (multiplicand[0]));
NOR2_X1 i_135 (.ZN (n_104), .A1 (n_124), .A2 (multiplicand[1]));
OAI21_X1 i_134 (.ZN (n_103), .A (n_106), .B1 (n_105), .B2 (n_104));
NAND2_X1 i_133 (.ZN (n_102), .A1 (n_123), .A2 (multiplicand[0]));
INV_X1 i_132 (.ZN (n_101), .A (n_102));
NOR2_X1 i_131 (.ZN (n_100), .A1 (n_125), .A2 (multiplicand[2]));
INV_X1 i_130 (.ZN (n_99), .A (n_100));
OAI221_X1 i_129 (.ZN (n_98), .A (n_103), .B1 (n_107), .B2 (n_99), .C1 (n_126), .C2 (multiplicand[3]));
AOI21_X1 i_128 (.ZN (n_97), .A (n_98), .B1 (n_106), .B2 (n_102));
NOR2_X1 i_127 (.ZN (n_96), .A1 (n_127), .A2 (multiplicand[4]));
NOR2_X1 i_126 (.ZN (n_95), .A1 (n_128), .A2 (multiplicand[5]));
NOR2_X1 i_125 (.ZN (n_94), .A1 (n_96), .A2 (n_95));
NOR2_X1 i_124 (.ZN (n_93), .A1 (n_129), .A2 (multiplicand[6]));
NAND2_X1 i_123 (.ZN (n_92), .A1 (n_114), .A2 (n_93));
NAND2_X1 i_122 (.ZN (n_91), .A1 (n_134), .A2 (multiplicand[17]));
INV_X1 i_121 (.ZN (n_90), .A (n_91));
AND2_X1 i_120 (.ZN (n_89), .A1 (n_135), .A2 (multiplicand[18]));
NOR2_X1 i_119 (.ZN (n_88), .A1 (n_133), .A2 (multiplicand[16]));
NOR2_X1 i_118 (.ZN (n_87), .A1 (n_134), .A2 (multiplicand[17]));
NOR2_X1 i_117 (.ZN (n_86), .A1 (n_88), .A2 (n_87));
NOR2_X1 i_116 (.ZN (n_85), .A1 (n_135), .A2 (multiplicand[18]));
INV_X1 i_115 (.ZN (n_84), .A (n_85));
NAND2_X1 i_114 (.ZN (n_83), .A1 (n_138), .A2 (multiplicand[21]));
INV_X1 i_113 (.ZN (n_82), .A (n_83));
AND2_X1 i_112 (.ZN (n_81), .A1 (n_139), .A2 (multiplicand[22]));
NOR2_X1 i_111 (.ZN (n_80), .A1 (n_138), .A2 (multiplicand[21]));
AOI21_X1 i_110 (.ZN (n_79), .A (n_80), .B1 (A[20]), .B2 (n_120));
NOR2_X1 i_109 (.ZN (n_78), .A1 (n_139), .A2 (multiplicand[22]));
INV_X1 i_108 (.ZN (n_77), .A (n_78));
NAND2_X1 i_107 (.ZN (n_76), .A1 (n_142), .A2 (multiplicand[25]));
INV_X1 i_106 (.ZN (n_75), .A (n_76));
AND2_X1 i_105 (.ZN (n_74), .A1 (n_143), .A2 (multiplicand[26]));
NOR2_X1 i_104 (.ZN (n_73), .A1 (n_142), .A2 (multiplicand[25]));
AOI21_X1 i_103 (.ZN (n_72), .A (n_73), .B1 (A[24]), .B2 (n_121));
NOR2_X1 i_102 (.ZN (n_71), .A1 (n_143), .A2 (multiplicand[26]));
INV_X1 i_101 (.ZN (n_70), .A (n_71));
NAND2_X1 i_100 (.ZN (n_69), .A1 (multiplicand[28]), .A2 (n_163));
OAI21_X1 i_99 (.ZN (n_68), .A (n_69), .B1 (A[28]), .B2 (n_164));
NAND2_X1 i_98 (.ZN (n_67), .A1 (A[31]), .A2 (n_122));
INV_X1 i_97 (.ZN (n_66), .A (n_67));
NAND2_X1 i_96 (.ZN (n_65), .A1 (n_145), .A2 (multiplicand[29]));
INV_X1 i_95 (.ZN (n_64), .A (n_65));
OAI21_X1 i_94 (.ZN (n_63), .A (n_65), .B1 (n_145), .B2 (multiplicand[29]));
INV_X1 i_93 (.ZN (n_62), .A (n_63));
NAND3_X1 i_92 (.ZN (n_61), .A1 (n_67), .A2 (n_62), .A3 (n_68));
OAI221_X1 i_91 (.ZN (n_60), .A (n_61), .B1 (A[31]), .B2 (n_122), .C1 (n_66), .C2 (n_65));
XOR2_X1 i_90 (.Z (n_59), .A (A[31]), .B (multiplicand[31]));
XOR2_X1 i_89 (.Z (p_0[31]), .A (n_60), .B (n_59));
OAI21_X1 i_88 (.ZN (n_58), .A (n_67), .B1 (A[31]), .B2 (n_122));
OAI22_X1 i_87 (.ZN (n_57), .A1 (n_145), .A2 (multiplicand[29]), .B1 (n_68), .B2 (n_64));
XNOR2_X1 i_86 (.ZN (p_0[30]), .A (n_58), .B (n_57));
XOR2_X1 i_85 (.Z (p_0[29]), .A (n_68), .B (n_63));
NOR2_X1 i_84 (.ZN (n_56), .A1 (n_147), .A2 (n_146));
OAI22_X1 i_83 (.ZN (n_55), .A1 (n_141), .A2 (multiplicand[24]), .B1 (n_148), .B2 (n_179));
OR2_X1 i_82 (.ZN (n_54), .A1 (n_75), .A2 (n_73));
NOR2_X1 i_81 (.ZN (n_53), .A1 (n_55), .A2 (n_54));
OAI21_X1 i_80 (.ZN (n_52), .A (n_70), .B1 (n_172), .B2 (n_53));
XOR2_X1 i_79 (.Z (p_0[27]), .A (n_56), .B (n_52));
NOR2_X1 i_78 (.ZN (n_51), .A1 (n_74), .A2 (n_71));
OAI21_X1 i_77 (.ZN (n_50), .A (n_76), .B1 (n_73), .B2 (n_55));
XNOR2_X1 i_76 (.ZN (p_0[26]), .A (n_51), .B (n_50));
AOI21_X1 i_75 (.ZN (n_49), .A (n_53), .B1 (n_55), .B2 (n_54));
INV_X1 i_74 (.ZN (p_0[25]), .A (n_49));
OAI22_X1 i_73 (.ZN (n_48), .A1 (A[24]), .A2 (n_121), .B1 (n_141), .B2 (multiplicand[24]));
XOR2_X1 i_72 (.Z (p_0[24]), .A (n_148), .B (n_48));
NOR2_X1 i_71 (.ZN (n_47), .A1 (n_150), .A2 (n_149));
OAI22_X1 i_70 (.ZN (n_46), .A1 (n_137), .A2 (multiplicand[20]), .B1 (n_152), .B2 (n_151));
OR2_X1 i_69 (.ZN (n_45), .A1 (n_82), .A2 (n_80));
NOR2_X1 i_68 (.ZN (n_44), .A1 (n_46), .A2 (n_45));
OAI21_X1 i_67 (.ZN (n_43), .A (n_77), .B1 (n_185), .B2 (n_44));
XOR2_X1 i_66 (.Z (p_0[23]), .A (n_47), .B (n_43));
NOR2_X1 i_65 (.ZN (n_42), .A1 (n_81), .A2 (n_78));
OAI21_X1 i_64 (.ZN (n_41), .A (n_83), .B1 (n_80), .B2 (n_46));
XNOR2_X1 i_63 (.ZN (p_0[22]), .A (n_42), .B (n_41));
AOI21_X1 i_62 (.ZN (n_40), .A (n_44), .B1 (n_46), .B2 (n_45));
INV_X1 i_61 (.ZN (p_0[21]), .A (n_40));
OAI22_X1 i_60 (.ZN (n_39), .A1 (A[20]), .A2 (n_120), .B1 (n_137), .B2 (multiplicand[20]));
XOR2_X1 i_59 (.Z (p_0[20]), .A (n_152), .B (n_39));
NOR2_X1 i_58 (.ZN (n_38), .A1 (n_240), .A2 (n_153));
OAI22_X1 i_57 (.ZN (n_37), .A1 (n_133), .A2 (multiplicand[16]), .B1 (n_156), .B2 (n_155));
OR2_X1 i_56 (.ZN (n_36), .A1 (n_90), .A2 (n_87));
NOR2_X1 i_55 (.ZN (n_35), .A1 (n_37), .A2 (n_36));
OAI21_X1 i_54 (.ZN (n_34), .A (n_84), .B1 (n_154), .B2 (n_35));
XOR2_X1 i_53 (.Z (p_0[19]), .A (n_38), .B (n_34));
NOR2_X1 i_52 (.ZN (n_33), .A1 (n_89), .A2 (n_85));
OAI21_X1 i_51 (.ZN (n_32), .A (n_91), .B1 (n_87), .B2 (n_37));
XNOR2_X1 i_50 (.ZN (p_0[18]), .A (n_33), .B (n_32));
AOI21_X1 i_49 (.ZN (n_31), .A (n_35), .B1 (n_37), .B2 (n_36));
INV_X1 i_48 (.ZN (p_0[17]), .A (n_31));
NOR2_X1 i_47 (.ZN (n_30), .A1 (n_155), .A2 (n_88));
XNOR2_X1 i_46 (.ZN (p_0[16]), .A (n_156), .B (n_30));
OAI21_X1 i_45 (.ZN (n_29), .A (n_207), .B1 (n_208), .B2 (multiplicand[15]));
NOR2_X1 i_44 (.ZN (n_28), .A1 (n_234), .A2 (n_233));
OAI21_X1 i_43 (.ZN (n_27), .A (n_215), .B1 (n_117), .B2 (n_28));
OAI21_X1 i_42 (.ZN (n_26), .A (n_213), .B1 (n_203), .B2 (n_27));
INV_X1 i_41 (.ZN (n_25), .A (n_26));
OAI21_X1 i_40 (.ZN (n_24), .A (n_209), .B1 (n_202), .B2 (n_25));
OAI21_X1 i_39 (.ZN (n_23), .A (n_157), .B1 (n_158), .B2 (n_24));
XNOR2_X1 i_38 (.ZN (p_0[15]), .A (n_29), .B (n_23));
NOR2_X1 i_37 (.ZN (n_22), .A1 (n_158), .A2 (n_200));
XNOR2_X1 i_36 (.ZN (p_0[14]), .A (n_24), .B (n_22));
NOR2_X1 i_35 (.ZN (n_21), .A1 (n_159), .A2 (n_202));
XNOR2_X1 i_34 (.ZN (p_0[13]), .A (n_26), .B (n_21));
OAI21_X1 i_33 (.ZN (n_20), .A (n_213), .B1 (n_132), .B2 (multiplicand[12]));
XNOR2_X1 i_32 (.ZN (p_0[12]), .A (n_27), .B (n_20));
OAI21_X1 i_31 (.ZN (n_19), .A (n_222), .B1 (n_230), .B2 (multiplicand[11]));
OAI22_X1 i_30 (.ZN (n_18), .A1 (n_131), .A2 (multiplicand[8]), .B1 (n_118), .B2 (n_28));
OAI21_X1 i_29 (.ZN (n_17), .A (n_223), .B1 (n_227), .B2 (n_18));
OAI21_X1 i_28 (.ZN (n_16), .A (n_160), .B1 (n_224), .B2 (n_17));
XNOR2_X1 i_27 (.ZN (p_0[11]), .A (n_19), .B (n_16));
NOR2_X1 i_26 (.ZN (n_15), .A1 (n_224), .A2 (n_218));
XNOR2_X1 i_25 (.ZN (p_0[10]), .A (n_17), .B (n_15));
NOR2_X1 i_24 (.ZN (n_14), .A1 (n_161), .A2 (n_227));
XOR2_X1 i_23 (.Z (p_0[9]), .A (n_18), .B (n_14));
NOR2_X1 i_22 (.ZN (n_13), .A1 (n_118), .A2 (n_229));
XNOR2_X1 i_21 (.ZN (p_0[8]), .A (n_28), .B (n_13));
OAI21_X1 i_20 (.ZN (n_12), .A (n_114), .B1 (n_130), .B2 (multiplicand[7]));
OAI22_X1 i_19 (.ZN (n_11), .A1 (n_112), .A2 (n_97), .B1 (n_127), .B2 (multiplicand[4]));
OAI21_X1 i_18 (.ZN (n_10), .A (n_115), .B1 (n_95), .B2 (n_11));
INV_X1 i_17 (.ZN (n_9), .A (n_10));
OAI21_X1 i_16 (.ZN (n_8), .A (n_116), .B1 (n_93), .B2 (n_9));
XOR2_X1 i_15 (.Z (p_0[7]), .A (n_12), .B (n_8));
OAI21_X1 i_14 (.ZN (n_7), .A (n_116), .B1 (n_129), .B2 (multiplicand[6]));
XNOR2_X1 i_13 (.ZN (p_0[6]), .A (n_9), .B (n_7));
OAI21_X1 i_12 (.ZN (n_6), .A (n_115), .B1 (n_128), .B2 (multiplicand[5]));
XNOR2_X1 i_11 (.ZN (p_0[5]), .A (n_11), .B (n_6));
NOR2_X1 i_10 (.ZN (n_5), .A1 (n_112), .A2 (n_96));
XNOR2_X1 i_9 (.ZN (p_0[4]), .A (n_97), .B (n_5));
OAI21_X1 i_8 (.ZN (n_4), .A (n_108), .B1 (n_126), .B2 (multiplicand[3]));
OAI22_X1 i_7 (.ZN (n_3), .A1 (n_124), .A2 (multiplicand[1]), .B1 (n_111), .B2 (n_101));
OAI21_X1 i_6 (.ZN (n_2), .A (n_110), .B1 (n_100), .B2 (n_3));
XOR2_X1 i_5 (.Z (p_0[3]), .A (n_4), .B (n_2));
NOR2_X1 i_4 (.ZN (n_1), .A1 (n_109), .A2 (n_100));
XOR2_X1 i_3 (.Z (p_0[2]), .A (n_3), .B (n_1));
NOR2_X1 i_2 (.ZN (n_0), .A1 (n_111), .A2 (n_104));
XNOR2_X1 i_1 (.ZN (p_0[1]), .A (n_101), .B (n_0));
OAI21_X1 i_0 (.ZN (p_0[0]), .A (n_102), .B1 (n_123), .B2 (multiplicand[0]));

endmodule //datapath__0_65

module datapath (p_0, a);

output [31:0] p_0;
input [31:0] a;
wire n_62;
wire n_60;
wire n_61;
wire n_58;
wire n_59;
wire n_5;
wire n_57;
wire n_1;
wire n_55;
wire n_0;
wire n_56;
wire n_11;
wire n_54;
wire n_7;
wire n_52;
wire n_6;
wire n_53;
wire n_17;
wire n_51;
wire n_13;
wire n_49;
wire n_12;
wire n_50;
wire n_23;
wire n_48;
wire n_21;
wire n_22;
wire n_19;
wire n_20;
wire n_45;
wire n_18;
wire n_46;
wire n_25;
wire n_44;
wire n_37;
wire n_38;
wire n_4;
wire n_74;
wire n_39;
wire n_29;
wire n_10;
wire n_26;
wire n_16;
wire n_24;
wire n_27;
wire n_28;
wire n_30;
wire n_32;
wire n_31;
wire n_33;
wire n_34;
wire n_40;
wire n_42;
wire n_41;
wire n_43;
wire n_47;
wire n_63;
wire n_84;
wire n_65;
wire n_64;
wire n_66;
wire n_83;
wire n_67;
wire n_85;
wire n_68;
wire n_69;
wire n_70;
wire n_82;
wire n_72;
wire n_80;
wire n_79;
wire n_75;
wire n_71;
wire n_78;
wire n_101;
wire n_73;
wire n_76;
wire n_77;
wire n_81;
wire n_100;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_99;
wire n_98;
wire n_97;
wire n_96;


INV_X1 i_132 (.ZN (n_101), .A (a[28]));
INV_X1 i_131 (.ZN (n_100), .A (a[23]));
INV_X1 i_130 (.ZN (n_99), .A (a[3]));
INV_X1 i_129 (.ZN (n_98), .A (a[2]));
INV_X1 i_128 (.ZN (n_97), .A (a[1]));
INV_X1 i_127 (.ZN (n_96), .A (a[0]));
NAND2_X1 i_126 (.ZN (n_61), .A1 (n_97), .A2 (n_96));
INV_X1 i_125 (.ZN (n_62), .A (n_61));
NAND2_X1 i_124 (.ZN (n_59), .A1 (n_62), .A2 (n_98));
INV_X1 i_123 (.ZN (n_60), .A (n_59));
NAND2_X1 i_122 (.ZN (n_57), .A1 (n_60), .A2 (n_99));
INV_X1 i_121 (.ZN (n_58), .A (n_57));
OR3_X1 i_120 (.ZN (n_56), .A1 (a[6]), .A2 (a[5]), .A3 (a[4]));
OR2_X1 i_119 (.ZN (n_95), .A1 (n_56), .A2 (a[7]));
INV_X1 i_118 (.ZN (n_94), .A (n_95));
NAND2_X1 i_117 (.ZN (n_54), .A1 (n_94), .A2 (n_58));
INV_X1 i_116 (.ZN (n_55), .A (n_54));
OR3_X1 i_115 (.ZN (n_53), .A1 (a[10]), .A2 (a[9]), .A3 (a[8]));
OR2_X1 i_114 (.ZN (n_93), .A1 (n_53), .A2 (a[11]));
INV_X1 i_113 (.ZN (n_92), .A (n_93));
NAND2_X1 i_112 (.ZN (n_51), .A1 (n_55), .A2 (n_92));
INV_X1 i_111 (.ZN (n_52), .A (n_51));
OR3_X1 i_110 (.ZN (n_50), .A1 (a[14]), .A2 (a[13]), .A3 (a[12]));
OR2_X1 i_109 (.ZN (n_91), .A1 (n_50), .A2 (a[15]));
INV_X1 i_108 (.ZN (n_90), .A (n_91));
NAND2_X1 i_107 (.ZN (n_48), .A1 (n_52), .A2 (n_90));
INV_X1 i_106 (.ZN (n_49), .A (n_48));
OR3_X1 i_105 (.ZN (n_46), .A1 (a[18]), .A2 (a[17]), .A3 (a[16]));
OR2_X1 i_104 (.ZN (n_89), .A1 (n_46), .A2 (a[19]));
INV_X1 i_103 (.ZN (n_88), .A (n_89));
NAND2_X1 i_102 (.ZN (n_44), .A1 (n_49), .A2 (n_88));
INV_X1 i_101 (.ZN (n_45), .A (n_44));
OR3_X1 i_100 (.ZN (n_87), .A1 (a[22]), .A2 (a[21]), .A3 (a[20]));
INV_X1 i_99 (.ZN (n_86), .A (n_87));
NAND2_X1 i_98 (.ZN (n_85), .A1 (n_45), .A2 (n_86));
INV_X1 i_97 (.ZN (n_84), .A (n_85));
NAND2_X1 i_96 (.ZN (n_83), .A1 (n_84), .A2 (n_100));
INV_X1 i_95 (.ZN (n_82), .A (n_83));
INV_X1 i_94 (.ZN (n_81), .A (a[26]));
INV_X1 i_93 (.ZN (n_80), .A (a[25]));
INV_X1 i_92 (.ZN (n_79), .A (a[24]));
NAND3_X1 i_91 (.ZN (n_78), .A1 (n_81), .A2 (n_80), .A3 (n_79));
OR2_X1 i_90 (.ZN (n_77), .A1 (n_78), .A2 (a[27]));
INV_X1 i_89 (.ZN (n_76), .A (n_77));
NAND2_X1 i_88 (.ZN (n_38), .A1 (n_82), .A2 (n_76));
INV_X1 i_87 (.ZN (n_75), .A (n_38));
NAND2_X1 i_86 (.ZN (n_74), .A1 (n_75), .A2 (n_101));
XNOR2_X1 i_85 (.ZN (n_73), .A (n_74), .B (a[29]));
INV_X1 i_84 (.ZN (p_0[29]), .A (n_73));
XNOR2_X1 i_83 (.ZN (p_0[28]), .A (n_38), .B (n_101));
INV_X1 i_82 (.ZN (n_72), .A (n_78));
NAND2_X1 i_81 (.ZN (n_71), .A1 (n_82), .A2 (n_72));
AOI21_X1 i_80 (.ZN (p_0[27]), .A (n_75), .B1 (n_71), .B2 (a[27]));
NAND3_X1 i_79 (.ZN (n_70), .A1 (n_82), .A2 (n_80), .A3 (n_79));
AOI22_X1 i_78 (.ZN (p_0[26]), .A1 (n_70), .A2 (a[26]), .B1 (n_82), .B2 (n_72));
OAI21_X1 i_77 (.ZN (n_69), .A (a[25]), .B1 (n_83), .B2 (a[24]));
AND2_X1 i_76 (.ZN (p_0[25]), .A1 (n_69), .A2 (n_70));
XNOR2_X1 i_75 (.ZN (n_68), .A (n_83), .B (a[24]));
INV_X1 i_74 (.ZN (p_0[24]), .A (n_68));
NAND2_X1 i_73 (.ZN (n_67), .A1 (n_85), .A2 (a[23]));
NAND2_X1 i_72 (.ZN (n_66), .A1 (n_83), .A2 (n_67));
INV_X1 i_71 (.ZN (p_0[23]), .A (n_66));
INV_X1 i_70 (.ZN (n_65), .A (a[21]));
INV_X1 i_69 (.ZN (n_64), .A (a[20]));
NAND3_X1 i_66 (.ZN (n_63), .A1 (n_45), .A2 (n_65), .A3 (n_64));
AOI21_X1 i_63 (.ZN (p_0[22]), .A (n_84), .B1 (n_63), .B2 (a[22]));
INV_X1 i_62 (.ZN (n_47), .A (n_25));
INV_X1 i_61 (.ZN (n_43), .A (n_63));
AOI21_X1 i_60 (.ZN (p_0[21]), .A (n_43), .B1 (n_47), .B2 (a[21]));
INV_X1 i_59 (.ZN (n_42), .A (a[13]));
INV_X1 i_58 (.ZN (n_41), .A (a[12]));
NAND2_X1 i_57 (.ZN (n_40), .A1 (n_52), .A2 (n_41));
INV_X1 i_56 (.ZN (n_17), .A (n_40));
NAND2_X1 i_55 (.ZN (n_39), .A1 (n_17), .A2 (n_42));
NAND2_X1 i_54 (.ZN (n_34), .A1 (n_40), .A2 (a[13]));
NAND2_X1 i_53 (.ZN (n_33), .A1 (n_39), .A2 (n_34));
INV_X1 i_52 (.ZN (p_0[13]), .A (n_33));
INV_X1 i_51 (.ZN (n_32), .A (a[9]));
INV_X1 i_50 (.ZN (n_31), .A (a[8]));
NAND2_X1 i_49 (.ZN (n_30), .A1 (n_55), .A2 (n_31));
INV_X1 i_48 (.ZN (n_11), .A (n_30));
NAND2_X1 i_47 (.ZN (n_29), .A1 (n_11), .A2 (n_32));
NAND2_X1 i_45 (.ZN (n_28), .A1 (n_30), .A2 (a[9]));
NAND2_X1 i_44 (.ZN (n_27), .A1 (n_29), .A2 (n_28));
INV_X1 i_32 (.ZN (p_0[9]), .A (n_27));
INV_X1 i_31 (.ZN (n_26), .A (a[5]));
INV_X1 i_30 (.ZN (n_24), .A (a[4]));
NAND2_X1 i_24 (.ZN (n_16), .A1 (n_58), .A2 (n_24));
XNOR2_X1 i_22 (.ZN (p_0[5]), .A (n_16), .B (n_26));
INV_X1 i_21 (.ZN (n_5), .A (n_16));
NAND2_X1 i_20 (.ZN (n_10), .A1 (n_5), .A2 (n_26));
OR2_X1 i_10 (.ZN (n_4), .A1 (n_74), .A2 (a[29]));
NOR4_X1 i_68 (.ZN (n_37), .A1 (a[29]), .A2 (a[28]), .A3 (a[30]), .A4 (n_38));
XNOR2_X1 i_67 (.ZN (p_0[31]), .A (a[31]), .B (n_37));
AOI21_X1 i_64 (.ZN (p_0[30]), .A (n_37), .B1 (a[30]), .B2 (n_4));
NOR2_X1 i_46 (.ZN (n_25), .A1 (a[20]), .A2 (n_44));
AOI21_X1 i_43 (.ZN (p_0[20]), .A (n_25), .B1 (a[20]), .B2 (n_44));
NOR2_X1 i_42 (.ZN (n_23), .A1 (a[16]), .A2 (n_48));
INV_X1 i_41 (.ZN (n_22), .A (n_23));
NOR2_X1 i_40 (.ZN (n_21), .A1 (a[17]), .A2 (n_22));
INV_X1 i_39 (.ZN (n_20), .A (n_21));
NOR2_X1 i_38 (.ZN (n_19), .A1 (n_48), .A2 (n_46));
INV_X1 i_37 (.ZN (n_18), .A (n_19));
AOI21_X1 i_36 (.ZN (p_0[19]), .A (n_45), .B1 (a[19]), .B2 (n_18));
AOI21_X1 i_35 (.ZN (p_0[18]), .A (n_19), .B1 (a[18]), .B2 (n_20));
AOI21_X1 i_34 (.ZN (p_0[17]), .A (n_21), .B1 (a[17]), .B2 (n_22));
AOI21_X1 i_33 (.ZN (p_0[16]), .A (n_23), .B1 (a[16]), .B2 (n_48));
NOR2_X1 i_28 (.ZN (n_13), .A1 (n_51), .A2 (n_50));
INV_X1 i_27 (.ZN (n_12), .A (n_13));
AOI21_X1 i_26 (.ZN (p_0[15]), .A (n_49), .B1 (a[15]), .B2 (n_12));
AOI21_X1 i_25 (.ZN (p_0[14]), .A (n_13), .B1 (a[14]), .B2 (n_39));
AOI21_X1 i_23 (.ZN (p_0[12]), .A (n_17), .B1 (a[12]), .B2 (n_51));
NOR2_X1 i_18 (.ZN (n_7), .A1 (n_54), .A2 (n_53));
INV_X1 i_17 (.ZN (n_6), .A (n_7));
AOI21_X1 i_16 (.ZN (p_0[11]), .A (n_52), .B1 (a[11]), .B2 (n_6));
AOI21_X1 i_15 (.ZN (p_0[10]), .A (n_7), .B1 (a[10]), .B2 (n_29));
AOI21_X1 i_13 (.ZN (p_0[8]), .A (n_11), .B1 (a[8]), .B2 (n_54));
NOR2_X1 i_8 (.ZN (n_1), .A1 (n_57), .A2 (n_56));
INV_X1 i_7 (.ZN (n_0), .A (n_1));
AOI21_X1 i_6 (.ZN (p_0[7]), .A (n_55), .B1 (a[7]), .B2 (n_0));
AOI21_X1 i_5 (.ZN (p_0[6]), .A (n_1), .B1 (a[6]), .B2 (n_10));
AOI21_X1 i_3 (.ZN (p_0[4]), .A (n_5), .B1 (a[4]), .B2 (n_57));
AOI21_X1 i_2 (.ZN (p_0[3]), .A (n_58), .B1 (a[3]), .B2 (n_59));
AOI21_X1 i_1 (.ZN (p_0[2]), .A (n_60), .B1 (a[2]), .B2 (n_61));
AOI21_X1 i_0 (.ZN (p_0[1]), .A (n_62), .B1 (a[1]), .B2 (a[0]));

endmodule //datapath

module booth_multiplier (clk, rst, en, a, b, c);

output [63:0] c;
input [31:0] a;
input [31:0] b;
input clk;
input en;
input rst;
wire CTS_n_tid0_336;
wire CTS_n_tid1_243;
wire n_64_3;
wire n_64_4;
wire n_64_5;
wire n_64_6;
wire n_64_7;
wire n_64_8;
wire n_64_9;
wire n_64_10;
wire n_64_11;
wire n_64_12;
wire n_64_13;
wire n_64_14;
wire n_64_15;
wire n_64_16;
wire n_64_17;
wire n_64_18;
wire n_64_19;
wire n_64_20;
wire n_64_21;
wire n_64_22;
wire n_64_23;
wire n_64_24;
wire n_64_25;
wire n_64_26;
wire n_64_27;
wire n_64_28;
wire n_64_29;
wire n_64_30;
wire n_64_31;
wire n_64_32;
wire n_64_33;
wire n_64_34;
wire n_64_35;
wire n_64_36;
wire n_64_37;
wire n_64_38;
wire n_64_39;
wire n_64_40;
wire n_64_41;
wire n_64_42;
wire n_64_43;
wire n_64_44;
wire n_64_45;
wire n_64_46;
wire n_64_47;
wire n_64_48;
wire n_64_49;
wire n_64_50;
wire n_64_51;
wire n_64_52;
wire n_64_53;
wire n_64_54;
wire n_64_55;
wire n_64_56;
wire n_64_57;
wire n_64_58;
wire n_64_59;
wire n_64_60;
wire n_64_61;
wire n_64_62;
wire n_64_63;
wire n_64_64;
wire n_64_65;
wire n_64_66;
wire n_64_67;
wire n_64_68;
wire n_64_69;
wire n_64_70;
wire n_64_71;
wire n_64_72;
wire n_64_73;
wire n_64_74;
wire n_64_75;
wire n_64_76;
wire n_64_77;
wire n_64_78;
wire n_64_79;
wire n_64_80;
wire n_64_81;
wire n_64_82;
wire n_64_83;
wire n_64_84;
wire n_64_85;
wire n_64_86;
wire n_64_87;
wire n_64_88;
wire n_64_89;
wire n_64_90;
wire n_64_91;
wire n_64_92;
wire n_64_93;
wire n_64_94;
wire n_64_95;
wire n_64_96;
wire n_64_97;
wire n_64_98;
wire n_64_99;
wire n_64_100;
wire n_64_101;
wire n_64_102;
wire n_64_103;
wire n_64_104;
wire n_64_105;
wire n_64_106;
wire n_64_107;
wire n_64_108;
wire n_64_109;
wire n_64_110;
wire n_64_111;
wire n_64_112;
wire n_64_113;
wire n_64_114;
wire n_64_115;
wire n_64_116;
wire n_64_117;
wire n_64_118;
wire n_64_119;
wire n_64_120;
wire n_64_121;
wire n_64_122;
wire n_64_123;
wire n_64_124;
wire n_64_125;
wire n_64_126;
wire n_64_127;
wire n_64_128;
wire n_64_129;
wire n_64_130;
wire n_64_131;
wire n_64_132;
wire n_64_133;
wire n_64_134;
wire n_64_135;
wire n_64_136;
wire n_64_137;
wire n_64_138;
wire n_64_139;
wire n_64_140;
wire n_64_141;
wire n_64_142;
wire n_64_143;
wire n_64_144;
wire n_64_145;
wire n_64_146;
wire n_64_147;
wire n_64_148;
wire n_64_149;
wire n_64_150;
wire n_64_151;
wire n_64_152;
wire n_64_153;
wire n_64_154;
wire n_64_155;
wire n_64_156;
wire n_64_157;
wire n_64_158;
wire n_64_159;
wire n_64_160;
wire n_64_161;
wire n_64_162;
wire n_64_163;
wire n_64_164;
wire n_64_165;
wire n_64_166;
wire n_64_167;
wire n_64_168;
wire n_64_169;
wire n_64_170;
wire n_64_171;
wire n_64_172;
wire n_64_173;
wire n_64_174;
wire n_64_175;
wire n_64_176;
wire n_64_177;
wire n_64_178;
wire n_64_179;
wire n_64_180;
wire n_64_181;
wire n_64_182;
wire n_64_183;
wire n_64_184;
wire n_64_185;
wire n_64_186;
wire n_64_187;
wire n_64_188;
wire n_64_189;
wire n_64_190;
wire n_64_191;
wire n_64_192;
wire \A[31] ;
wire \A[29] ;
wire \A[28] ;
wire \A[27] ;
wire \A[26] ;
wire \A[25] ;
wire \A[24] ;
wire \A[23] ;
wire \A[22] ;
wire \A[21] ;
wire \A[20] ;
wire \A[19] ;
wire \A[18] ;
wire \A[17] ;
wire \A[16] ;
wire \A[15] ;
wire \A[14] ;
wire \A[13] ;
wire \A[12] ;
wire \A[11] ;
wire \A[10] ;
wire \A[9] ;
wire \A[8] ;
wire \A[7] ;
wire \A[6] ;
wire \A[5] ;
wire \A[4] ;
wire \A[3] ;
wire \A[2] ;
wire \A[1] ;
wire \A[0] ;
wire \SC[6] ;
wire \SC[5] ;
wire \SC[4] ;
wire \SC[3] ;
wire \SC[2] ;
wire \SC[1] ;
wire \SC[0] ;
wire \multiplicand[31] ;
wire \multiplicand[30] ;
wire \multiplicand[29] ;
wire \multiplicand[28] ;
wire \multiplicand[27] ;
wire \multiplicand[26] ;
wire \multiplicand[25] ;
wire \multiplicand[24] ;
wire \multiplicand[23] ;
wire \multiplicand[22] ;
wire \multiplicand[21] ;
wire \multiplicand[20] ;
wire \multiplicand[19] ;
wire \multiplicand[18] ;
wire \multiplicand[17] ;
wire \multiplicand[16] ;
wire \multiplicand[15] ;
wire \multiplicand[14] ;
wire \multiplicand[13] ;
wire \multiplicand[12] ;
wire \multiplicand[11] ;
wire \multiplicand[10] ;
wire \multiplicand[9] ;
wire \multiplicand[8] ;
wire \multiplicand[7] ;
wire \multiplicand[6] ;
wire \multiplicand[5] ;
wire \multiplicand[4] ;
wire \multiplicand[3] ;
wire \multiplicand[2] ;
wire \multiplicand[1] ;
wire \multiplicand[0] ;
wire \Q[32] ;
wire \Q[31] ;
wire \Q[30] ;
wire \Q[29] ;
wire \Q[28] ;
wire \Q[27] ;
wire \Q[26] ;
wire \Q[25] ;
wire \Q[24] ;
wire \Q[23] ;
wire \Q[22] ;
wire \Q[21] ;
wire \Q[20] ;
wire \Q[19] ;
wire \Q[18] ;
wire \Q[17] ;
wire \Q[16] ;
wire \Q[15] ;
wire \Q[14] ;
wire \Q[13] ;
wire \Q[12] ;
wire \Q[11] ;
wire \Q[10] ;
wire \Q[9] ;
wire \Q[8] ;
wire \Q[7] ;
wire \Q[6] ;
wire \Q[5] ;
wire \Q[4] ;
wire \Q[3] ;
wire \Q[2] ;
wire \Q[1] ;
wire \Q[0] ;
wire out_sign;
wire CLOCK_slh__n427;
wire CTS_n_tid1_109;
wire n_64_1_5;
wire n_64_1_0;
wire n_64_1_6;
wire n_64_1_1;
wire n_64_1_7;
wire n_64_1_2;
wire n_64_1_8;
wire n_64_1_3;
wire n_64_1_9;
wire n_64_1_4;
wire n_64_193;
wire n_64_194;
wire n_64_195;
wire n_64_196;
wire n_64_197;
wire n_64_198;
wire n_64_199;
wire n_64_1_10;
wire n_64_1_11;
wire n_64_1_12;
wire n_64_200;
wire n_64_1_13;
wire n_64_1_14;
wire n_64_1_15;
wire n_64_201;
wire n_64_1_16;
wire n_64_202;
wire n_64_1_17;
wire n_64_203;
wire n_64_1_18;
wire n_64_204;
wire n_64_1_19;
wire n_64_205;
wire n_64_1_20;
wire n_64_206;
wire n_64_1_21;
wire n_64_207;
wire n_64_1_22;
wire n_64_208;
wire n_64_1_23;
wire n_64_209;
wire n_64_1_24;
wire n_64_210;
wire n_64_1_25;
wire n_64_211;
wire n_64_1_26;
wire n_64_212;
wire n_64_1_27;
wire n_64_213;
wire n_64_1_28;
wire n_64_214;
wire n_64_1_29;
wire n_64_215;
wire n_64_1_30;
wire n_64_216;
wire n_64_1_31;
wire n_64_217;
wire n_64_1_32;
wire n_64_218;
wire n_64_1_33;
wire n_64_219;
wire n_64_1_34;
wire n_64_220;
wire n_64_1_35;
wire n_64_221;
wire n_64_1_36;
wire n_64_222;
wire n_64_1_37;
wire n_64_223;
wire n_64_1_38;
wire n_64_224;
wire n_64_1_39;
wire n_64_225;
wire n_64_1_40;
wire n_64_226;
wire n_64_1_41;
wire n_64_227;
wire n_64_1_42;
wire n_64_228;
wire n_64_1_43;
wire n_64_229;
wire n_64_1_44;
wire n_64_230;
wire n_64_1_45;
wire n_64_231;
wire n_64_1_46;
wire n_64_232;
wire n_64_1_47;
wire n_64_233;
wire n_64_1_48;
wire n_64_234;
wire n_64_1_49;
wire n_64_235;
wire n_64_1_50;
wire n_64_236;
wire n_64_1_51;
wire n_64_237;
wire n_64_1_52;
wire n_64_238;
wire n_64_1_53;
wire n_64_239;
wire n_64_1_54;
wire n_64_240;
wire n_64_1_55;
wire n_64_241;
wire n_64_1_56;
wire n_64_242;
wire n_64_1_57;
wire n_64_243;
wire n_64_1_58;
wire n_64_244;
wire n_64_1_59;
wire n_64_245;
wire n_64_1_60;
wire n_64_246;
wire n_64_1_61;
wire n_64_247;
wire n_64_1_62;
wire n_64_248;
wire n_64_1_63;
wire n_64_249;
wire n_64_1_64;
wire n_64_250;
wire n_64_1_65;
wire n_64_251;
wire n_64_1_66;
wire n_64_252;
wire n_64_1_67;
wire n_64_253;
wire n_64_1_68;
wire n_64_254;
wire n_64_1_69;
wire n_64_255;
wire n_64_1_70;
wire n_64_256;
wire n_64_1_71;
wire n_64_257;
wire n_64_1_72;
wire n_64_258;
wire n_64_1_73;
wire n_64_259;
wire n_64_1_74;
wire n_64_260;
wire n_64_1_75;
wire n_64_265;
wire n_64_266;
wire n_64_267;
wire n_64_268;
wire n_64_269;
wire n_64_270;
wire n_64_271;
wire n_64_272;
wire n_64_273;
wire n_64_274;
wire n_64_275;
wire n_64_276;
wire n_64_277;
wire n_64_278;
wire n_64_279;
wire n_64_280;
wire n_64_281;
wire n_64_282;
wire n_64_283;
wire n_64_284;
wire n_64_285;
wire n_64_286;
wire n_64_287;
wire n_64_288;
wire n_64_289;
wire n_64_290;
wire n_64_291;
wire n_64_292;
wire n_64_293;
wire n_64_294;
wire n_64_295;
wire n_64_296;
wire n_64_300;
wire n_64_1_81;
wire n_64_301;
wire n_64_1_82;
wire n_64_302;
wire n_64_1_83;
wire n_64_303;
wire n_64_1_84;
wire n_64_310;
wire n_64_1_91;
wire n_64_311;
wire n_64_1_92;
wire n_64_312;
wire n_64_1_93;
wire n_64_313;
wire n_64_1_94;
wire n_64_314;
wire n_64_1_95;
wire n_64_315;
wire n_64_1_96;
wire n_64_316;
wire n_64_1_97;
wire n_64_317;
wire n_64_1_98;
wire n_64_318;
wire n_64_1_99;
wire n_64_319;
wire n_64_1_100;
wire n_64_320;
wire n_64_1_101;
wire n_64_321;
wire n_64_1_102;
wire n_64_322;
wire n_64_1_103;
wire n_64_323;
wire n_64_1_104;
wire n_64_324;
wire n_64_1_105;
wire n_64_325;
wire n_64_1_106;
wire n_64_326;
wire n_64_1_107;
wire n_64_327;
wire n_64_1_108;
wire n_64_328;
wire n_64_1_110;
wire n_64_1_111;
wire n_64_329;
wire n_64_1_113;
wire n_64_330;
wire n_64_1_114;
wire n_64_331;
wire n_64_1_115;
wire n_64_332;
wire n_64_1_116;
wire n_64_333;
wire n_64_1_117;
wire n_64_334;
wire n_64_1_118;
wire n_64_335;
wire n_64_1_119;
wire n_64_336;
wire n_64_1_120;
wire n_64_337;
wire n_64_1_121;
wire n_64_338;
wire n_64_1_122;
wire n_64_339;
wire n_64_1_123;
wire n_64_340;
wire n_64_1_124;
wire n_64_341;
wire n_64_1_125;
wire n_64_342;
wire n_64_1_126;
wire n_64_343;
wire n_64_1_127;
wire n_64_344;
wire n_64_1_128;
wire n_64_345;
wire n_64_1_129;
wire n_64_346;
wire n_64_1_130;
wire n_64_347;
wire n_64_1_131;
wire n_64_348;
wire n_64_1_132;
wire n_64_349;
wire n_64_1_133;
wire n_64_350;
wire n_64_1_134;
wire n_64_351;
wire n_64_1_135;
wire n_64_352;
wire n_64_1_136;
wire n_64_353;
wire n_64_1_137;
wire n_64_354;
wire n_64_1_138;
wire n_64_355;
wire n_64_1_139;
wire n_64_356;
wire n_64_1_140;
wire n_64_357;
wire n_64_1_141;
wire n_64_358;
wire n_64_1_142;
wire n_64_359;
wire hfn_ipo_n19;
wire n_64_1_145;
wire n_64_1_146;
wire n_64_1_147;
wire n_64_1_148;
wire n_64_297;
wire n_64_1_149;
wire n_64_361;
wire n_64_1_150;
wire n_64_362;
wire n_64_1_151;
wire n_64_363;
wire n_64_1_152;
wire n_64_364;
wire n_64_1_153;
wire n_64_365;
wire n_64_1_154;
wire n_64_366;
wire n_64_1_155;
wire n_64_367;
wire n_64_1_156;
wire n_64_368;
wire n_64_1_157;
wire n_64_369;
wire n_64_1_158;
wire n_64_370;
wire n_64_1_159;
wire n_64_371;
wire n_64_1_160;
wire n_64_372;
wire n_64_1_161;
wire n_64_373;
wire n_64_1_162;
wire n_64_374;
wire n_64_1_163;
wire n_64_375;
wire n_64_1_164;
wire n_64_376;
wire n_64_1_165;
wire n_64_377;
wire n_64_1_166;
wire n_64_378;
wire n_64_1_167;
wire n_64_379;
wire n_64_1_168;
wire n_64_380;
wire n_64_1_169;
wire n_64_381;
wire n_64_1_170;
wire n_64_382;
wire n_64_1_171;
wire n_64_383;
wire n_64_1_172;
wire n_64_384;
wire n_64_1_173;
wire n_64_385;
wire n_64_1_174;
wire n_64_386;
wire n_64_1_175;
wire n_64_387;
wire n_64_1_176;
wire n_64_388;
wire n_64_1_177;
wire n_64_389;
wire n_64_1_178;
wire n_64_390;
wire n_64_1_179;
wire n_64_391;
wire n_64_1_180;
wire n_64_1_181;
wire n_64_392;
wire n_64_1_182;
wire n_64_1_183;
wire n_64_1_186;
wire n_64_1_187;
wire n_64_393;
wire n_64_394;
wire n_64_1_188;
wire n_64_1_189;
wire n_64_1_190;
wire n_64_1_191;
wire n_64_1_192;
wire n_64_264;
wire n_64_1_193;
wire n_64_1_194;
wire n_64_1_144;
wire n_64_261;
wire n_64_1_143;
wire n_64_1_76;
wire n_64_262;
wire n_64_1_77;
wire n_64_1_79;
wire n_64_1_195;
wire n_64_1_196;
wire n_64_1_197;
wire n_64_1_198;
wire n_64_1_199;
wire n_64_1_200;
wire n_64_263;
wire n_64_1_201;
wire n_64_1_78;
wire n_64_1_202;
wire n_64_298;
wire n_64_1_203;
wire n_64_1_204;
wire n_64_299;
wire n_64_1_80;
wire n_64_1_205;
wire n_64_304;
wire n_64_1_85;
wire n_64_1_206;
wire n_64_305;
wire n_64_1_86;
wire n_64_1_207;
wire n_64_306;
wire n_64_1_87;
wire n_64_1_208;
wire n_64_307;
wire n_64_1_88;
wire n_64_1_209;
wire n_64_308;
wire n_64_1_89;
wire n_64_1_210;
wire n_64_309;
wire n_64_1_90;
wire n_64_1_211;
wire n_64_1_109;
wire n_64_1_212;
wire n_64_1_112;
wire n_64_1_184;
wire n_64_1_185;
wire n_64;
wire n_0;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire hfn_ipo_n20;
wire hfn_ipo_n21;
wire drc_ipo_n22;
wire CTS_n_tid1_111;
wire CTS_n_tid0_338;
wire hfn_ipo_n17;
wire hfn_ipo_n18;
wire drc_ipo_n24;
wire drc_ipo_n25;
wire drc_ipo_n26;
wire drc_ipo_n27;
wire drc_ipo_n28;
wire drc_ipo_n29;
wire drc_ipo_n30;
wire drc_ipo_n31;
wire drc_ipo_n32;
wire drc_ipo_n33;
wire drc_ipo_n34;
wire drc_ipo_n35;
wire drc_ipo_n36;
wire drc_ipo_n37;
wire drc_ipo_n38;
wire drc_ipo_n39;
wire drc_ipo_n40;
wire drc_ipo_n41;
wire drc_ipo_n42;
wire drc_ipo_n43;
wire drc_ipo_n44;
wire drc_ipo_n45;
wire drc_ipo_n46;
wire drc_ipo_n47;
wire drc_ipo_n48;
wire drc_ipo_n49;
wire drc_ipo_n50;
wire drc_ipo_n51;
wire drc_ipo_n52;
wire drc_ipo_n53;
wire drc_ipo_n54;
wire drc_ipo_n55;
wire drc_ipo_n56;
wire drc_ipo_n57;
wire drc_ipo_n58;
wire drc_ipo_n59;
wire drc_ipo_n60;
wire drc_ipo_n61;
wire drc_ipo_n62;
wire drc_ipo_n63;
wire drc_ipo_n64;
wire drc_ipo_n65;
wire drc_ipo_n66;
wire drc_ipo_n67;
wire drc_ipo_n68;
wire drc_ipo_n69;
wire drc_ipo_n70;
wire drc_ipo_n71;
wire drc_ipo_n72;
wire drc_ipo_n73;
wire drc_ipo_n74;
wire drc_ipo_n75;
wire drc_ipo_n76;
wire drc_ipo_n77;
wire drc_ipo_n78;
wire drc_ipo_n79;
wire drc_ipo_n80;
wire drc_ipo_n81;
wire drc_ipo_n82;
wire drc_ipo_n83;
wire drc_ipo_n84;
wire drc_ipo_n85;
wire drc_ipo_n86;
wire drc_ipo_n87;
wire drc_ipo_n88;
wire drc_ipo_n89;
wire CTS_n_tid0_339;
wire CTS_n_tid1_244;
wire CTS_n_tid0_337;
wire CTS_n_tid0_234;
wire CLOCK_slh__n439;
wire CTS_n_tid0_128;
wire CLOCK_slh__n428;
wire CLOCK_slh__n440;
wire CLOCK_slh__n443;
wire CTS_n_tid0_136;
wire CLOCK_slh__n444;
wire CLOCK_slh__n447;
wire CLOCK_slh__n448;
wire CLOCK_slh__n431;
wire CLOCK_slh__n432;
wire CLOCK_slh__n435;
wire CLOCK_slh__n436;
wire CLOCK_slh__n451;
wire CLOCK_slh__n452;
wire CLOCK_slh__n455;
wire CLOCK_slh__n456;
wire CLOCK_slh__n459;
wire CLOCK_slh__n460;
wire CLOCK_slh__n463;
wire CLOCK_slh__n464;
wire CLOCK_slh__n467;
wire CLOCK_slh__n468;
wire CLOCK_slh__n471;
wire CLOCK_slh__n472;
wire CLOCK_slh__n475;
wire CLOCK_slh__n476;
wire CLOCK_slh__n479;
wire CLOCK_slh__n480;
wire CLOCK_slh__n483;
wire CLOCK_slh__n484;
wire CLOCK_slh__n487;
wire CLOCK_slh__n488;
wire CLOCK_slh__n491;
wire CLOCK_slh__n492;
wire CLOCK_slh__n495;
wire CLOCK_slh__n496;
wire CLOCK_slh__n499;
wire CLOCK_slh__n500;
wire CLOCK_slh__n503;
wire CLOCK_slh__n504;
wire CLOCK_slh__n507;
wire CLOCK_slh__n508;
wire CLOCK_slh__n511;
wire CLOCK_slh__n513;
wire CLOCK_slh__n515;
wire CLOCK_slh__n517;
wire CLOCK_slh__n519;
wire CLOCK_slh__n520;
wire CLOCK_slh__n521;
wire CLOCK_slh__n522;


NAND2_X4 i_64_1_409 (.ZN (n_64_1_185), .A1 (n_64_1_186), .A2 (n_64_1_187));
INV_X4 i_64_1_408 (.ZN (n_64_1_184), .A (n_64_1_185));
NAND2_X2 i_64_1_407 (.ZN (n_64_1_112), .A1 (n_64_1_184), .A2 (drc_ipo_n55));
NOR2_X1 i_64_1_406 (.ZN (n_64_1_212), .A1 (drc_ipo_n55), .A2 (n_64_1_185));
INV_X2 i_64_1_405 (.ZN (n_64_1_109), .A (n_64_1_212));
OR2_X1 i_64_1_404 (.ZN (n_64_1_211), .A1 (n_64_1_109), .A2 (drc_ipo_n36));
OAI221_X1 i_64_1_403 (.ZN (n_64_1_90), .A (n_64_1_211), .B1 (\Q[13] ), .B2 (n_64_1_184)
    , .C1 (n_64_110), .C2 (n_64_1_112));
INV_X1 i_64_1_402 (.ZN (n_64_309), .A (n_64_1_90));
OR2_X1 i_64_1_401 (.ZN (n_64_1_210), .A1 (n_64_1_109), .A2 (drc_ipo_n35));
OAI221_X1 i_64_1_400 (.ZN (n_64_1_89), .A (n_64_1_210), .B1 (\Q[12] ), .B2 (n_64_1_184)
    , .C1 (n_64_109), .C2 (n_64_1_112));
INV_X1 i_64_1_399 (.ZN (n_64_308), .A (n_64_1_89));
OR2_X1 i_64_1_398 (.ZN (n_64_1_209), .A1 (n_64_1_109), .A2 (drc_ipo_n34));
OAI221_X1 i_64_1_397 (.ZN (n_64_1_88), .A (n_64_1_209), .B1 (\Q[11] ), .B2 (n_64_1_184)
    , .C1 (n_64_108), .C2 (n_64_1_112));
INV_X1 i_64_1_396 (.ZN (n_64_307), .A (n_64_1_88));
OR2_X1 i_64_1_395 (.ZN (n_64_1_208), .A1 (n_64_1_109), .A2 (drc_ipo_n33));
OAI221_X1 i_64_1_394 (.ZN (n_64_1_87), .A (n_64_1_208), .B1 (\Q[10] ), .B2 (n_64_1_184)
    , .C1 (n_64_107), .C2 (n_64_1_112));
INV_X1 i_64_1_393 (.ZN (n_64_306), .A (n_64_1_87));
OR2_X1 i_64_1_392 (.ZN (n_64_1_207), .A1 (n_64_1_109), .A2 (drc_ipo_n32));
OAI221_X1 i_64_1_379 (.ZN (n_64_1_86), .A (n_64_1_207), .B1 (\Q[9] ), .B2 (n_64_1_184)
    , .C1 (n_64_106), .C2 (n_64_1_112));
INV_X1 i_64_1_378 (.ZN (n_64_305), .A (n_64_1_86));
OR2_X1 i_64_1_305 (.ZN (n_64_1_206), .A1 (n_64_1_109), .A2 (drc_ipo_n31));
OAI221_X1 i_64_1_303 (.ZN (n_64_1_85), .A (n_64_1_206), .B1 (\Q[8] ), .B2 (n_64_1_184)
    , .C1 (n_64_105), .C2 (n_64_1_112));
INV_X1 i_64_1_241 (.ZN (n_64_304), .A (n_64_1_85));
OR2_X1 i_64_1_237 (.ZN (n_64_1_205), .A1 (n_64_1_109), .A2 (drc_ipo_n26));
OAI221_X1 i_64_1_200 (.ZN (n_64_1_80), .A (n_64_1_205), .B1 (\Q[3] ), .B2 (n_64_1_184)
    , .C1 (n_64_100), .C2 (n_64_1_112));
INV_X1 i_64_1_199 (.ZN (n_64_299), .A (n_64_1_80));
NOR2_X1 i_64_1_198 (.ZN (n_64_1_204), .A1 (n_64_99), .A2 (n_64_1_112));
OAI22_X1 i_64_1_197 (.ZN (n_64_1_203), .A1 (n_64_1_109), .A2 (drc_ipo_n25), .B1 (\Q[2] ), .B2 (n_64_1_184));
NOR2_X1 i_64_1_196 (.ZN (CLOCK_slh__n487), .A1 (n_64_1_204), .A2 (n_64_1_203));
NOR2_X1 i_64_1_195 (.ZN (n_64_1_202), .A1 (n_64_1_189), .A2 (out_sign));
INV_X1 i_64_1_194 (.ZN (n_64_1_78), .A (n_64_1_202));
NAND2_X1 i_64_1_193 (.ZN (n_64_1_201), .A1 (n_64_192), .A2 (hfn_ipo_n17));
INV_X1 i_64_1_192 (.ZN (n_64_263), .A (n_64_1_201));
NAND2_X1 i_64_1_191 (.ZN (n_64_1_200), .A1 (n_64_191), .A2 (hfn_ipo_n17));
INV_X1 i_64_1_190 (.ZN (n_64_1_199), .A (n_64_66));
INV_X1 i_64_1_189 (.ZN (n_64_1_198), .A (n_64_98));
INV_X1 i_64_1_180 (.ZN (n_64_1_197), .A (drc_ipo_n22));
INV_X1 i_64_1_179 (.ZN (n_64_1_196), .A (n_64_1_148));
INV_X1 i_64_1_178 (.ZN (n_64_1_195), .A (n_64_1_145));
OAI221_X1 i_64_1_177 (.ZN (n_64_1_79), .A (n_64_1_195), .B1 (n_64_1_199), .B2 (n_64_1_196)
    , .C1 (n_64_1_198), .C2 (n_64_1_197));
NAND2_X1 i_64_1_144 (.ZN (n_64_1_77), .A1 (n_64_1_79), .A2 (n_64_1_202));
NAND2_X1 i_64_1_143 (.ZN (n_64_262), .A1 (n_64_1_200), .A2 (n_64_1_77));
NAND2_X1 i_64_1_142 (.ZN (n_64_1_76), .A1 (n_64_190), .A2 (hfn_ipo_n17));
AOI221_X1 i_64_1_141 (.ZN (n_64_1_143), .A (n_64_1_145), .B1 (n_64_65), .B2 (n_64_1_148)
    , .C1 (n_64_97), .C2 (drc_ipo_n22));
OAI21_X1 i_64_1_140 (.ZN (n_64_261), .A (n_64_1_76), .B1 (hfn_ipo_n18), .B2 (n_64_1_143));
INV_X1 i_64_1_139 (.ZN (n_64_1_144), .A (n_64_1_79));
INV_X1 i_64_1_391 (.ZN (n_64_1_194), .A (drc_ipo_n88));
INV_X1 i_64_1_390 (.ZN (n_64_1_193), .A (\Q[0] ));
NOR2_X1 i_64_1_389 (.ZN (n_64_264), .A1 (drc_ipo_n89), .A2 (n_64_1_194));
NAND3_X1 i_64_1_388 (.ZN (n_64_1_192), .A1 (\SC[2] ), .A2 (\SC[1] ), .A3 (\SC[0] ));
NAND2_X1 i_64_1_387 (.ZN (n_64_1_191), .A1 (\SC[4] ), .A2 (\SC[3] ));
NOR4_X1 i_64_1_386 (.ZN (n_64_1_190), .A1 (\SC[6] ), .A2 (\SC[5] ), .A3 (n_64_1_191), .A4 (n_64_1_192));
INV_X1 i_64_1_385 (.ZN (n_64_1_189), .A (n_64_1_190));
OAI21_X1 i_64_1_384 (.ZN (n_64_1_188), .A (n_64_264), .B1 (n_64_3), .B2 (n_64_1_190));
INV_X1 i_64_1_383 (.ZN (n_64_394), .A (n_64_1_188));
NAND2_X1 i_64_1_382 (.ZN (n_64_393), .A1 (n_64_264), .A2 (n_64_1_189));
NOR3_X1 i_64_1_381 (.ZN (n_64_1_187), .A1 (\SC[2] ), .A2 (\SC[1] ), .A3 (\SC[0] ));
NOR4_X1 i_64_1_380 (.ZN (n_64_1_186), .A1 (\SC[6] ), .A2 (\SC[5] ), .A3 (\SC[4] ), .A4 (\SC[3] ));
AND2_X4 i_64_1_377 (.ZN (n_64_1_183), .A1 (drc_ipo_n87), .A2 (n_64_1_184));
AOI22_X1 i_64_1_376 (.ZN (n_64_1_182), .A1 (\multiplicand[31] ), .A2 (n_64_1_185)
    , .B1 (n_64_34), .B2 (n_64_1_183));
INV_X1 i_64_1_375 (.ZN (n_64_392), .A (n_64_1_182));
NOR2_X4 i_64_1_374 (.ZN (n_64_1_181), .A1 (drc_ipo_n87), .A2 (n_64_1_185));
AOI222_X1 i_64_1_373 (.ZN (n_64_1_180), .A1 (drc_ipo_n86), .A2 (n_64_1_181), .B1 (\multiplicand[30] )
    , .B2 (n_64_1_185), .C1 (n_64_33), .C2 (n_64_1_183));
INV_X1 i_64_1_372 (.ZN (n_64_391), .A (n_64_1_180));
AOI222_X1 i_64_1_371 (.ZN (n_64_1_179), .A1 (drc_ipo_n85), .A2 (n_64_1_181), .B1 (\multiplicand[29] )
    , .B2 (n_64_1_185), .C1 (n_64_32), .C2 (n_64_1_183));
INV_X1 i_64_1_370 (.ZN (n_64_390), .A (n_64_1_179));
AOI222_X1 i_64_1_369 (.ZN (n_64_1_178), .A1 (drc_ipo_n84), .A2 (n_64_1_181), .B1 (\multiplicand[28] )
    , .B2 (n_64_1_185), .C1 (n_64_31), .C2 (n_64_1_183));
INV_X1 i_64_1_368 (.ZN (n_64_389), .A (n_64_1_178));
AOI222_X1 i_64_1_367 (.ZN (n_64_1_177), .A1 (drc_ipo_n83), .A2 (n_64_1_181), .B1 (\multiplicand[27] )
    , .B2 (n_64_1_185), .C1 (n_64_30), .C2 (n_64_1_183));
INV_X1 i_64_1_366 (.ZN (n_64_388), .A (n_64_1_177));
AOI222_X1 i_64_1_365 (.ZN (n_64_1_176), .A1 (drc_ipo_n82), .A2 (n_64_1_181), .B1 (\multiplicand[26] )
    , .B2 (n_64_1_185), .C1 (n_64_29), .C2 (n_64_1_183));
INV_X1 i_64_1_364 (.ZN (n_64_387), .A (n_64_1_176));
AOI222_X1 i_64_1_363 (.ZN (n_64_1_175), .A1 (drc_ipo_n81), .A2 (n_64_1_181), .B1 (\multiplicand[25] )
    , .B2 (n_64_1_185), .C1 (n_64_28), .C2 (n_64_1_183));
INV_X1 i_64_1_362 (.ZN (n_64_386), .A (n_64_1_175));
AOI222_X1 i_64_1_361 (.ZN (n_64_1_174), .A1 (drc_ipo_n80), .A2 (n_64_1_181), .B1 (\multiplicand[24] )
    , .B2 (n_64_1_185), .C1 (n_64_27), .C2 (n_64_1_183));
INV_X1 i_64_1_360 (.ZN (n_64_385), .A (n_64_1_174));
AOI222_X1 i_64_1_359 (.ZN (n_64_1_173), .A1 (drc_ipo_n79), .A2 (n_64_1_181), .B1 (\multiplicand[23] )
    , .B2 (n_64_1_185), .C1 (n_64_26), .C2 (n_64_1_183));
INV_X1 i_64_1_358 (.ZN (n_64_384), .A (n_64_1_173));
AOI222_X1 i_64_1_357 (.ZN (n_64_1_172), .A1 (drc_ipo_n78), .A2 (n_64_1_181), .B1 (\multiplicand[22] )
    , .B2 (n_64_1_185), .C1 (n_64_25), .C2 (n_64_1_183));
INV_X1 i_64_1_356 (.ZN (n_64_383), .A (n_64_1_172));
AOI222_X1 i_64_1_355 (.ZN (n_64_1_171), .A1 (drc_ipo_n77), .A2 (n_64_1_181), .B1 (\multiplicand[21] )
    , .B2 (n_64_1_185), .C1 (n_64_24), .C2 (n_64_1_183));
INV_X1 i_64_1_354 (.ZN (n_64_382), .A (n_64_1_171));
AOI222_X1 i_64_1_353 (.ZN (n_64_1_170), .A1 (drc_ipo_n76), .A2 (n_64_1_181), .B1 (\multiplicand[20] )
    , .B2 (n_64_1_185), .C1 (n_64_23), .C2 (n_64_1_183));
INV_X1 i_64_1_352 (.ZN (n_64_381), .A (n_64_1_170));
AOI222_X1 i_64_1_351 (.ZN (n_64_1_169), .A1 (drc_ipo_n75), .A2 (n_64_1_181), .B1 (\multiplicand[19] )
    , .B2 (n_64_1_185), .C1 (n_64_22), .C2 (n_64_1_183));
INV_X1 i_64_1_350 (.ZN (n_64_380), .A (n_64_1_169));
AOI222_X1 i_64_1_349 (.ZN (n_64_1_168), .A1 (drc_ipo_n74), .A2 (n_64_1_181), .B1 (\multiplicand[18] )
    , .B2 (n_64_1_185), .C1 (n_64_21), .C2 (n_64_1_183));
INV_X1 i_64_1_348 (.ZN (n_64_379), .A (n_64_1_168));
AOI222_X1 i_64_1_347 (.ZN (n_64_1_167), .A1 (drc_ipo_n73), .A2 (n_64_1_181), .B1 (\multiplicand[17] )
    , .B2 (n_64_1_185), .C1 (n_64_20), .C2 (n_64_1_183));
INV_X1 i_64_1_346 (.ZN (n_64_378), .A (n_64_1_167));
AOI222_X1 i_64_1_345 (.ZN (n_64_1_166), .A1 (drc_ipo_n72), .A2 (n_64_1_181), .B1 (\multiplicand[16] )
    , .B2 (n_64_1_185), .C1 (n_64_19), .C2 (n_64_1_183));
INV_X1 i_64_1_344 (.ZN (n_64_377), .A (n_64_1_166));
AOI222_X1 i_64_1_343 (.ZN (n_64_1_165), .A1 (drc_ipo_n71), .A2 (n_64_1_181), .B1 (\multiplicand[15] )
    , .B2 (n_64_1_185), .C1 (n_64_18), .C2 (n_64_1_183));
INV_X1 i_64_1_342 (.ZN (n_64_376), .A (n_64_1_165));
AOI222_X1 i_64_1_341 (.ZN (n_64_1_164), .A1 (drc_ipo_n70), .A2 (n_64_1_181), .B1 (\multiplicand[14] )
    , .B2 (n_64_1_185), .C1 (n_64_17), .C2 (n_64_1_183));
INV_X1 i_64_1_340 (.ZN (n_64_375), .A (n_64_1_164));
AOI222_X1 i_64_1_339 (.ZN (n_64_1_163), .A1 (drc_ipo_n69), .A2 (n_64_1_181), .B1 (\multiplicand[13] )
    , .B2 (n_64_1_185), .C1 (n_64_16), .C2 (n_64_1_183));
INV_X1 i_64_1_338 (.ZN (n_64_374), .A (n_64_1_163));
AOI222_X1 i_64_1_337 (.ZN (n_64_1_162), .A1 (drc_ipo_n68), .A2 (n_64_1_181), .B1 (\multiplicand[12] )
    , .B2 (n_64_1_185), .C1 (n_64_15), .C2 (n_64_1_183));
INV_X1 i_64_1_336 (.ZN (n_64_373), .A (n_64_1_162));
AOI222_X1 i_64_1_335 (.ZN (n_64_1_161), .A1 (drc_ipo_n67), .A2 (n_64_1_181), .B1 (\multiplicand[11] )
    , .B2 (n_64_1_185), .C1 (n_64_14), .C2 (n_64_1_183));
INV_X1 i_64_1_334 (.ZN (n_64_372), .A (n_64_1_161));
AOI222_X1 i_64_1_333 (.ZN (n_64_1_160), .A1 (drc_ipo_n66), .A2 (n_64_1_181), .B1 (\multiplicand[10] )
    , .B2 (n_64_1_185), .C1 (n_64_13), .C2 (n_64_1_183));
INV_X1 i_64_1_332 (.ZN (n_64_371), .A (n_64_1_160));
AOI222_X1 i_64_1_331 (.ZN (n_64_1_159), .A1 (drc_ipo_n65), .A2 (n_64_1_181), .B1 (\multiplicand[9] )
    , .B2 (n_64_1_185), .C1 (n_64_12), .C2 (n_64_1_183));
INV_X1 i_64_1_330 (.ZN (n_64_370), .A (n_64_1_159));
AOI222_X1 i_64_1_329 (.ZN (n_64_1_158), .A1 (drc_ipo_n64), .A2 (n_64_1_181), .B1 (\multiplicand[8] )
    , .B2 (n_64_1_185), .C1 (n_64_11), .C2 (n_64_1_183));
INV_X1 i_64_1_328 (.ZN (n_64_369), .A (n_64_1_158));
AOI222_X1 i_64_1_327 (.ZN (n_64_1_157), .A1 (drc_ipo_n63), .A2 (n_64_1_181), .B1 (\multiplicand[7] )
    , .B2 (n_64_1_185), .C1 (n_64_10), .C2 (n_64_1_183));
INV_X1 i_64_1_326 (.ZN (n_64_368), .A (n_64_1_157));
AOI222_X1 i_64_1_325 (.ZN (n_64_1_156), .A1 (drc_ipo_n62), .A2 (n_64_1_181), .B1 (\multiplicand[6] )
    , .B2 (n_64_1_185), .C1 (n_64_9), .C2 (n_64_1_183));
INV_X1 i_64_1_324 (.ZN (n_64_367), .A (n_64_1_156));
AOI222_X1 i_64_1_323 (.ZN (n_64_1_155), .A1 (drc_ipo_n61), .A2 (n_64_1_181), .B1 (\multiplicand[5] )
    , .B2 (n_64_1_185), .C1 (n_64_8), .C2 (n_64_1_183));
INV_X1 i_64_1_322 (.ZN (n_64_366), .A (n_64_1_155));
AOI222_X1 i_64_1_321 (.ZN (n_64_1_154), .A1 (drc_ipo_n60), .A2 (n_64_1_181), .B1 (\multiplicand[4] )
    , .B2 (n_64_1_185), .C1 (n_64_7), .C2 (n_64_1_183));
INV_X1 i_64_1_320 (.ZN (n_64_365), .A (n_64_1_154));
AOI222_X1 i_64_1_319 (.ZN (n_64_1_153), .A1 (drc_ipo_n59), .A2 (n_64_1_181), .B1 (\multiplicand[3] )
    , .B2 (n_64_1_185), .C1 (n_64_6), .C2 (n_64_1_183));
INV_X1 i_64_1_318 (.ZN (n_64_364), .A (n_64_1_153));
AOI222_X1 i_64_1_317 (.ZN (n_64_1_152), .A1 (drc_ipo_n58), .A2 (n_64_1_181), .B1 (\multiplicand[2] )
    , .B2 (n_64_1_185), .C1 (n_64_5), .C2 (n_64_1_183));
INV_X1 i_64_1_316 (.ZN (n_64_363), .A (n_64_1_152));
AOI222_X1 i_64_1_315 (.ZN (n_64_1_151), .A1 (drc_ipo_n57), .A2 (n_64_1_181), .B1 (\multiplicand[1] )
    , .B2 (n_64_1_185), .C1 (n_64_4), .C2 (n_64_1_183));
INV_X1 i_64_1_314 (.ZN (n_64_362), .A (n_64_1_151));
AOI22_X1 i_64_1_313 (.ZN (n_64_1_150), .A1 (\multiplicand[0] ), .A2 (n_64_1_185), .B1 (drc_ipo_n56), .B2 (n_64_1_184));
INV_X1 i_64_1_312 (.ZN (n_64_361), .A (n_64_1_150));
OAI22_X1 i_64_1_311 (.ZN (n_64_1_149), .A1 (\Q[1] ), .A2 (n_64_1_184), .B1 (drc_ipo_n24), .B2 (n_64_1_185));
INV_X1 i_64_1_310 (.ZN (n_64_297), .A (n_64_1_149));
AOI21_X4 i_64_1_309 (.ZN (n_64_1_148), .A (n_64_1_149), .B1 (\Q[0] ), .B2 (n_64_1_185));
NOR3_X1 i_64_1_308 (.ZN (n_64_1_147), .A1 (n_64_1_193), .A2 (n_64_1_184), .A3 (\Q[1] ));
NOR2_X4 i_64_1_307 (.ZN (n_64_1_146), .A1 (n_64_1_148), .A2 (drc_ipo_n22));
AND2_X1 i_64_1_306 (.ZN (n_64_1_145), .A1 (\A[31] ), .A2 (n_64_1_146));
BUF_X2 hfn_ipo_c19 (.Z (hfn_ipo_n19), .A (n_64_1_78));
INV_X1 i_64_1_302 (.ZN (n_64_359), .A (n_64_1_143));
AOI222_X1 i_64_1_301 (.ZN (n_64_1_142), .A1 (n_64_96), .A2 (drc_ipo_n22), .B1 (n_64_64)
    , .B2 (n_64_1_148), .C1 (\A[29] ), .C2 (n_64_1_146));
INV_X1 i_64_1_300 (.ZN (n_64_358), .A (n_64_1_142));
AOI222_X1 i_64_1_299 (.ZN (n_64_1_141), .A1 (n_64_95), .A2 (drc_ipo_n22), .B1 (n_64_63)
    , .B2 (n_64_1_148), .C1 (\A[28] ), .C2 (n_64_1_146));
INV_X1 i_64_1_298 (.ZN (n_64_357), .A (n_64_1_141));
AOI222_X1 i_64_1_297 (.ZN (n_64_1_140), .A1 (n_64_94), .A2 (drc_ipo_n22), .B1 (n_64_62)
    , .B2 (n_64_1_148), .C1 (\A[27] ), .C2 (n_64_1_146));
INV_X1 i_64_1_296 (.ZN (n_64_356), .A (n_64_1_140));
AOI222_X1 i_64_1_295 (.ZN (n_64_1_139), .A1 (n_64_93), .A2 (drc_ipo_n22), .B1 (n_64_61)
    , .B2 (n_64_1_148), .C1 (\A[26] ), .C2 (n_64_1_146));
INV_X1 i_64_1_294 (.ZN (n_64_355), .A (n_64_1_139));
AOI222_X1 i_64_1_293 (.ZN (n_64_1_138), .A1 (n_64_92), .A2 (drc_ipo_n22), .B1 (n_64_60)
    , .B2 (n_64_1_148), .C1 (\A[25] ), .C2 (n_64_1_146));
INV_X1 i_64_1_292 (.ZN (n_64_354), .A (n_64_1_138));
AOI222_X1 i_64_1_291 (.ZN (n_64_1_137), .A1 (n_64_91), .A2 (drc_ipo_n22), .B1 (n_64_59)
    , .B2 (n_64_1_148), .C1 (\A[24] ), .C2 (n_64_1_146));
INV_X1 i_64_1_290 (.ZN (n_64_353), .A (n_64_1_137));
AOI222_X1 i_64_1_289 (.ZN (n_64_1_136), .A1 (n_64_90), .A2 (drc_ipo_n22), .B1 (n_64_58)
    , .B2 (n_64_1_148), .C1 (\A[23] ), .C2 (n_64_1_146));
INV_X1 i_64_1_288 (.ZN (n_64_352), .A (n_64_1_136));
AOI222_X1 i_64_1_287 (.ZN (n_64_1_135), .A1 (n_64_89), .A2 (drc_ipo_n22), .B1 (n_64_57)
    , .B2 (n_64_1_148), .C1 (\A[22] ), .C2 (n_64_1_146));
INV_X1 i_64_1_286 (.ZN (n_64_351), .A (n_64_1_135));
AOI222_X1 i_64_1_285 (.ZN (n_64_1_134), .A1 (n_64_88), .A2 (drc_ipo_n22), .B1 (n_64_56)
    , .B2 (n_64_1_148), .C1 (\A[21] ), .C2 (n_64_1_146));
INV_X1 i_64_1_284 (.ZN (n_64_350), .A (n_64_1_134));
AOI222_X1 i_64_1_283 (.ZN (n_64_1_133), .A1 (n_64_87), .A2 (drc_ipo_n22), .B1 (n_64_55)
    , .B2 (n_64_1_148), .C1 (\A[20] ), .C2 (n_64_1_146));
INV_X1 i_64_1_282 (.ZN (n_64_349), .A (n_64_1_133));
AOI222_X1 i_64_1_281 (.ZN (n_64_1_132), .A1 (n_64_86), .A2 (drc_ipo_n22), .B1 (n_64_54)
    , .B2 (n_64_1_148), .C1 (\A[19] ), .C2 (n_64_1_146));
INV_X1 i_64_1_280 (.ZN (n_64_348), .A (n_64_1_132));
AOI222_X1 i_64_1_279 (.ZN (n_64_1_131), .A1 (n_64_85), .A2 (drc_ipo_n22), .B1 (n_64_53)
    , .B2 (n_64_1_148), .C1 (\A[18] ), .C2 (n_64_1_146));
INV_X1 i_64_1_278 (.ZN (n_64_347), .A (n_64_1_131));
AOI222_X1 i_64_1_277 (.ZN (n_64_1_130), .A1 (n_64_84), .A2 (drc_ipo_n22), .B1 (n_64_52)
    , .B2 (n_64_1_148), .C1 (\A[17] ), .C2 (n_64_1_146));
INV_X1 i_64_1_276 (.ZN (n_64_346), .A (n_64_1_130));
AOI222_X1 i_64_1_275 (.ZN (n_64_1_129), .A1 (n_64_83), .A2 (drc_ipo_n22), .B1 (n_64_51)
    , .B2 (n_64_1_148), .C1 (\A[16] ), .C2 (n_64_1_146));
INV_X1 i_64_1_274 (.ZN (n_64_345), .A (n_64_1_129));
AOI222_X1 i_64_1_273 (.ZN (n_64_1_128), .A1 (n_64_82), .A2 (drc_ipo_n22), .B1 (n_64_50)
    , .B2 (n_64_1_148), .C1 (\A[15] ), .C2 (n_64_1_146));
INV_X1 i_64_1_272 (.ZN (n_64_344), .A (n_64_1_128));
AOI222_X1 i_64_1_271 (.ZN (n_64_1_127), .A1 (n_64_81), .A2 (drc_ipo_n22), .B1 (n_64_49)
    , .B2 (n_64_1_148), .C1 (\A[14] ), .C2 (n_64_1_146));
INV_X1 i_64_1_270 (.ZN (n_64_343), .A (n_64_1_127));
AOI222_X1 i_64_1_269 (.ZN (n_64_1_126), .A1 (n_64_80), .A2 (drc_ipo_n22), .B1 (n_64_48)
    , .B2 (n_64_1_148), .C1 (\A[13] ), .C2 (n_64_1_146));
INV_X1 i_64_1_268 (.ZN (n_64_342), .A (n_64_1_126));
AOI222_X1 i_64_1_267 (.ZN (n_64_1_125), .A1 (n_64_79), .A2 (drc_ipo_n22), .B1 (n_64_47)
    , .B2 (n_64_1_148), .C1 (\A[12] ), .C2 (n_64_1_146));
INV_X1 i_64_1_266 (.ZN (n_64_341), .A (n_64_1_125));
AOI222_X1 i_64_1_265 (.ZN (n_64_1_124), .A1 (n_64_78), .A2 (drc_ipo_n22), .B1 (n_64_46)
    , .B2 (n_64_1_148), .C1 (\A[11] ), .C2 (n_64_1_146));
INV_X1 i_64_1_264 (.ZN (n_64_340), .A (n_64_1_124));
AOI222_X1 i_64_1_263 (.ZN (n_64_1_123), .A1 (n_64_77), .A2 (drc_ipo_n22), .B1 (n_64_45)
    , .B2 (n_64_1_148), .C1 (\A[10] ), .C2 (n_64_1_146));
INV_X1 i_64_1_262 (.ZN (n_64_339), .A (n_64_1_123));
AOI222_X1 i_64_1_261 (.ZN (n_64_1_122), .A1 (n_64_76), .A2 (drc_ipo_n22), .B1 (n_64_44)
    , .B2 (n_64_1_148), .C1 (\A[9] ), .C2 (n_64_1_146));
INV_X1 i_64_1_260 (.ZN (n_64_338), .A (n_64_1_122));
AOI222_X1 i_64_1_259 (.ZN (n_64_1_121), .A1 (n_64_75), .A2 (drc_ipo_n22), .B1 (n_64_43)
    , .B2 (n_64_1_148), .C1 (\A[8] ), .C2 (n_64_1_146));
INV_X1 i_64_1_258 (.ZN (n_64_337), .A (n_64_1_121));
AOI222_X1 i_64_1_257 (.ZN (n_64_1_120), .A1 (n_64_74), .A2 (drc_ipo_n22), .B1 (n_64_42)
    , .B2 (n_64_1_148), .C1 (\A[7] ), .C2 (n_64_1_146));
INV_X1 i_64_1_256 (.ZN (n_64_336), .A (n_64_1_120));
AOI222_X1 i_64_1_255 (.ZN (n_64_1_119), .A1 (n_64_73), .A2 (drc_ipo_n22), .B1 (n_64_41)
    , .B2 (n_64_1_148), .C1 (\A[6] ), .C2 (n_64_1_146));
INV_X1 i_64_1_254 (.ZN (n_64_335), .A (n_64_1_119));
AOI222_X1 i_64_1_253 (.ZN (n_64_1_118), .A1 (n_64_72), .A2 (drc_ipo_n22), .B1 (n_64_40)
    , .B2 (n_64_1_148), .C1 (\A[5] ), .C2 (n_64_1_146));
INV_X1 i_64_1_252 (.ZN (n_64_334), .A (n_64_1_118));
AOI222_X1 i_64_1_251 (.ZN (n_64_1_117), .A1 (n_64_71), .A2 (drc_ipo_n22), .B1 (n_64_39)
    , .B2 (n_64_1_148), .C1 (\A[4] ), .C2 (n_64_1_146));
INV_X1 i_64_1_250 (.ZN (n_64_333), .A (n_64_1_117));
AOI222_X1 i_64_1_249 (.ZN (n_64_1_116), .A1 (n_64_70), .A2 (drc_ipo_n22), .B1 (n_64_38)
    , .B2 (n_64_1_148), .C1 (\A[3] ), .C2 (n_64_1_146));
INV_X1 i_64_1_248 (.ZN (n_64_332), .A (n_64_1_116));
AOI222_X1 i_64_1_247 (.ZN (n_64_1_115), .A1 (n_64_69), .A2 (drc_ipo_n22), .B1 (n_64_37)
    , .B2 (n_64_1_148), .C1 (\A[2] ), .C2 (n_64_1_146));
INV_X1 i_64_1_246 (.ZN (n_64_331), .A (n_64_1_115));
AOI222_X1 i_64_1_245 (.ZN (n_64_1_114), .A1 (n_64_68), .A2 (drc_ipo_n22), .B1 (n_64_36)
    , .B2 (n_64_1_148), .C1 (\A[1] ), .C2 (n_64_1_146));
INV_X1 i_64_1_244 (.ZN (n_64_330), .A (n_64_1_114));
AOI222_X1 i_64_1_243 (.ZN (n_64_1_113), .A1 (n_64_67), .A2 (drc_ipo_n22), .B1 (n_64_35)
    , .B2 (n_64_1_148), .C1 (\A[0] ), .C2 (n_64_1_146));
INV_X1 i_64_1_242 (.ZN (n_64_329), .A (n_64_1_113));
INV_X1 i_64_1_240 (.ZN (n_64_1_111), .A (n_64_1_112));
AOI22_X1 i_64_1_239 (.ZN (n_64_1_110), .A1 (\Q[32] ), .A2 (n_64_1_185), .B1 (n_64_129), .B2 (n_64_1_111));
INV_X1 i_64_1_238 (.ZN (n_64_328), .A (n_64_1_110));
OAI222_X1 i_64_1_236 (.ZN (n_64_1_108), .A1 (\Q[31] ), .A2 (n_64_1_184), .B1 (n_64_128)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n54), .C2 (n_64_1_109));
INV_X1 i_64_1_235 (.ZN (n_64_327), .A (n_64_1_108));
OAI222_X1 i_64_1_234 (.ZN (n_64_1_107), .A1 (\Q[30] ), .A2 (n_64_1_184), .B1 (n_64_127)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n53), .C2 (n_64_1_109));
INV_X1 i_64_1_233 (.ZN (n_64_326), .A (n_64_1_107));
OAI222_X1 i_64_1_232 (.ZN (n_64_1_106), .A1 (\Q[29] ), .A2 (n_64_1_184), .B1 (n_64_126)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n52), .C2 (n_64_1_109));
INV_X1 i_64_1_231 (.ZN (n_64_325), .A (n_64_1_106));
OAI222_X1 i_64_1_230 (.ZN (n_64_1_105), .A1 (\Q[28] ), .A2 (n_64_1_184), .B1 (n_64_125)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n51), .C2 (n_64_1_109));
INV_X1 i_64_1_229 (.ZN (n_64_324), .A (n_64_1_105));
OAI222_X1 i_64_1_228 (.ZN (n_64_1_104), .A1 (\Q[27] ), .A2 (n_64_1_184), .B1 (n_64_124)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n50), .C2 (n_64_1_109));
INV_X1 i_64_1_227 (.ZN (n_64_323), .A (n_64_1_104));
OAI222_X1 i_64_1_226 (.ZN (n_64_1_103), .A1 (\Q[26] ), .A2 (n_64_1_184), .B1 (n_64_123)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n49), .C2 (n_64_1_109));
INV_X1 i_64_1_225 (.ZN (n_64_322), .A (n_64_1_103));
OAI222_X1 i_64_1_224 (.ZN (n_64_1_102), .A1 (\Q[25] ), .A2 (n_64_1_184), .B1 (n_64_122)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n48), .C2 (n_64_1_109));
INV_X1 i_64_1_223 (.ZN (n_64_321), .A (n_64_1_102));
OAI222_X1 i_64_1_222 (.ZN (n_64_1_101), .A1 (\Q[24] ), .A2 (n_64_1_184), .B1 (n_64_121)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n47), .C2 (n_64_1_109));
INV_X1 i_64_1_221 (.ZN (n_64_320), .A (n_64_1_101));
OAI222_X1 i_64_1_220 (.ZN (n_64_1_100), .A1 (\Q[23] ), .A2 (n_64_1_184), .B1 (n_64_120)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n46), .C2 (n_64_1_109));
INV_X1 i_64_1_219 (.ZN (n_64_319), .A (n_64_1_100));
OAI222_X1 i_64_1_218 (.ZN (n_64_1_99), .A1 (\Q[22] ), .A2 (n_64_1_184), .B1 (n_64_119)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n45), .C2 (n_64_1_109));
INV_X1 i_64_1_217 (.ZN (n_64_318), .A (n_64_1_99));
OAI222_X1 i_64_1_216 (.ZN (n_64_1_98), .A1 (\Q[21] ), .A2 (n_64_1_184), .B1 (n_64_118)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n44), .C2 (n_64_1_109));
INV_X1 i_64_1_215 (.ZN (n_64_317), .A (n_64_1_98));
OAI222_X1 i_64_1_214 (.ZN (n_64_1_97), .A1 (\Q[20] ), .A2 (n_64_1_184), .B1 (n_64_117)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n43), .C2 (n_64_1_109));
INV_X1 i_64_1_213 (.ZN (n_64_316), .A (n_64_1_97));
OAI222_X1 i_64_1_212 (.ZN (n_64_1_96), .A1 (\Q[19] ), .A2 (n_64_1_184), .B1 (n_64_116)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n42), .C2 (n_64_1_109));
INV_X1 i_64_1_211 (.ZN (n_64_315), .A (n_64_1_96));
OAI222_X1 i_64_1_210 (.ZN (n_64_1_95), .A1 (\Q[18] ), .A2 (n_64_1_184), .B1 (n_64_115)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n41), .C2 (n_64_1_109));
INV_X1 i_64_1_209 (.ZN (n_64_314), .A (n_64_1_95));
OAI222_X1 i_64_1_208 (.ZN (n_64_1_94), .A1 (\Q[17] ), .A2 (n_64_1_184), .B1 (n_64_114)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n40), .C2 (n_64_1_109));
INV_X1 i_64_1_207 (.ZN (n_64_313), .A (n_64_1_94));
OAI222_X1 i_64_1_206 (.ZN (n_64_1_93), .A1 (\Q[16] ), .A2 (n_64_1_184), .B1 (n_64_113)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n39), .C2 (n_64_1_109));
INV_X1 i_64_1_205 (.ZN (n_64_312), .A (n_64_1_93));
OAI222_X1 i_64_1_204 (.ZN (n_64_1_92), .A1 (\Q[15] ), .A2 (n_64_1_184), .B1 (n_64_112)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n38), .C2 (n_64_1_109));
INV_X1 i_64_1_203 (.ZN (n_64_311), .A (n_64_1_92));
OAI222_X1 i_64_1_202 (.ZN (n_64_1_91), .A1 (\Q[14] ), .A2 (n_64_1_184), .B1 (n_64_111)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n37), .C2 (n_64_1_109));
INV_X1 i_64_1_201 (.ZN (n_64_310), .A (n_64_1_91));
OAI222_X1 i_64_1_188 (.ZN (n_64_1_84), .A1 (\Q[7] ), .A2 (n_64_1_184), .B1 (n_64_104)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n30), .C2 (n_64_1_109));
INV_X1 i_64_1_187 (.ZN (n_64_303), .A (n_64_1_84));
OAI222_X1 i_64_1_186 (.ZN (n_64_1_83), .A1 (\Q[6] ), .A2 (n_64_1_184), .B1 (n_64_103)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n29), .C2 (n_64_1_109));
INV_X1 i_64_1_185 (.ZN (n_64_302), .A (n_64_1_83));
OAI222_X1 i_64_1_184 (.ZN (n_64_1_82), .A1 (\Q[5] ), .A2 (n_64_1_184), .B1 (n_64_102)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n28), .C2 (n_64_1_109));
INV_X1 i_64_1_183 (.ZN (n_64_301), .A (n_64_1_82));
OAI222_X1 i_64_1_182 (.ZN (n_64_1_81), .A1 (\Q[4] ), .A2 (n_64_1_184), .B1 (n_64_101)
    , .B2 (n_64_1_112), .C1 (drc_ipo_n27), .C2 (n_64_1_109));
INV_X1 i_64_1_181 (.ZN (n_64_300), .A (n_64_1_81));
OR2_X1 i_64_1_176 (.ZN (n_64_296), .A1 (drc_ipo_n89), .A2 (drc_ipo_n88));
NOR2_X1 i_64_1_175 (.ZN (n_64_295), .A1 (drc_ipo_n89), .A2 (n_64_1_144));
NOR2_X1 i_64_1_174 (.ZN (n_64_294), .A1 (drc_ipo_n89), .A2 (n_64_1_143));
NOR2_X1 i_64_1_173 (.ZN (n_64_293), .A1 (drc_ipo_n89), .A2 (n_64_1_142));
NOR2_X1 i_64_1_172 (.ZN (n_64_292), .A1 (drc_ipo_n89), .A2 (n_64_1_141));
NOR2_X1 i_64_1_171 (.ZN (n_64_291), .A1 (drc_ipo_n89), .A2 (n_64_1_140));
NOR2_X1 i_64_1_170 (.ZN (n_64_290), .A1 (drc_ipo_n89), .A2 (n_64_1_139));
NOR2_X1 i_64_1_169 (.ZN (n_64_289), .A1 (drc_ipo_n89), .A2 (n_64_1_138));
NOR2_X1 i_64_1_168 (.ZN (n_64_288), .A1 (drc_ipo_n89), .A2 (n_64_1_137));
NOR2_X1 i_64_1_167 (.ZN (n_64_287), .A1 (drc_ipo_n89), .A2 (n_64_1_136));
NOR2_X1 i_64_1_166 (.ZN (n_64_286), .A1 (drc_ipo_n89), .A2 (n_64_1_135));
NOR2_X1 i_64_1_165 (.ZN (n_64_285), .A1 (drc_ipo_n89), .A2 (n_64_1_134));
NOR2_X1 i_64_1_164 (.ZN (n_64_284), .A1 (drc_ipo_n89), .A2 (n_64_1_133));
NOR2_X1 i_64_1_163 (.ZN (n_64_283), .A1 (drc_ipo_n89), .A2 (n_64_1_132));
NOR2_X1 i_64_1_162 (.ZN (n_64_282), .A1 (drc_ipo_n89), .A2 (n_64_1_131));
NOR2_X1 i_64_1_161 (.ZN (n_64_281), .A1 (drc_ipo_n89), .A2 (n_64_1_130));
NOR2_X1 i_64_1_160 (.ZN (n_64_280), .A1 (drc_ipo_n89), .A2 (n_64_1_129));
NOR2_X1 i_64_1_159 (.ZN (n_64_279), .A1 (drc_ipo_n89), .A2 (n_64_1_128));
NOR2_X1 i_64_1_158 (.ZN (n_64_278), .A1 (drc_ipo_n89), .A2 (n_64_1_127));
NOR2_X1 i_64_1_157 (.ZN (n_64_277), .A1 (drc_ipo_n89), .A2 (n_64_1_126));
NOR2_X1 i_64_1_156 (.ZN (n_64_276), .A1 (drc_ipo_n89), .A2 (n_64_1_125));
NOR2_X1 i_64_1_155 (.ZN (n_64_275), .A1 (drc_ipo_n89), .A2 (n_64_1_124));
NOR2_X1 i_64_1_154 (.ZN (n_64_274), .A1 (drc_ipo_n89), .A2 (n_64_1_123));
NOR2_X1 i_64_1_153 (.ZN (n_64_273), .A1 (drc_ipo_n89), .A2 (n_64_1_122));
NOR2_X1 i_64_1_152 (.ZN (n_64_272), .A1 (drc_ipo_n89), .A2 (n_64_1_121));
NOR2_X1 i_64_1_151 (.ZN (n_64_271), .A1 (drc_ipo_n89), .A2 (n_64_1_120));
NOR2_X1 i_64_1_150 (.ZN (n_64_270), .A1 (drc_ipo_n89), .A2 (n_64_1_119));
NOR2_X1 i_64_1_149 (.ZN (n_64_269), .A1 (drc_ipo_n89), .A2 (n_64_1_118));
NOR2_X1 i_64_1_148 (.ZN (n_64_268), .A1 (drc_ipo_n89), .A2 (n_64_1_117));
NOR2_X1 i_64_1_147 (.ZN (n_64_267), .A1 (drc_ipo_n89), .A2 (n_64_1_116));
NOR2_X1 i_64_1_146 (.ZN (n_64_266), .A1 (drc_ipo_n89), .A2 (n_64_1_115));
NOR2_X1 i_64_1_145 (.ZN (n_64_265), .A1 (drc_ipo_n89), .A2 (n_64_1_114));
NAND2_X1 i_64_1_138 (.ZN (n_64_1_75), .A1 (n_64_189), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_137 (.ZN (n_64_260), .A (n_64_1_75), .B1 (n_64_1_142), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_136 (.ZN (n_64_1_74), .A1 (n_64_188), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_135 (.ZN (n_64_259), .A (n_64_1_74), .B1 (n_64_1_141), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_134 (.ZN (n_64_1_73), .A1 (n_64_187), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_133 (.ZN (n_64_258), .A (n_64_1_73), .B1 (n_64_1_140), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_132 (.ZN (n_64_1_72), .A1 (n_64_186), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_131 (.ZN (n_64_257), .A (n_64_1_72), .B1 (n_64_1_139), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_130 (.ZN (n_64_1_71), .A1 (n_64_185), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_129 (.ZN (n_64_256), .A (n_64_1_71), .B1 (n_64_1_138), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_128 (.ZN (n_64_1_70), .A1 (n_64_184), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_127 (.ZN (n_64_255), .A (n_64_1_70), .B1 (n_64_1_137), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_126 (.ZN (n_64_1_69), .A1 (n_64_183), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_125 (.ZN (n_64_254), .A (n_64_1_69), .B1 (n_64_1_136), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_124 (.ZN (n_64_1_68), .A1 (n_64_182), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_123 (.ZN (n_64_253), .A (n_64_1_68), .B1 (n_64_1_135), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_122 (.ZN (n_64_1_67), .A1 (n_64_181), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_121 (.ZN (n_64_252), .A (n_64_1_67), .B1 (n_64_1_134), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_120 (.ZN (n_64_1_66), .A1 (n_64_180), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_119 (.ZN (n_64_251), .A (n_64_1_66), .B1 (n_64_1_133), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_118 (.ZN (n_64_1_65), .A1 (n_64_179), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_117 (.ZN (n_64_250), .A (n_64_1_65), .B1 (n_64_1_132), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_116 (.ZN (n_64_1_64), .A1 (n_64_178), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_115 (.ZN (n_64_249), .A (n_64_1_64), .B1 (n_64_1_131), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_114 (.ZN (n_64_1_63), .A1 (n_64_177), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_113 (.ZN (n_64_248), .A (n_64_1_63), .B1 (n_64_1_130), .B2 (hfn_ipo_n17));
NAND2_X1 i_64_1_112 (.ZN (n_64_1_62), .A1 (n_64_176), .A2 (hfn_ipo_n17));
OAI21_X1 i_64_1_111 (.ZN (n_64_247), .A (n_64_1_62), .B1 (n_64_1_129), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_110 (.ZN (n_64_1_61), .A1 (n_64_175), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_109 (.ZN (n_64_246), .A (n_64_1_61), .B1 (n_64_1_128), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_108 (.ZN (n_64_1_60), .A1 (n_64_174), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_107 (.ZN (n_64_245), .A (n_64_1_60), .B1 (n_64_1_127), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_106 (.ZN (n_64_1_59), .A1 (n_64_173), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_105 (.ZN (n_64_244), .A (n_64_1_59), .B1 (n_64_1_126), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_104 (.ZN (n_64_1_58), .A1 (n_64_172), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_103 (.ZN (n_64_243), .A (n_64_1_58), .B1 (n_64_1_125), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_102 (.ZN (n_64_1_57), .A1 (n_64_171), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_101 (.ZN (n_64_242), .A (n_64_1_57), .B1 (n_64_1_124), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_100 (.ZN (n_64_1_56), .A1 (n_64_170), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_99 (.ZN (n_64_241), .A (n_64_1_56), .B1 (n_64_1_123), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_98 (.ZN (n_64_1_55), .A1 (n_64_169), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_97 (.ZN (n_64_240), .A (n_64_1_55), .B1 (n_64_1_122), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_96 (.ZN (n_64_1_54), .A1 (n_64_168), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_95 (.ZN (n_64_239), .A (n_64_1_54), .B1 (n_64_1_121), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_94 (.ZN (n_64_1_53), .A1 (n_64_167), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_93 (.ZN (n_64_238), .A (n_64_1_53), .B1 (n_64_1_120), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_92 (.ZN (n_64_1_52), .A1 (n_64_166), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_91 (.ZN (n_64_237), .A (n_64_1_52), .B1 (n_64_1_119), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_90 (.ZN (n_64_1_51), .A1 (n_64_165), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_89 (.ZN (n_64_236), .A (n_64_1_51), .B1 (n_64_1_118), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_88 (.ZN (n_64_1_50), .A1 (n_64_164), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_87 (.ZN (n_64_235), .A (n_64_1_50), .B1 (n_64_1_117), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_86 (.ZN (n_64_1_49), .A1 (n_64_163), .A2 (hfn_ipo_n18));
OAI21_X1 i_64_1_85 (.ZN (n_64_234), .A (n_64_1_49), .B1 (n_64_1_116), .B2 (hfn_ipo_n18));
NAND2_X1 i_64_1_84 (.ZN (n_64_1_48), .A1 (n_64_162), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_83 (.ZN (n_64_233), .A (n_64_1_48), .B1 (n_64_1_115), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_82 (.ZN (n_64_1_47), .A1 (n_64_161), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_81 (.ZN (n_64_232), .A (n_64_1_47), .B1 (n_64_1_114), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_80 (.ZN (n_64_1_46), .A1 (n_64_160), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_79 (.ZN (n_64_231), .A (n_64_1_46), .B1 (n_64_1_113), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_78 (.ZN (n_64_1_45), .A1 (n_64_159), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_77 (.ZN (n_64_230), .A (n_64_1_45), .B1 (n_64_1_110), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_76 (.ZN (n_64_1_44), .A1 (n_64_158), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_75 (.ZN (CLOCK_slh__n463), .A (n_64_1_44), .B1 (n_64_1_108), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_74 (.ZN (n_64_1_43), .A1 (n_64_157), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_73 (.ZN (CLOCK_slh__n491), .A (n_64_1_43), .B1 (n_64_1_107), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_72 (.ZN (n_64_1_42), .A1 (n_64_156), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_71 (.ZN (CLOCK_slh__n513), .A (n_64_1_42), .B1 (n_64_1_106), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_70 (.ZN (n_64_1_41), .A1 (n_64_155), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_69 (.ZN (CLOCK_slh__n467), .A (n_64_1_41), .B1 (n_64_1_105), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_68 (.ZN (n_64_1_40), .A1 (n_64_154), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_67 (.ZN (CLOCK_slh__n439), .A (n_64_1_40), .B1 (n_64_1_104), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_66 (.ZN (n_64_1_39), .A1 (n_64_153), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_65 (.ZN (CLOCK_slh__n479), .A (n_64_1_39), .B1 (n_64_1_103), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_64 (.ZN (n_64_1_38), .A1 (n_64_152), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_63 (.ZN (CLOCK_slh__n499), .A (n_64_1_38), .B1 (n_64_1_102), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_62 (.ZN (n_64_1_37), .A1 (n_64_151), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_61 (.ZN (CLOCK_slh__n443), .A (n_64_1_37), .B1 (n_64_1_101), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_60 (.ZN (n_64_1_36), .A1 (n_64_150), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_59 (.ZN (CLOCK_slh__n451), .A (n_64_1_36), .B1 (n_64_1_100), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_58 (.ZN (n_64_1_35), .A1 (n_64_149), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_57 (.ZN (CLOCK_slh__n471), .A (n_64_1_35), .B1 (n_64_1_99), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_56 (.ZN (n_64_1_34), .A1 (n_64_148), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_55 (.ZN (CLOCK_slh__n517), .A (n_64_1_34), .B1 (n_64_1_98), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_54 (.ZN (n_64_1_33), .A1 (n_64_147), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_53 (.ZN (CLOCK_slh__n455), .A (n_64_1_33), .B1 (n_64_1_97), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_52 (.ZN (n_64_1_32), .A1 (n_64_146), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_51 (.ZN (CLOCK_slh__n459), .A (n_64_1_32), .B1 (n_64_1_96), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_50 (.ZN (n_64_1_31), .A1 (n_64_145), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_49 (.ZN (CLOCK_slh__n495), .A (n_64_1_31), .B1 (n_64_1_95), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_48 (.ZN (n_64_1_30), .A1 (n_64_144), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_47 (.ZN (n_64_215), .A (n_64_1_30), .B1 (n_64_1_94), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_46 (.ZN (n_64_1_29), .A1 (n_64_143), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_45 (.ZN (CLOCK_slh__n431), .A (n_64_1_29), .B1 (n_64_1_93), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_44 (.ZN (n_64_1_28), .A1 (n_64_142), .A2 (hfn_ipo_n19));
OAI21_X1 i_64_1_43 (.ZN (CLOCK_slh__n427), .A (n_64_1_28), .B1 (n_64_1_92), .B2 (hfn_ipo_n19));
NAND2_X1 i_64_1_42 (.ZN (n_64_1_27), .A1 (n_64_141), .A2 (n_64_1_78));
OAI21_X1 i_64_1_41 (.ZN (CLOCK_slh__n475), .A (n_64_1_27), .B1 (n_64_1_91), .B2 (n_64_1_78));
NAND2_X1 i_64_1_40 (.ZN (n_64_1_26), .A1 (n_64_140), .A2 (n_64_1_78));
OAI21_X1 i_64_1_39 (.ZN (CLOCK_slh__n522), .A (n_64_1_26), .B1 (n_64_1_90), .B2 (n_64_1_78));
NAND2_X1 i_64_1_38 (.ZN (n_64_1_25), .A1 (n_64_139), .A2 (n_64_1_78));
OAI21_X1 i_64_1_37 (.ZN (CLOCK_slh__n511), .A (n_64_1_25), .B1 (n_64_1_89), .B2 (n_64_1_78));
NAND2_X1 i_64_1_36 (.ZN (n_64_1_24), .A1 (n_64_138), .A2 (n_64_1_78));
OAI21_X1 i_64_1_35 (.ZN (CLOCK_slh__n507), .A (n_64_1_24), .B1 (n_64_1_88), .B2 (n_64_1_78));
NAND2_X1 i_64_1_34 (.ZN (n_64_1_23), .A1 (n_64_137), .A2 (n_64_1_78));
OAI21_X1 i_64_1_33 (.ZN (CLOCK_slh__n520), .A (n_64_1_23), .B1 (n_64_1_87), .B2 (n_64_1_78));
NAND2_X1 i_64_1_32 (.ZN (n_64_1_22), .A1 (n_64_136), .A2 (n_64_1_78));
OAI21_X1 i_64_1_31 (.ZN (CLOCK_slh__n521), .A (n_64_1_22), .B1 (n_64_1_86), .B2 (n_64_1_78));
NAND2_X1 i_64_1_30 (.ZN (n_64_1_21), .A1 (n_64_135), .A2 (n_64_1_78));
OAI21_X1 i_64_1_29 (.ZN (CLOCK_slh__n515), .A (n_64_1_21), .B1 (n_64_1_85), .B2 (n_64_1_78));
NAND2_X1 i_64_1_28 (.ZN (n_64_1_20), .A1 (n_64_134), .A2 (n_64_1_78));
OAI21_X1 i_64_1_27 (.ZN (CLOCK_slh__n435), .A (n_64_1_20), .B1 (n_64_1_84), .B2 (n_64_1_78));
NAND2_X1 i_64_1_26 (.ZN (n_64_1_19), .A1 (n_64_133), .A2 (n_64_1_78));
OAI21_X1 i_64_1_25 (.ZN (CLOCK_slh__n447), .A (n_64_1_19), .B1 (n_64_1_83), .B2 (n_64_1_78));
NAND2_X1 i_64_1_24 (.ZN (n_64_1_18), .A1 (n_64_132), .A2 (n_64_1_78));
OAI21_X1 i_64_1_23 (.ZN (CLOCK_slh__n503), .A (n_64_1_18), .B1 (n_64_1_82), .B2 (n_64_1_78));
NAND2_X1 i_64_1_22 (.ZN (n_64_1_17), .A1 (n_64_131), .A2 (n_64_1_78));
OAI21_X1 i_64_1_21 (.ZN (CLOCK_slh__n483), .A (n_64_1_17), .B1 (n_64_1_81), .B2 (n_64_1_78));
NAND2_X1 i_64_1_20 (.ZN (n_64_1_16), .A1 (n_64_130), .A2 (n_64_1_78));
OAI21_X1 i_64_1_19 (.ZN (CLOCK_slh__n519), .A (n_64_1_16), .B1 (n_64_1_80), .B2 (n_64_1_78));
AOI21_X1 i_64_1_18 (.ZN (n_64_1_15), .A (out_sign), .B1 (drc_ipo_n88), .B2 (n_64_1_184));
NAND2_X1 i_64_1_17 (.ZN (n_64_1_14), .A1 (drc_ipo_n55), .A2 (n_64_1_183));
OAI21_X1 i_64_1_16 (.ZN (n_64_1_13), .A (n_64_1_14), .B1 (drc_ipo_n87), .B2 (n_64_1_109));
AOI21_X1 i_64_1_15 (.ZN (n_64_200), .A (n_64_1_15), .B1 (drc_ipo_n88), .B2 (n_64_1_13));
OAI21_X1 i_64_1_14 (.ZN (n_64_1_12), .A (n_64_296), .B1 (drc_ipo_n89), .B2 (n_64_1_190));
NAND2_X1 i_64_1_13 (.ZN (n_64_1_11), .A1 (\SC[6] ), .A2 (n_64_1_4));
OAI211_X1 i_64_1_12 (.ZN (n_64_1_10), .A (n_64_1_12), .B (n_64_1_11), .C1 (\SC[6] ), .C2 (n_64_1_4));
INV_X1 i_64_1_11 (.ZN (n_64_199), .A (n_64_1_10));
AND2_X1 i_64_1_10 (.ZN (n_64_198), .A1 (n_64_1_9), .A2 (n_64_1_12));
AND2_X1 i_64_1_9 (.ZN (n_64_197), .A1 (n_64_1_8), .A2 (n_64_1_12));
AND2_X1 i_64_1_8 (.ZN (n_64_196), .A1 (n_64_1_7), .A2 (n_64_1_12));
AND2_X1 i_64_1_7 (.ZN (n_64_195), .A1 (n_64_1_6), .A2 (n_64_1_12));
AND2_X1 i_64_1_6 (.ZN (n_64_194), .A1 (n_64_1_5), .A2 (n_64_1_12));
NOR2_X1 i_64_1_5 (.ZN (n_64_193), .A1 (drc_ipo_n89), .A2 (\SC[0] ));
HA_X1 i_64_1_4 (.CO (n_64_1_4), .S (n_64_1_9), .A (\SC[5] ), .B (n_64_1_3));
HA_X1 i_64_1_3 (.CO (n_64_1_3), .S (n_64_1_8), .A (\SC[4] ), .B (n_64_1_2));
HA_X1 i_64_1_2 (.CO (n_64_1_2), .S (n_64_1_7), .A (\SC[3] ), .B (n_64_1_1));
HA_X1 i_64_1_1 (.CO (n_64_1_1), .S (n_64_1_6), .A (\SC[2] ), .B (n_64_1_0));
HA_X1 i_64_1_0 (.CO (n_64_1_0), .S (n_64_1_5), .A (\SC[1] ), .B (\SC[0] ));
CLKGATETST_X8 clk_gate_out_sign_reg (.GCK (CTS_n_tid0_234), .CK (CTS_n_tid0_339), .E (n_64_264), .SE (1'b0 ));
CLKGATETST_X8 clk_gate_SC_reg (.GCK (CTS_n_tid1_111), .CK (CTS_n_tid0_339), .E (n_64_296), .SE (1'b0 ));
DFF_X1 out_sign_reg (.Q (out_sign), .CK (CTS_n_tid0_128), .D (n_64_200));
DFF_X1 \Q_reg[0]  (.Q (\Q[0] ), .CK (CTS_n_tid0_128), .D (n_64_297));
DFF_X1 \Q_reg[1]  (.Q (\Q[1] ), .CK (CTS_n_tid0_128), .D (n_64_298));
DFF_X1 \Q_reg[2]  (.Q (\Q[2] ), .CK (CTS_n_tid0_128), .D (n_64_299));
DFF_X1 \Q_reg[3]  (.Q (\Q[3] ), .CK (CTS_n_tid0_128), .D (n_64_300));
DFF_X1 \Q_reg[4]  (.Q (\Q[4] ), .CK (CTS_n_tid0_128), .D (n_64_301));
DFF_X1 \Q_reg[5]  (.Q (\Q[5] ), .CK (CTS_n_tid0_128), .D (n_64_302));
DFF_X1 \Q_reg[6]  (.Q (\Q[6] ), .CK (CTS_n_tid0_128), .D (n_64_303));
DFF_X1 \Q_reg[7]  (.Q (\Q[7] ), .CK (CTS_n_tid0_128), .D (n_64_304));
DFF_X1 \Q_reg[8]  (.Q (\Q[8] ), .CK (CTS_n_tid0_128), .D (n_64_305));
DFF_X1 \Q_reg[9]  (.Q (\Q[9] ), .CK (CTS_n_tid0_128), .D (n_64_306));
DFF_X1 \Q_reg[10]  (.Q (\Q[10] ), .CK (CTS_n_tid0_128), .D (n_64_307));
DFF_X1 \Q_reg[11]  (.Q (\Q[11] ), .CK (CTS_n_tid0_128), .D (n_64_308));
DFF_X1 \Q_reg[12]  (.Q (\Q[12] ), .CK (CTS_n_tid0_128), .D (n_64_309));
DFF_X1 \Q_reg[13]  (.Q (\Q[13] ), .CK (CTS_n_tid0_128), .D (n_64_310));
DFF_X1 \Q_reg[14]  (.Q (\Q[14] ), .CK (CTS_n_tid0_128), .D (n_64_311));
DFF_X1 \Q_reg[15]  (.Q (\Q[15] ), .CK (CTS_n_tid0_128), .D (n_64_312));
DFF_X1 \Q_reg[16]  (.Q (\Q[16] ), .CK (CTS_n_tid0_128), .D (n_64_313));
DFF_X1 \Q_reg[17]  (.Q (\Q[17] ), .CK (CTS_n_tid0_128), .D (n_64_314));
DFF_X1 \Q_reg[18]  (.Q (\Q[18] ), .CK (CTS_n_tid0_128), .D (n_64_315));
DFF_X1 \Q_reg[19]  (.Q (\Q[19] ), .CK (CTS_n_tid0_128), .D (n_64_316));
DFF_X1 \Q_reg[20]  (.Q (\Q[20] ), .CK (CTS_n_tid0_128), .D (n_64_317));
DFF_X1 \Q_reg[21]  (.Q (\Q[21] ), .CK (CTS_n_tid0_128), .D (n_64_318));
DFF_X1 \Q_reg[22]  (.Q (\Q[22] ), .CK (CTS_n_tid0_128), .D (n_64_319));
DFF_X1 \Q_reg[23]  (.Q (\Q[23] ), .CK (CTS_n_tid0_128), .D (n_64_320));
DFF_X1 \Q_reg[24]  (.Q (\Q[24] ), .CK (CTS_n_tid0_128), .D (n_64_321));
DFF_X1 \Q_reg[25]  (.Q (\Q[25] ), .CK (CTS_n_tid0_128), .D (n_64_322));
DFF_X1 \Q_reg[26]  (.Q (\Q[26] ), .CK (CTS_n_tid0_128), .D (n_64_323));
DFF_X1 \Q_reg[27]  (.Q (\Q[27] ), .CK (CTS_n_tid0_128), .D (n_64_324));
DFF_X1 \Q_reg[28]  (.Q (\Q[28] ), .CK (CTS_n_tid0_128), .D (n_64_325));
DFF_X1 \Q_reg[29]  (.Q (\Q[29] ), .CK (CTS_n_tid0_128), .D (n_64_326));
DFF_X1 \Q_reg[30]  (.Q (\Q[30] ), .CK (CTS_n_tid0_128), .D (n_64_327));
DFF_X1 \Q_reg[31]  (.Q (\Q[31] ), .CK (CTS_n_tid0_128), .D (n_64_328));
DFF_X1 \Q_reg[32]  (.Q (\Q[32] ), .CK (CTS_n_tid0_128), .D (n_64_329));
DFF_X1 \multiplicand_reg[0]  (.Q (\multiplicand[0] ), .CK (CTS_n_tid0_128), .D (n_64_361));
DFF_X1 \multiplicand_reg[1]  (.Q (\multiplicand[1] ), .CK (CTS_n_tid0_136), .D (n_64_362));
DFF_X1 \multiplicand_reg[2]  (.Q (\multiplicand[2] ), .CK (CTS_n_tid0_136), .D (n_64_363));
DFF_X1 \multiplicand_reg[3]  (.Q (\multiplicand[3] ), .CK (CTS_n_tid0_136), .D (n_64_364));
DFF_X1 \multiplicand_reg[4]  (.Q (\multiplicand[4] ), .CK (CTS_n_tid0_136), .D (n_64_365));
DFF_X1 \multiplicand_reg[5]  (.Q (\multiplicand[5] ), .CK (CTS_n_tid0_136), .D (n_64_366));
DFF_X1 \multiplicand_reg[6]  (.Q (\multiplicand[6] ), .CK (CTS_n_tid0_136), .D (n_64_367));
DFF_X1 \multiplicand_reg[7]  (.Q (\multiplicand[7] ), .CK (CTS_n_tid0_136), .D (n_64_368));
DFF_X1 \multiplicand_reg[8]  (.Q (\multiplicand[8] ), .CK (CTS_n_tid0_136), .D (n_64_369));
DFF_X1 \multiplicand_reg[9]  (.Q (\multiplicand[9] ), .CK (CTS_n_tid0_136), .D (n_64_370));
DFF_X1 \multiplicand_reg[10]  (.Q (\multiplicand[10] ), .CK (CTS_n_tid0_136), .D (n_64_371));
DFF_X1 \multiplicand_reg[11]  (.Q (\multiplicand[11] ), .CK (CTS_n_tid0_136), .D (n_64_372));
DFF_X1 \multiplicand_reg[12]  (.Q (\multiplicand[12] ), .CK (CTS_n_tid0_136), .D (n_64_373));
DFF_X1 \multiplicand_reg[13]  (.Q (\multiplicand[13] ), .CK (CTS_n_tid0_136), .D (n_64_374));
DFF_X1 \multiplicand_reg[14]  (.Q (\multiplicand[14] ), .CK (CTS_n_tid0_136), .D (n_64_375));
DFF_X1 \multiplicand_reg[15]  (.Q (\multiplicand[15] ), .CK (CTS_n_tid0_136), .D (n_64_376));
DFF_X1 \multiplicand_reg[16]  (.Q (\multiplicand[16] ), .CK (CTS_n_tid0_136), .D (n_64_377));
DFF_X1 \multiplicand_reg[17]  (.Q (\multiplicand[17] ), .CK (CTS_n_tid0_136), .D (n_64_378));
DFF_X1 \multiplicand_reg[18]  (.Q (\multiplicand[18] ), .CK (CTS_n_tid0_136), .D (n_64_379));
DFF_X1 \multiplicand_reg[19]  (.Q (\multiplicand[19] ), .CK (CTS_n_tid0_136), .D (n_64_380));
DFF_X1 \multiplicand_reg[20]  (.Q (\multiplicand[20] ), .CK (CTS_n_tid0_136), .D (n_64_381));
DFF_X1 \multiplicand_reg[21]  (.Q (\multiplicand[21] ), .CK (CTS_n_tid0_136), .D (n_64_382));
DFF_X1 \multiplicand_reg[22]  (.Q (\multiplicand[22] ), .CK (CTS_n_tid0_136), .D (n_64_383));
DFF_X1 \multiplicand_reg[23]  (.Q (\multiplicand[23] ), .CK (CTS_n_tid0_136), .D (n_64_384));
DFF_X1 \multiplicand_reg[24]  (.Q (\multiplicand[24] ), .CK (CTS_n_tid0_136), .D (n_64_385));
DFF_X1 \multiplicand_reg[25]  (.Q (\multiplicand[25] ), .CK (CTS_n_tid0_136), .D (n_64_386));
DFF_X1 \multiplicand_reg[26]  (.Q (\multiplicand[26] ), .CK (CTS_n_tid0_136), .D (n_64_387));
DFF_X1 \multiplicand_reg[27]  (.Q (\multiplicand[27] ), .CK (CTS_n_tid0_128), .D (n_64_388));
DFF_X1 \multiplicand_reg[28]  (.Q (\multiplicand[28] ), .CK (CTS_n_tid0_136), .D (n_64_389));
DFF_X1 \multiplicand_reg[29]  (.Q (\multiplicand[29] ), .CK (CTS_n_tid0_128), .D (n_64_390));
DFF_X1 \multiplicand_reg[30]  (.Q (\multiplicand[30] ), .CK (CTS_n_tid0_128), .D (n_64_391));
DFF_X1 \multiplicand_reg[31]  (.Q (\multiplicand[31] ), .CK (CTS_n_tid0_128), .D (n_64_392));
DFF_X1 \SC_reg[0]  (.Q (\SC[0] ), .CK (CTS_n_tid1_109), .D (n_64_193));
DFF_X1 \SC_reg[1]  (.Q (\SC[1] ), .CK (CTS_n_tid1_109), .D (n_64_194));
DFF_X1 \SC_reg[2]  (.Q (\SC[2] ), .CK (CTS_n_tid1_109), .D (n_64_195));
DFF_X1 \SC_reg[3]  (.Q (\SC[3] ), .CK (CTS_n_tid1_109), .D (n_64_196));
DFF_X1 \SC_reg[4]  (.Q (\SC[4] ), .CK (CTS_n_tid1_109), .D (n_64_197));
DFF_X1 \SC_reg[5]  (.Q (\SC[5] ), .CK (CTS_n_tid1_109), .D (n_64_198));
DFF_X1 \SC_reg[6]  (.Q (\SC[6] ), .CK (CTS_n_tid1_109), .D (n_64_199));
DFF_X1 \A_reg[0]  (.Q (\A[0] ), .CK (CTS_n_tid1_109), .D (n_64_265));
DFF_X1 \A_reg[1]  (.Q (\A[1] ), .CK (CTS_n_tid1_109), .D (n_64_266));
DFF_X1 \A_reg[2]  (.Q (\A[2] ), .CK (CTS_n_tid1_109), .D (n_64_267));
DFF_X1 \A_reg[3]  (.Q (\A[3] ), .CK (CTS_n_tid1_109), .D (n_64_268));
DFF_X1 \A_reg[4]  (.Q (\A[4] ), .CK (CTS_n_tid1_109), .D (n_64_269));
DFF_X1 \A_reg[5]  (.Q (\A[5] ), .CK (CTS_n_tid1_109), .D (n_64_270));
DFF_X1 \A_reg[6]  (.Q (\A[6] ), .CK (CTS_n_tid1_109), .D (n_64_271));
DFF_X1 \A_reg[7]  (.Q (\A[7] ), .CK (CTS_n_tid1_109), .D (n_64_272));
DFF_X1 \A_reg[8]  (.Q (\A[8] ), .CK (CTS_n_tid1_109), .D (n_64_273));
DFF_X1 \A_reg[9]  (.Q (\A[9] ), .CK (CTS_n_tid1_109), .D (n_64_274));
DFF_X1 \A_reg[10]  (.Q (\A[10] ), .CK (CTS_n_tid1_109), .D (n_64_275));
DFF_X1 \A_reg[11]  (.Q (\A[11] ), .CK (CTS_n_tid1_109), .D (n_64_276));
DFF_X1 \A_reg[12]  (.Q (\A[12] ), .CK (CTS_n_tid1_109), .D (n_64_277));
DFF_X1 \A_reg[13]  (.Q (\A[13] ), .CK (CTS_n_tid1_109), .D (n_64_278));
DFF_X1 \A_reg[14]  (.Q (\A[14] ), .CK (CTS_n_tid1_109), .D (n_64_279));
DFF_X1 \A_reg[15]  (.Q (\A[15] ), .CK (CTS_n_tid1_109), .D (n_64_280));
DFF_X1 \A_reg[16]  (.Q (\A[16] ), .CK (CTS_n_tid1_109), .D (n_64_281));
DFF_X1 \A_reg[17]  (.Q (\A[17] ), .CK (CTS_n_tid1_109), .D (n_64_282));
DFF_X1 \A_reg[18]  (.Q (\A[18] ), .CK (CTS_n_tid1_109), .D (n_64_283));
DFF_X1 \A_reg[19]  (.Q (\A[19] ), .CK (CTS_n_tid1_109), .D (n_64_284));
DFF_X1 \A_reg[20]  (.Q (\A[20] ), .CK (CTS_n_tid1_109), .D (n_64_285));
DFF_X1 \A_reg[21]  (.Q (\A[21] ), .CK (CTS_n_tid1_109), .D (n_64_286));
DFF_X1 \A_reg[22]  (.Q (\A[22] ), .CK (CTS_n_tid1_109), .D (n_64_287));
DFF_X1 \A_reg[23]  (.Q (\A[23] ), .CK (CTS_n_tid1_109), .D (n_64_288));
DFF_X1 \A_reg[24]  (.Q (\A[24] ), .CK (CTS_n_tid1_109), .D (n_64_289));
DFF_X1 \A_reg[25]  (.Q (\A[25] ), .CK (CTS_n_tid1_109), .D (n_64_290));
DFF_X1 \A_reg[26]  (.Q (\A[26] ), .CK (CTS_n_tid1_109), .D (n_64_291));
DFF_X1 \A_reg[27]  (.Q (\A[27] ), .CK (CTS_n_tid1_109), .D (n_64_292));
DFF_X1 \A_reg[28]  (.Q (\A[28] ), .CK (CTS_n_tid1_109), .D (n_64_293));
DFF_X1 \A_reg[29]  (.Q (\A[29] ), .CK (CTS_n_tid1_109), .D (n_64_294));
DFF_X1 \A_reg[31]  (.Q (\A[31] ), .CK (CTS_n_tid1_109), .D (n_64_295));
datapath__0_72 i_64_203 (.p_0 ({n_64_192, n_64_191, n_64_190, n_64_189, n_64_188, 
    n_64_187, n_64_186, n_64_185, n_64_184, n_64_183, n_64_182, n_64_181, n_64_180, 
    n_64_179, n_64_178, n_64_177, n_64_176, n_64_175, n_64_174, n_64_173, n_64_172, 
    n_64_171, n_64_170, n_64_169, n_64_168, n_64_167, n_64_166, n_64_165, n_64_164, 
    n_64_163, n_64_162, n_64_161, n_64_160, n_64_159, n_64_158, n_64_157, n_64_156, 
    n_64_155, n_64_154, n_64_153, n_64_152, n_64_151, n_64_150, n_64_149, n_64_148, 
    n_64_147, n_64_146, n_64_145, n_64_144, n_64_143, n_64_142, n_64_141, n_64_140, 
    n_64_139, n_64_138, n_64_137, n_64_136, n_64_135, n_64_134, n_64_133, n_64_132, 
    n_64_131, n_64_130, uc_4}), .p_1 ({uc_5, n_64_1_79, n_64_359, n_64_358, n_64_357, 
    n_64_356, n_64_355, n_64_354, n_64_353, n_64_352, n_64_351, n_64_350, n_64_349, 
    n_64_348, n_64_347, n_64_346, n_64_345, n_64_344, n_64_343, n_64_342, n_64_341, 
    n_64_340, n_64_339, n_64_338, n_64_337, n_64_336, n_64_335, n_64_334, n_64_333, 
    n_64_332, n_64_331, n_64_330, n_64_329, n_64_328, n_64_327, n_64_326, n_64_325, 
    n_64_324, n_64_323, n_64_322, n_64_321, n_64_320, n_64_319, n_64_318, n_64_317, 
    n_64_316, n_64_315, n_64_314, n_64_313, n_64_312, n_64_311, n_64_310, n_64_309, 
    n_64_308, n_64_307, n_64_306, n_64_305, n_64_304, n_64_303, n_64_302, n_64_301, 
    n_64_300, n_64_299, n_64_298}));
datapath__0_67 i_64_198 (.p_0 ({n_64_129, n_64_128, n_64_127, n_64_126, n_64_125, 
    n_64_124, n_64_123, n_64_122, n_64_121, n_64_120, n_64_119, n_64_118, n_64_117, 
    n_64_116, n_64_115, n_64_114, n_64_113, n_64_112, n_64_111, n_64_110, n_64_109, 
    n_64_108, n_64_107, n_64_106, n_64_105, n_64_104, n_64_103, n_64_102, n_64_101, 
    n_64_100, n_64_99, uc_3}), .b ({drc_ipo_n55, drc_ipo_n54, drc_ipo_n53, drc_ipo_n52, 
    drc_ipo_n51, drc_ipo_n50, drc_ipo_n49, drc_ipo_n48, drc_ipo_n47, drc_ipo_n46, 
    drc_ipo_n45, drc_ipo_n44, drc_ipo_n43, drc_ipo_n42, drc_ipo_n41, drc_ipo_n40, 
    drc_ipo_n39, drc_ipo_n38, drc_ipo_n37, drc_ipo_n36, drc_ipo_n35, drc_ipo_n34, 
    drc_ipo_n33, drc_ipo_n32, drc_ipo_n31, drc_ipo_n30, drc_ipo_n29, drc_ipo_n28, 
    drc_ipo_n27, drc_ipo_n26, drc_ipo_n25, drc_ipo_n24}));
datapath__0_66 i_64_197 (.p_0 ({n_64_98, n_64_97, n_64_96, n_64_95, n_64_94, n_64_93, 
    n_64_92, n_64_91, n_64_90, n_64_89, n_64_88, n_64_87, n_64_86, n_64_85, n_64_84, 
    n_64_83, n_64_82, n_64_81, n_64_80, n_64_79, n_64_78, n_64_77, n_64_76, n_64_75, 
    n_64_74, n_64_73, n_64_72, n_64_71, n_64_70, n_64_69, n_64_68, n_64_67}), .A ({
    \A[31] , uc_2, \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] , 
    \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] , \A[15] , \A[14] , 
    \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , 
    \A[3] , \A[2] , \A[1] , \A[0] }), .multiplicand ({n_64_392, n_64_391, n_64_390, 
    n_64_389, n_64_388, n_64_387, n_64_386, n_64_385, n_64_384, n_64_383, n_64_382, 
    n_64_381, n_64_380, n_64_379, n_64_378, n_64_377, n_64_376, n_64_375, n_64_374, 
    n_64_373, n_64_372, n_64_371, n_64_370, n_64_369, n_64_368, n_64_367, n_64_366, 
    n_64_365, n_64_364, n_64_363, n_64_362, n_64_361}));
datapath__0_65 i_64_196 (.p_0 ({n_64_66, n_64_65, n_64_64, n_64_63, n_64_62, n_64_61, 
    n_64_60, n_64_59, n_64_58, n_64_57, n_64_56, n_64_55, n_64_54, n_64_53, n_64_52, 
    n_64_51, n_64_50, n_64_49, n_64_48, n_64_47, n_64_46, n_64_45, n_64_44, n_64_43, 
    n_64_42, n_64_41, n_64_40, n_64_39, n_64_38, n_64_37, n_64_36, n_64_35}), .A ({
    \A[31] , uc_1, \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] , 
    \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] , \A[15] , \A[14] , 
    \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , 
    \A[3] , \A[2] , \A[1] , \A[0] }), .multiplicand ({n_64_392, n_64_391, n_64_390, 
    n_64_389, n_64_388, n_64_387, n_64_386, n_64_385, n_64_384, n_64_383, n_64_382, 
    n_64_381, n_64_380, n_64_379, n_64_378, n_64_377, n_64_376, n_64_375, n_64_374, 
    n_64_373, n_64_372, n_64_371, n_64_370, n_64_369, n_64_368, n_64_367, n_64_366, 
    n_64_365, n_64_364, n_64_363, n_64_362, n_64_361}));
datapath i_64_194 (.p_0 ({n_64_34, n_64_33, n_64_32, n_64_31, n_64_30, n_64_29, n_64_28, 
    n_64_27, n_64_26, n_64_25, n_64_24, n_64_23, n_64_22, n_64_21, n_64_20, n_64_19, 
    n_64_18, n_64_17, n_64_16, n_64_15, n_64_14, n_64_13, n_64_12, n_64_11, n_64_10, 
    n_64_9, n_64_8, n_64_7, n_64_6, n_64_5, n_64_4, uc_0}), .a ({drc_ipo_n87, drc_ipo_n86, 
    drc_ipo_n85, drc_ipo_n84, drc_ipo_n83, drc_ipo_n82, drc_ipo_n81, drc_ipo_n80, 
    drc_ipo_n79, drc_ipo_n78, drc_ipo_n77, drc_ipo_n76, drc_ipo_n75, drc_ipo_n74, 
    drc_ipo_n73, drc_ipo_n72, drc_ipo_n71, drc_ipo_n70, drc_ipo_n69, drc_ipo_n68, 
    drc_ipo_n67, drc_ipo_n66, drc_ipo_n65, drc_ipo_n64, drc_ipo_n63, drc_ipo_n62, 
    drc_ipo_n61, drc_ipo_n60, drc_ipo_n59, drc_ipo_n58, drc_ipo_n57, drc_ipo_n56}));
DFF_X1 i_64_64 (.Q (n_64_3), .CK (CTS_n_tid0_336), .D (n_64_394));
DFF_X1 \c_reg[0]  (.Q (n_64), .CK (CTS_n_tid1_243), .D (n_64_298));
DFF_X1 \c_reg[1]  (.Q (n_63), .CK (CTS_n_tid1_243), .D (n_64_201));
DFF_X1 \c_reg[2]  (.Q (n_62), .CK (CTS_n_tid1_243), .D (n_64_202));
DFF_X1 \c_reg[3]  (.Q (n_61), .CK (CTS_n_tid1_243), .D (n_64_203));
DFF_X1 \c_reg[4]  (.Q (n_60), .CK (CTS_n_tid1_243), .D (n_64_204));
DFF_X1 \c_reg[5]  (.Q (n_59), .CK (CTS_n_tid1_243), .D (n_64_205));
DFF_X1 \c_reg[6]  (.Q (n_58), .CK (CTS_n_tid1_243), .D (n_64_206));
DFF_X1 \c_reg[7]  (.Q (n_57), .CK (CTS_n_tid1_243), .D (n_64_207));
DFF_X1 \c_reg[8]  (.Q (n_56), .CK (CTS_n_tid1_243), .D (n_64_208));
DFF_X1 \c_reg[9]  (.Q (n_55), .CK (CTS_n_tid1_243), .D (n_64_209));
DFF_X1 \c_reg[10]  (.Q (n_54), .CK (CTS_n_tid1_243), .D (n_64_210));
DFF_X1 \c_reg[11]  (.Q (n_53), .CK (CTS_n_tid1_243), .D (n_64_211));
DFF_X1 \c_reg[12]  (.Q (n_52), .CK (CTS_n_tid1_243), .D (n_64_212));
DFF_X1 \c_reg[13]  (.Q (n_51), .CK (CTS_n_tid1_243), .D (n_64_213));
DFF_X1 \c_reg[14]  (.Q (n_50), .CK (CTS_n_tid1_243), .D (n_64_214));
DFF_X1 \c_reg[15]  (.Q (n_49), .CK (CTS_n_tid1_243), .D (n_64_215));
DFF_X1 \c_reg[16]  (.Q (n_48), .CK (CTS_n_tid1_243), .D (n_64_216));
DFF_X1 \c_reg[17]  (.Q (n_47), .CK (CTS_n_tid1_243), .D (n_64_217));
DFF_X1 \c_reg[18]  (.Q (n_46), .CK (CTS_n_tid1_243), .D (n_64_218));
DFF_X1 \c_reg[19]  (.Q (n_45), .CK (CTS_n_tid1_243), .D (n_64_219));
DFF_X1 \c_reg[20]  (.Q (n_44), .CK (CTS_n_tid1_243), .D (n_64_220));
DFF_X1 \c_reg[21]  (.Q (n_43), .CK (CTS_n_tid1_243), .D (n_64_221));
DFF_X1 \c_reg[22]  (.Q (n_42), .CK (CTS_n_tid1_243), .D (n_64_222));
DFF_X1 \c_reg[23]  (.Q (n_41), .CK (CTS_n_tid1_243), .D (n_64_223));
DFF_X1 \c_reg[24]  (.Q (n_40), .CK (CTS_n_tid1_243), .D (n_64_224));
DFF_X1 \c_reg[25]  (.Q (n_39), .CK (CTS_n_tid1_243), .D (n_64_225));
DFF_X1 \c_reg[26]  (.Q (n_38), .CK (CTS_n_tid1_243), .D (n_64_226));
DFF_X1 \c_reg[27]  (.Q (n_37), .CK (CTS_n_tid1_243), .D (n_64_227));
DFF_X1 \c_reg[28]  (.Q (n_36), .CK (CTS_n_tid1_243), .D (n_64_228));
DFF_X1 \c_reg[29]  (.Q (n_35), .CK (CTS_n_tid1_243), .D (n_64_229));
DFF_X1 \c_reg[30]  (.Q (n_34), .CK (CTS_n_tid1_243), .D (n_64_230));
DFF_X1 \c_reg[31]  (.Q (n_33), .CK (CTS_n_tid1_243), .D (n_64_231));
DFF_X1 \c_reg[32]  (.Q (n_32), .CK (CTS_n_tid1_243), .D (n_64_232));
DFF_X1 \c_reg[33]  (.Q (n_31), .CK (CTS_n_tid1_243), .D (n_64_233));
DFF_X1 \c_reg[34]  (.Q (n_30), .CK (CTS_n_tid1_243), .D (n_64_234));
DFF_X1 \c_reg[35]  (.Q (n_29), .CK (CTS_n_tid1_243), .D (n_64_235));
DFF_X1 \c_reg[36]  (.Q (n_28), .CK (CTS_n_tid1_243), .D (n_64_236));
DFF_X1 \c_reg[37]  (.Q (n_27), .CK (CTS_n_tid1_243), .D (n_64_237));
DFF_X1 \c_reg[38]  (.Q (n_26), .CK (CTS_n_tid1_243), .D (n_64_238));
DFF_X1 \c_reg[39]  (.Q (n_25), .CK (CTS_n_tid1_243), .D (n_64_239));
DFF_X1 \c_reg[40]  (.Q (n_24), .CK (CTS_n_tid1_243), .D (n_64_240));
DFF_X1 \c_reg[41]  (.Q (n_23), .CK (CTS_n_tid1_243), .D (n_64_241));
DFF_X1 \c_reg[42]  (.Q (n_22), .CK (CTS_n_tid1_243), .D (n_64_242));
DFF_X1 \c_reg[43]  (.Q (n_21), .CK (CTS_n_tid1_243), .D (n_64_243));
DFF_X1 \c_reg[44]  (.Q (n_20), .CK (CTS_n_tid1_243), .D (n_64_244));
DFF_X1 \c_reg[45]  (.Q (n_19), .CK (CTS_n_tid1_243), .D (n_64_245));
DFF_X1 \c_reg[46]  (.Q (n_18), .CK (CTS_n_tid1_243), .D (n_64_246));
DFF_X1 \c_reg[47]  (.Q (n_17), .CK (CTS_n_tid1_243), .D (n_64_247));
DFF_X1 \c_reg[48]  (.Q (n_16), .CK (CTS_n_tid1_243), .D (n_64_248));
DFF_X1 \c_reg[49]  (.Q (n_15), .CK (CTS_n_tid1_243), .D (n_64_249));
DFF_X1 \c_reg[50]  (.Q (n_14), .CK (CTS_n_tid1_243), .D (n_64_250));
DFF_X1 \c_reg[51]  (.Q (n_13), .CK (CTS_n_tid1_243), .D (n_64_251));
DFF_X1 \c_reg[52]  (.Q (n_12), .CK (CTS_n_tid1_243), .D (n_64_252));
DFF_X1 \c_reg[53]  (.Q (n_11), .CK (CTS_n_tid1_243), .D (n_64_253));
DFF_X1 \c_reg[54]  (.Q (n_10), .CK (CTS_n_tid1_243), .D (n_64_254));
DFF_X1 \c_reg[55]  (.Q (n_9), .CK (CTS_n_tid1_243), .D (n_64_255));
DFF_X1 \c_reg[56]  (.Q (n_8), .CK (CTS_n_tid1_243), .D (n_64_256));
DFF_X1 \c_reg[57]  (.Q (n_7), .CK (CTS_n_tid1_243), .D (n_64_257));
DFF_X1 \c_reg[58]  (.Q (n_6), .CK (CTS_n_tid1_243), .D (n_64_258));
DFF_X1 \c_reg[59]  (.Q (n_5), .CK (CTS_n_tid1_243), .D (n_64_259));
DFF_X1 \c_reg[60]  (.Q (n_4), .CK (CTS_n_tid1_243), .D (n_64_260));
DFF_X1 \c_reg[61]  (.Q (n_3), .CK (CTS_n_tid1_243), .D (n_64_261));
DFF_X1 \c_reg[62]  (.Q (n_2), .CK (CTS_n_tid1_243), .D (n_64_262));
DFF_X1 \c_reg[63]  (.Q (n_1), .CK (CTS_n_tid1_243), .D (n_64_263));
CLKGATETST_X8 clk_gate_c_reg (.GCK (CTS_n_tid1_244), .CK (CTS_n_tid0_339), .E (n_64_393), .SE (1'b0 ));
INV_X1 i_64_0 (.ZN (n_0), .A (n_64_3));
TBUF_X1 i_63 (.Z (c[63]), .A (n_1), .EN (hfn_ipo_n20));
TBUF_X1 i_62 (.Z (c[62]), .A (n_2), .EN (hfn_ipo_n21));
TBUF_X1 i_61 (.Z (c[61]), .A (n_3), .EN (hfn_ipo_n20));
TBUF_X1 i_60 (.Z (c[60]), .A (n_4), .EN (hfn_ipo_n20));
TBUF_X1 i_59 (.Z (c[59]), .A (n_5), .EN (hfn_ipo_n20));
TBUF_X1 i_58 (.Z (c[58]), .A (n_6), .EN (hfn_ipo_n20));
TBUF_X1 i_57 (.Z (c[57]), .A (n_7), .EN (hfn_ipo_n20));
TBUF_X1 i_56 (.Z (c[56]), .A (n_8), .EN (hfn_ipo_n20));
TBUF_X1 i_55 (.Z (c[55]), .A (n_9), .EN (hfn_ipo_n20));
TBUF_X1 i_54 (.Z (c[54]), .A (n_10), .EN (hfn_ipo_n20));
TBUF_X1 i_53 (.Z (c[53]), .A (n_11), .EN (hfn_ipo_n20));
TBUF_X1 i_52 (.Z (c[52]), .A (n_12), .EN (hfn_ipo_n20));
TBUF_X1 i_51 (.Z (c[51]), .A (n_13), .EN (hfn_ipo_n20));
TBUF_X1 i_50 (.Z (c[50]), .A (n_14), .EN (hfn_ipo_n20));
TBUF_X1 i_49 (.Z (c[49]), .A (n_15), .EN (hfn_ipo_n20));
TBUF_X1 i_48 (.Z (c[48]), .A (n_16), .EN (hfn_ipo_n20));
TBUF_X1 i_47 (.Z (c[47]), .A (n_17), .EN (hfn_ipo_n20));
TBUF_X1 i_46 (.Z (c[46]), .A (n_18), .EN (hfn_ipo_n20));
TBUF_X1 i_45 (.Z (c[45]), .A (n_19), .EN (hfn_ipo_n20));
TBUF_X1 i_44 (.Z (c[44]), .A (n_20), .EN (hfn_ipo_n20));
TBUF_X1 i_43 (.Z (c[43]), .A (n_21), .EN (hfn_ipo_n20));
TBUF_X1 i_42 (.Z (c[42]), .A (n_22), .EN (hfn_ipo_n20));
TBUF_X1 i_41 (.Z (c[41]), .A (n_23), .EN (hfn_ipo_n20));
TBUF_X1 i_40 (.Z (c[40]), .A (n_24), .EN (hfn_ipo_n20));
TBUF_X1 i_39 (.Z (c[39]), .A (n_25), .EN (hfn_ipo_n20));
TBUF_X1 i_38 (.Z (c[38]), .A (n_26), .EN (hfn_ipo_n20));
TBUF_X1 i_37 (.Z (c[37]), .A (n_27), .EN (hfn_ipo_n21));
TBUF_X1 i_36 (.Z (c[36]), .A (n_28), .EN (hfn_ipo_n21));
TBUF_X1 i_35 (.Z (c[35]), .A (n_29), .EN (hfn_ipo_n21));
TBUF_X1 i_34 (.Z (c[34]), .A (n_30), .EN (hfn_ipo_n21));
TBUF_X1 i_33 (.Z (c[33]), .A (n_31), .EN (hfn_ipo_n21));
TBUF_X1 i_32 (.Z (c[32]), .A (n_32), .EN (hfn_ipo_n21));
TBUF_X1 i_31 (.Z (c[31]), .A (n_33), .EN (hfn_ipo_n21));
TBUF_X1 i_30 (.Z (c[30]), .A (n_34), .EN (hfn_ipo_n21));
TBUF_X1 i_29 (.Z (c[29]), .A (n_35), .EN (hfn_ipo_n21));
TBUF_X1 i_28 (.Z (c[28]), .A (n_36), .EN (hfn_ipo_n21));
TBUF_X1 i_27 (.Z (c[27]), .A (n_37), .EN (hfn_ipo_n21));
TBUF_X1 i_26 (.Z (c[26]), .A (n_38), .EN (hfn_ipo_n21));
TBUF_X1 i_25 (.Z (c[25]), .A (n_39), .EN (hfn_ipo_n21));
TBUF_X1 i_24 (.Z (c[24]), .A (n_40), .EN (hfn_ipo_n21));
TBUF_X1 i_23 (.Z (c[23]), .A (n_41), .EN (hfn_ipo_n21));
TBUF_X1 i_22 (.Z (c[22]), .A (n_42), .EN (hfn_ipo_n21));
TBUF_X1 i_21 (.Z (c[21]), .A (n_43), .EN (hfn_ipo_n21));
TBUF_X1 i_20 (.Z (c[20]), .A (n_44), .EN (hfn_ipo_n21));
TBUF_X1 i_19 (.Z (c[19]), .A (n_45), .EN (hfn_ipo_n21));
TBUF_X1 i_18 (.Z (c[18]), .A (n_46), .EN (hfn_ipo_n21));
TBUF_X1 i_17 (.Z (c[17]), .A (n_47), .EN (hfn_ipo_n21));
TBUF_X1 i_16 (.Z (c[16]), .A (n_48), .EN (hfn_ipo_n21));
TBUF_X1 i_15 (.Z (c[15]), .A (n_49), .EN (hfn_ipo_n21));
TBUF_X1 i_14 (.Z (c[14]), .A (n_50), .EN (hfn_ipo_n21));
TBUF_X1 i_13 (.Z (c[13]), .A (n_51), .EN (hfn_ipo_n21));
TBUF_X1 i_12 (.Z (c[12]), .A (n_52), .EN (hfn_ipo_n21));
TBUF_X1 i_11 (.Z (c[11]), .A (n_53), .EN (hfn_ipo_n20));
TBUF_X1 i_10 (.Z (c[10]), .A (n_54), .EN (hfn_ipo_n20));
TBUF_X1 i_9 (.Z (c[9]), .A (n_55), .EN (hfn_ipo_n20));
TBUF_X1 i_8 (.Z (c[8]), .A (n_56), .EN (hfn_ipo_n20));
TBUF_X1 i_7 (.Z (c[7]), .A (n_57), .EN (hfn_ipo_n20));
TBUF_X1 i_6 (.Z (c[6]), .A (n_58), .EN (hfn_ipo_n20));
TBUF_X1 i_5 (.Z (c[5]), .A (n_59), .EN (hfn_ipo_n20));
TBUF_X1 i_4 (.Z (c[4]), .A (n_60), .EN (hfn_ipo_n20));
TBUF_X1 i_3 (.Z (c[3]), .A (n_61), .EN (hfn_ipo_n20));
TBUF_X1 i_2 (.Z (c[2]), .A (n_62), .EN (hfn_ipo_n20));
TBUF_X1 i_1 (.Z (c[1]), .A (n_63), .EN (hfn_ipo_n20));
TBUF_X1 i_0 (.Z (c[0]), .A (n_64), .EN (hfn_ipo_n20));
BUF_X4 hfn_ipo_c20 (.Z (hfn_ipo_n20), .A (n_0));
CLKBUF_X2 hfn_ipo_c21 (.Z (hfn_ipo_n21), .A (n_0));
BUF_X4 drc_ipo_c22 (.Z (drc_ipo_n22), .A (n_64_1_147));
CLKBUF_X3 CTS_L3_c_tid1_111 (.Z (CTS_n_tid1_109), .A (CTS_n_tid1_111));
CLKBUF_X1 CTS_L4_c_tid0_287 (.Z (CTS_n_tid0_336), .A (CTS_n_tid0_337));
CLKBUF_X2 hfn_ipo_c17 (.Z (hfn_ipo_n17), .A (n_64_1_78));
CLKBUF_X1 hfn_ipo_c18 (.Z (hfn_ipo_n18), .A (n_64_1_78));
CLKBUF_X1 drc_ipo_c24 (.Z (drc_ipo_n24), .A (b[0]));
CLKBUF_X1 drc_ipo_c25 (.Z (drc_ipo_n25), .A (b[1]));
CLKBUF_X1 drc_ipo_c26 (.Z (drc_ipo_n26), .A (b[2]));
CLKBUF_X1 drc_ipo_c27 (.Z (drc_ipo_n27), .A (b[3]));
CLKBUF_X1 drc_ipo_c28 (.Z (drc_ipo_n28), .A (b[4]));
CLKBUF_X1 drc_ipo_c29 (.Z (drc_ipo_n29), .A (b[5]));
CLKBUF_X1 drc_ipo_c30 (.Z (drc_ipo_n30), .A (b[6]));
CLKBUF_X1 drc_ipo_c31 (.Z (drc_ipo_n31), .A (b[7]));
CLKBUF_X1 drc_ipo_c32 (.Z (drc_ipo_n32), .A (b[8]));
CLKBUF_X1 drc_ipo_c33 (.Z (drc_ipo_n33), .A (b[9]));
CLKBUF_X1 drc_ipo_c34 (.Z (drc_ipo_n34), .A (b[10]));
CLKBUF_X1 drc_ipo_c35 (.Z (drc_ipo_n35), .A (b[11]));
CLKBUF_X1 drc_ipo_c36 (.Z (drc_ipo_n36), .A (b[12]));
CLKBUF_X1 drc_ipo_c37 (.Z (drc_ipo_n37), .A (b[13]));
CLKBUF_X1 drc_ipo_c38 (.Z (drc_ipo_n38), .A (b[14]));
CLKBUF_X1 drc_ipo_c39 (.Z (drc_ipo_n39), .A (b[15]));
CLKBUF_X1 drc_ipo_c40 (.Z (drc_ipo_n40), .A (b[16]));
CLKBUF_X1 drc_ipo_c41 (.Z (drc_ipo_n41), .A (b[17]));
CLKBUF_X1 drc_ipo_c42 (.Z (drc_ipo_n42), .A (b[18]));
CLKBUF_X1 drc_ipo_c43 (.Z (drc_ipo_n43), .A (b[19]));
CLKBUF_X1 drc_ipo_c44 (.Z (drc_ipo_n44), .A (b[20]));
CLKBUF_X1 drc_ipo_c45 (.Z (drc_ipo_n45), .A (b[21]));
CLKBUF_X1 drc_ipo_c46 (.Z (drc_ipo_n46), .A (b[22]));
CLKBUF_X1 drc_ipo_c47 (.Z (drc_ipo_n47), .A (b[23]));
CLKBUF_X1 drc_ipo_c48 (.Z (drc_ipo_n48), .A (b[24]));
CLKBUF_X1 drc_ipo_c49 (.Z (drc_ipo_n49), .A (b[25]));
CLKBUF_X1 drc_ipo_c50 (.Z (drc_ipo_n50), .A (b[26]));
CLKBUF_X1 drc_ipo_c51 (.Z (drc_ipo_n51), .A (b[27]));
CLKBUF_X1 drc_ipo_c52 (.Z (drc_ipo_n52), .A (b[28]));
CLKBUF_X1 drc_ipo_c53 (.Z (drc_ipo_n53), .A (b[29]));
CLKBUF_X1 drc_ipo_c54 (.Z (drc_ipo_n54), .A (b[30]));
CLKBUF_X1 drc_ipo_c55 (.Z (drc_ipo_n55), .A (b[31]));
CLKBUF_X1 drc_ipo_c56 (.Z (drc_ipo_n56), .A (a[0]));
CLKBUF_X1 drc_ipo_c57 (.Z (drc_ipo_n57), .A (a[1]));
CLKBUF_X1 drc_ipo_c58 (.Z (drc_ipo_n58), .A (a[2]));
CLKBUF_X1 drc_ipo_c59 (.Z (drc_ipo_n59), .A (a[3]));
CLKBUF_X1 drc_ipo_c60 (.Z (drc_ipo_n60), .A (a[4]));
CLKBUF_X1 drc_ipo_c61 (.Z (drc_ipo_n61), .A (a[5]));
CLKBUF_X1 drc_ipo_c62 (.Z (drc_ipo_n62), .A (a[6]));
CLKBUF_X1 drc_ipo_c63 (.Z (drc_ipo_n63), .A (a[7]));
CLKBUF_X1 drc_ipo_c64 (.Z (drc_ipo_n64), .A (a[8]));
CLKBUF_X1 drc_ipo_c65 (.Z (drc_ipo_n65), .A (a[9]));
CLKBUF_X1 drc_ipo_c66 (.Z (drc_ipo_n66), .A (a[10]));
CLKBUF_X1 drc_ipo_c67 (.Z (drc_ipo_n67), .A (a[11]));
CLKBUF_X1 drc_ipo_c68 (.Z (drc_ipo_n68), .A (a[12]));
CLKBUF_X1 drc_ipo_c69 (.Z (drc_ipo_n69), .A (a[13]));
CLKBUF_X1 drc_ipo_c70 (.Z (drc_ipo_n70), .A (a[14]));
CLKBUF_X1 drc_ipo_c71 (.Z (drc_ipo_n71), .A (a[15]));
CLKBUF_X1 drc_ipo_c72 (.Z (drc_ipo_n72), .A (a[16]));
CLKBUF_X1 drc_ipo_c73 (.Z (drc_ipo_n73), .A (a[17]));
CLKBUF_X1 drc_ipo_c74 (.Z (drc_ipo_n74), .A (a[18]));
CLKBUF_X1 drc_ipo_c75 (.Z (drc_ipo_n75), .A (a[19]));
CLKBUF_X1 drc_ipo_c76 (.Z (drc_ipo_n76), .A (a[20]));
CLKBUF_X1 drc_ipo_c77 (.Z (drc_ipo_n77), .A (a[21]));
CLKBUF_X1 drc_ipo_c78 (.Z (drc_ipo_n78), .A (a[22]));
CLKBUF_X1 drc_ipo_c79 (.Z (drc_ipo_n79), .A (a[23]));
CLKBUF_X1 drc_ipo_c80 (.Z (drc_ipo_n80), .A (a[24]));
CLKBUF_X1 drc_ipo_c81 (.Z (drc_ipo_n81), .A (a[25]));
CLKBUF_X1 drc_ipo_c82 (.Z (drc_ipo_n82), .A (a[26]));
CLKBUF_X1 drc_ipo_c83 (.Z (drc_ipo_n83), .A (a[27]));
CLKBUF_X1 drc_ipo_c84 (.Z (drc_ipo_n84), .A (a[28]));
CLKBUF_X1 drc_ipo_c85 (.Z (drc_ipo_n85), .A (a[29]));
CLKBUF_X1 drc_ipo_c86 (.Z (drc_ipo_n86), .A (a[30]));
CLKBUF_X1 drc_ipo_c87 (.Z (drc_ipo_n87), .A (a[31]));
CLKBUF_X1 drc_ipo_c88 (.Z (drc_ipo_n88), .A (en));
BUF_X4 drc_ipo_c89 (.Z (drc_ipo_n89), .A (rst));
CLKBUF_X1 CTS_L3_c_tid0_290 (.Z (CTS_n_tid0_337), .A (CTS_n_tid0_338));
CLKBUF_X1 CTS_L2_c_tid0_293 (.Z (CTS_n_tid0_338), .A (CTS_n_tid0_339));
CLKBUF_X3 CTS_L3_c_tid1_211 (.Z (CTS_n_tid1_243), .A (CTS_n_tid1_244));
CLKBUF_X1 CLOCK_slh__c344 (.Z (CLOCK_slh__n436), .A (CLOCK_slh__n435));
CLKBUF_X3 CTS_L3_c_tid0_124 (.Z (CTS_n_tid0_128), .A (CTS_n_tid0_234));
CLKBUF_X1 CLOCK_slh__c345 (.Z (n_64_205), .A (CLOCK_slh__n436));
CLKBUF_X3 CTS_L1_c_tid0_294 (.Z (CTS_n_tid0_339), .A (clk));
CLKBUF_X1 CLOCK_slh__c348 (.Z (CLOCK_slh__n440), .A (CLOCK_slh__n439));
CLKBUF_X2 CTS_L3_c_tid0_131 (.Z (CTS_n_tid0_136), .A (CTS_n_tid0_234));
CLKBUF_X1 CLOCK_slh__c349 (.Z (n_64_225), .A (CLOCK_slh__n440));
CLKBUF_X1 CLOCK_slh__c352 (.Z (CLOCK_slh__n444), .A (CLOCK_slh__n443));
CLKBUF_X1 CLOCK_slh__c353 (.Z (n_64_222), .A (CLOCK_slh__n444));
CLKBUF_X1 CLOCK_slh__c336 (.Z (CLOCK_slh__n428), .A (CLOCK_slh__n427));
CLKBUF_X1 CLOCK_slh__c340 (.Z (CLOCK_slh__n432), .A (CLOCK_slh__n431));
CLKBUF_X1 CLOCK_slh__c337 (.Z (n_64_213), .A (CLOCK_slh__n428));
CLKBUF_X1 CLOCK_slh__c341 (.Z (n_64_214), .A (CLOCK_slh__n432));
CLKBUF_X1 CLOCK_slh__c356 (.Z (CLOCK_slh__n448), .A (CLOCK_slh__n447));
CLKBUF_X1 CLOCK_slh__c357 (.Z (n_64_204), .A (CLOCK_slh__n448));
CLKBUF_X1 CLOCK_slh__c360 (.Z (CLOCK_slh__n452), .A (CLOCK_slh__n451));
CLKBUF_X1 CLOCK_slh__c361 (.Z (n_64_221), .A (CLOCK_slh__n452));
CLKBUF_X1 CLOCK_slh__c364 (.Z (CLOCK_slh__n456), .A (CLOCK_slh__n455));
CLKBUF_X1 CLOCK_slh__c365 (.Z (n_64_218), .A (CLOCK_slh__n456));
CLKBUF_X1 CLOCK_slh__c368 (.Z (CLOCK_slh__n460), .A (CLOCK_slh__n459));
CLKBUF_X1 CLOCK_slh__c369 (.Z (n_64_217), .A (CLOCK_slh__n460));
CLKBUF_X1 CLOCK_slh__c372 (.Z (CLOCK_slh__n464), .A (CLOCK_slh__n463));
CLKBUF_X1 CLOCK_slh__c373 (.Z (n_64_229), .A (CLOCK_slh__n464));
CLKBUF_X1 CLOCK_slh__c376 (.Z (CLOCK_slh__n468), .A (CLOCK_slh__n467));
CLKBUF_X1 CLOCK_slh__c377 (.Z (n_64_226), .A (CLOCK_slh__n468));
CLKBUF_X1 CLOCK_slh__c380 (.Z (CLOCK_slh__n472), .A (CLOCK_slh__n471));
CLKBUF_X1 CLOCK_slh__c381 (.Z (n_64_220), .A (CLOCK_slh__n472));
CLKBUF_X1 CLOCK_slh__c384 (.Z (CLOCK_slh__n476), .A (CLOCK_slh__n475));
CLKBUF_X1 CLOCK_slh__c385 (.Z (n_64_212), .A (CLOCK_slh__n476));
CLKBUF_X1 CLOCK_slh__c388 (.Z (CLOCK_slh__n480), .A (CLOCK_slh__n479));
CLKBUF_X1 CLOCK_slh__c389 (.Z (n_64_224), .A (CLOCK_slh__n480));
CLKBUF_X1 CLOCK_slh__c392 (.Z (CLOCK_slh__n484), .A (CLOCK_slh__n483));
CLKBUF_X1 CLOCK_slh__c393 (.Z (n_64_202), .A (CLOCK_slh__n484));
CLKBUF_X1 CLOCK_slh__c396 (.Z (CLOCK_slh__n488), .A (CLOCK_slh__n487));
CLKBUF_X1 CLOCK_slh__c397 (.Z (n_64_298), .A (CLOCK_slh__n488));
CLKBUF_X1 CLOCK_slh__c400 (.Z (CLOCK_slh__n492), .A (CLOCK_slh__n491));
CLKBUF_X1 CLOCK_slh__c401 (.Z (n_64_228), .A (CLOCK_slh__n492));
CLKBUF_X1 CLOCK_slh__c404 (.Z (CLOCK_slh__n496), .A (CLOCK_slh__n495));
CLKBUF_X1 CLOCK_slh__c405 (.Z (n_64_216), .A (CLOCK_slh__n496));
CLKBUF_X1 CLOCK_slh__c408 (.Z (CLOCK_slh__n500), .A (CLOCK_slh__n499));
CLKBUF_X1 CLOCK_slh__c409 (.Z (n_64_223), .A (CLOCK_slh__n500));
CLKBUF_X1 CLOCK_slh__c412 (.Z (CLOCK_slh__n504), .A (CLOCK_slh__n503));
CLKBUF_X1 CLOCK_slh__c413 (.Z (n_64_203), .A (CLOCK_slh__n504));
CLKBUF_X1 CLOCK_slh__c416 (.Z (CLOCK_slh__n508), .A (CLOCK_slh__n507));
CLKBUF_X1 CLOCK_slh__c417 (.Z (n_64_209), .A (CLOCK_slh__n508));
CLKBUF_X1 CLOCK_slh__c420 (.Z (n_64_210), .A (CLOCK_slh__n511));
CLKBUF_X1 CLOCK_slh__c422 (.Z (n_64_227), .A (CLOCK_slh__n513));
CLKBUF_X1 CLOCK_slh__c424 (.Z (n_64_206), .A (CLOCK_slh__n515));
CLKBUF_X1 CLOCK_slh__c426 (.Z (n_64_219), .A (CLOCK_slh__n517));
CLKBUF_X1 CLOCK_slh__c428 (.Z (n_64_201), .A (CLOCK_slh__n519));
CLKBUF_X1 CLOCK_slh__c429 (.Z (n_64_208), .A (CLOCK_slh__n520));
CLKBUF_X1 CLOCK_slh__c430 (.Z (n_64_207), .A (CLOCK_slh__n521));
CLKBUF_X1 CLOCK_slh__c431 (.Z (n_64_211), .A (CLOCK_slh__n522));

endmodule //booth_multiplier


