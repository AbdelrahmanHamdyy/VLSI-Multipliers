/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 18:15:59 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3142015809 */

module buffer__0_65(clk, rst, D, Q);
   input clk;
   input rst;
   input [31:0]D;
   output [31:0]Q;

   wire n_0_0;

   DFF_X1 \Q_reg[31]  (.D(n_31), .CK(clk), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_30), .CK(clk), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_29), .CK(clk), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_28), .CK(clk), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_27), .CK(clk), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_26), .CK(clk), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_25), .CK(clk), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_24), .CK(clk), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_23), .CK(clk), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_22), .CK(clk), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_21), .CK(clk), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_20), .CK(clk), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_19), .CK(clk), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_18), .CK(clk), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_17), .CK(clk), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_16), .CK(clk), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(clk), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(clk), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(clk), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(clk), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(clk), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(clk), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(clk), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(clk), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(clk), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(clk), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(clk), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(clk), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(clk), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(clk), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(clk), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(clk), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_1 (.A1(n_0_0), .A2(D[0]), .ZN(n_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[1]), .ZN(n_1));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[2]), .ZN(n_2));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[3]), .ZN(n_3));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[4]), .ZN(n_4));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[5]), .ZN(n_5));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[6]), .ZN(n_6));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[7]), .ZN(n_7));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[8]), .ZN(n_8));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[9]), .ZN(n_9));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[10]), .ZN(n_10));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[11]), .ZN(n_11));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[12]), .ZN(n_12));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[13]), .ZN(n_13));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[14]), .ZN(n_14));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[15]), .ZN(n_15));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[16]), .ZN(n_16));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[17]), .ZN(n_17));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[18]), .ZN(n_18));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[19]), .ZN(n_19));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[20]), .ZN(n_20));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[21]), .ZN(n_21));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[22]), .ZN(n_22));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[23]), .ZN(n_23));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[24]), .ZN(n_24));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[25]), .ZN(n_25));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[26]), .ZN(n_26));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[27]), .ZN(n_27));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[28]), .ZN(n_28));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[29]), .ZN(n_29));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[30]), .ZN(n_30));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[31]), .ZN(n_31));
endmodule

module buffer(clk, rst, D, Q);
   input clk;
   input rst;
   input [31:0]D;
   output [31:0]Q;

   wire n_0_0;

   DFF_X1 \Q_reg[31]  (.D(n_31), .CK(clk), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_30), .CK(clk), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_29), .CK(clk), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_28), .CK(clk), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_27), .CK(clk), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_26), .CK(clk), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_25), .CK(clk), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_24), .CK(clk), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_23), .CK(clk), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_22), .CK(clk), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_21), .CK(clk), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_20), .CK(clk), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_19), .CK(clk), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_18), .CK(clk), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_17), .CK(clk), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_16), .CK(clk), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(clk), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(clk), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(clk), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(clk), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(clk), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(clk), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(clk), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(clk), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(clk), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(clk), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(clk), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(clk), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(clk), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(clk), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(clk), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(clk), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_1 (.A1(n_0_0), .A2(D[0]), .ZN(n_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[1]), .ZN(n_1));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[2]), .ZN(n_2));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[3]), .ZN(n_3));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[4]), .ZN(n_4));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[5]), .ZN(n_5));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[6]), .ZN(n_6));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[7]), .ZN(n_7));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[8]), .ZN(n_8));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[9]), .ZN(n_9));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[10]), .ZN(n_10));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[11]), .ZN(n_11));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[12]), .ZN(n_12));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[13]), .ZN(n_13));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[14]), .ZN(n_14));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[15]), .ZN(n_15));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[16]), .ZN(n_16));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[17]), .ZN(n_17));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[18]), .ZN(n_18));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[19]), .ZN(n_19));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[20]), .ZN(n_20));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[21]), .ZN(n_21));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[22]), .ZN(n_22));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[23]), .ZN(n_23));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[24]), .ZN(n_24));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[25]), .ZN(n_25));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[26]), .ZN(n_26));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[27]), .ZN(n_27));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[28]), .ZN(n_28));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[29]), .ZN(n_29));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[30]), .ZN(n_30));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[31]), .ZN(n_31));
endmodule

module datapath(b, a, p_0);
   input [31:0]b;
   input [31:0]a;
   output [63:0]p_0;

   HA_X1 i_1052 (.A(n_1030), .B(n_1045), .CO(n_1053), .S(n_1052));
   FA_X1 i_1067 (.A(n_1040), .B(n_1046), .CI(n_1063), .CO(n_1069), .S(n_1068));
   HA_X1 i_1068 (.A(n_1056), .B(n_1053), .CO(n_1071), .S(n_1070));
   FA_X1 i_1091 (.A(n_1081), .B(n_1074), .CI(n_1088), .CO(n_1095), .S(n_1094));
   HA_X1 i_1092 (.A(n_1071), .B(n_1069), .CO(n_1097), .S(n_1096));
   FA_X1 i_1115 (.A(n_1075), .B(n_1089), .CI(n_1113), .CO(n_1121), .S(n_1120));
   FA_X1 i_1116 (.A(n_1107), .B(n_1100), .CI(n_1097), .CO(n_1123), .S(n_1122));
   HA_X1 i_1117 (.A(n_1120), .B(n_1095), .CO(n_1125), .S(n_1124));
   FA_X1 i_1139 (.A(n_1108), .B(n_1101), .CI(n_1114), .CO(n_1148), .S(n_1147));
   FA_X1 i_1140 (.A(n_1142), .B(n_1135), .CI(n_1128), .CO(n_1150), .S(n_1149));
   FA_X1 i_1141 (.A(n_1147), .B(n_1121), .CI(n_1125), .CO(n_1152), .S(n_1151));
   HA_X1 i_1142 (.A(n_1123), .B(n_1149), .CO(n_1154), .S(n_1153));
   FA_X1 i_1172 (.A(n_1129), .B(n_1171), .CI(n_1164), .CO(n_1185), .S(n_1184));
   FA_X1 i_1173 (.A(n_1157), .B(n_1148), .CI(n_1178), .CO(n_1187), .S(n_1186));
   FA_X1 i_1174 (.A(n_1150), .B(n_1184), .CI(n_1186), .CO(n_1189), .S(n_1188));
   HA_X1 i_1175 (.A(n_1154), .B(n_1152), .CO(n_1191), .S(n_1190));
   FA_X1 i_1205 (.A(n_1165), .B(n_1158), .CI(n_1179), .CO(n_1222), .S(n_1221));
   FA_X1 i_1206 (.A(n_1214), .B(n_1208), .CI(n_1201), .CO(n_1224), .S(n_1223));
   FA_X1 i_1207 (.A(n_1194), .B(n_1221), .CI(n_1185), .CO(n_1226), .S(n_1225));
   FA_X1 i_1208 (.A(n_1187), .B(n_1223), .CI(n_1225), .CO(n_1228), .S(n_1227));
   HA_X1 i_1209 (.A(n_1191), .B(n_1189), .CO(n_1230), .S(n_1229));
   FA_X1 i_1238 (.A(n_1209), .B(n_1202), .CI(n_1195), .CO(n_1260), .S(n_1259));
   FA_X1 i_1239 (.A(n_1215), .B(n_1254), .CI(n_1247), .CO(n_1262), .S(n_1261));
   FA_X1 i_1240 (.A(n_1240), .B(n_1233), .CI(n_1222), .CO(n_1264), .S(n_1263));
   FA_X1 i_1241 (.A(n_1259), .B(n_1224), .CI(n_1226), .CO(n_1266), .S(n_1265));
   FA_X1 i_1242 (.A(n_1263), .B(n_1261), .CI(n_1265), .CO(n_1268), .S(n_1267));
   HA_X1 i_1243 (.A(n_1230), .B(n_1228), .CO(n_1270), .S(n_1269));
   FA_X1 i_1280 (.A(n_1241), .B(n_1234), .CI(n_1260), .CO(n_1308), .S(n_1307));
   FA_X1 i_1281 (.A(n_1294), .B(n_1287), .CI(n_1280), .CO(n_1310), .S(n_1309));
   FA_X1 i_1282 (.A(n_1273), .B(n_1307), .CI(n_1301), .CO(n_1312), .S(n_1311));
   FA_X1 i_1283 (.A(n_1262), .B(n_1264), .CI(n_1309), .CO(n_1314), .S(n_1313));
   FA_X1 i_1284 (.A(n_1266), .B(n_1311), .CI(n_1313), .CO(n_1316), .S(n_1315));
   HA_X1 i_1285 (.A(n_1268), .B(n_1270), .CO(n_1318), .S(n_1317));
   FA_X1 i_1322 (.A(n_1288), .B(n_1281), .CI(n_1274), .CO(n_1356), .S(n_1355));
   FA_X1 i_1323 (.A(n_1302), .B(n_1348), .CI(n_1342), .CO(n_1358), .S(n_1357));
   FA_X1 i_1324 (.A(n_1335), .B(n_1328), .CI(n_1321), .CO(n_1360), .S(n_1359));
   FA_X1 i_1325 (.A(n_1308), .B(n_1355), .CI(n_1310), .CO(n_1362), .S(n_1361));
   FA_X1 i_1326 (.A(n_1312), .B(n_1359), .CI(n_1357), .CO(n_1364), .S(n_1363));
   FA_X1 i_1327 (.A(n_1361), .B(n_1314), .CI(n_1316), .CO(n_1366), .S(n_1365));
   HA_X1 i_1328 (.A(n_1363), .B(n_1318), .CO(n_1368), .S(n_1367));
   FA_X1 i_1364 (.A(n_1343), .B(n_1336), .CI(n_1329), .CO(n_1405), .S(n_1404));
   FA_X1 i_1365 (.A(n_1322), .B(n_1356), .CI(n_1349), .CO(n_1407), .S(n_1406));
   FA_X1 i_1366 (.A(n_1399), .B(n_1392), .CI(n_1385), .CO(n_1409), .S(n_1408));
   FA_X1 i_1367 (.A(n_1378), .B(n_1371), .CI(n_1404), .CO(n_1411), .S(n_1410));
   FA_X1 i_1368 (.A(n_1360), .B(n_1358), .CI(n_1406), .CO(n_1413), .S(n_1412));
   FA_X1 i_1369 (.A(n_1362), .B(n_1410), .CI(n_1408), .CO(n_1415), .S(n_1414));
   FA_X1 i_1370 (.A(n_1412), .B(n_1364), .CI(n_1414), .CO(n_1417), .S(n_1416));
   HA_X1 i_1371 (.A(n_1366), .B(n_1368), .CO(n_1419), .S(n_1418));
   FA_X1 i_1415 (.A(n_1386), .B(n_1379), .CI(n_1372), .CO(n_1464), .S(n_1463));
   FA_X1 i_1416 (.A(n_1405), .B(n_1450), .CI(n_1443), .CO(n_1466), .S(n_1465));
   FA_X1 i_1417 (.A(n_1436), .B(n_1429), .CI(n_1422), .CO(n_1468), .S(n_1467));
   FA_X1 i_1418 (.A(n_1407), .B(n_1463), .CI(n_1457), .CO(n_1470), .S(n_1469));
   FA_X1 i_1419 (.A(n_1409), .B(n_1411), .CI(n_1467), .CO(n_1472), .S(n_1471));
   FA_X1 i_1420 (.A(n_1465), .B(n_1413), .CI(n_1469), .CO(n_1474), .S(n_1473));
   FA_X1 i_1421 (.A(n_1415), .B(n_1471), .CI(n_1473), .CO(n_1476), .S(n_1475));
   HA_X1 i_1422 (.A(n_1417), .B(n_1419), .CO(n_1478), .S(n_1477));
   FA_X1 i_1466 (.A(n_1444), .B(n_1437), .CI(n_1430), .CO(n_1523), .S(n_1522));
   FA_X1 i_1467 (.A(n_1423), .B(n_1464), .CI(n_1458), .CO(n_1525), .S(n_1524));
   FA_X1 i_1468 (.A(n_1515), .B(n_1509), .CI(n_1502), .CO(n_1527), .S(n_1526));
   FA_X1 i_1469 (.A(n_1495), .B(n_1488), .CI(n_1481), .CO(n_1529), .S(n_1528));
   FA_X1 i_1470 (.A(n_1522), .B(n_1468), .CI(n_1466), .CO(n_1531), .S(n_1530));
   FA_X1 i_1471 (.A(n_1524), .B(n_1470), .CI(n_1528), .CO(n_1533), .S(n_1532));
   FA_X1 i_1472 (.A(n_1526), .B(n_1530), .CI(n_1472), .CO(n_1535), .S(n_1534));
   FA_X1 i_1473 (.A(n_1532), .B(n_1474), .CI(n_1534), .CO(n_1537), .S(n_1536));
   HA_X1 i_1474 (.A(n_1476), .B(n_1478), .CO(n_1539), .S(n_1538));
   FA_X1 i_1517 (.A(n_1510), .B(n_1503), .CI(n_1496), .CO(n_1583), .S(n_1582));
   FA_X1 i_1518 (.A(n_1489), .B(n_1482), .CI(n_1523), .CO(n_1585), .S(n_1584));
   FA_X1 i_1519 (.A(n_1516), .B(n_1577), .CI(n_1570), .CO(n_1587), .S(n_1586));
   FA_X1 i_1520 (.A(n_1563), .B(n_1556), .CI(n_1549), .CO(n_1589), .S(n_1588));
   FA_X1 i_1521 (.A(n_1542), .B(n_1525), .CI(n_1584), .CO(n_1591), .S(n_1590));
   FA_X1 i_1522 (.A(n_1582), .B(n_1529), .CI(n_1527), .CO(n_1593), .S(n_1592));
   FA_X1 i_1523 (.A(n_1531), .B(n_1588), .CI(n_1586), .CO(n_1595), .S(n_1594));
   FA_X1 i_1524 (.A(n_1590), .B(n_1592), .CI(n_1533), .CO(n_1597), .S(n_1596));
   FA_X1 i_1525 (.A(n_1535), .B(n_1594), .CI(n_1596), .CO(n_1599), .S(n_1598));
   HA_X1 i_1526 (.A(n_1537), .B(n_1539), .CO(n_1601), .S(n_1600));
   FA_X1 i_1577 (.A(n_1564), .B(n_1557), .CI(n_1550), .CO(n_1653), .S(n_1652));
   FA_X1 i_1578 (.A(n_1543), .B(n_1583), .CI(n_1639), .CO(n_1655), .S(n_1654));
   FA_X1 i_1579 (.A(n_1632), .B(n_1625), .CI(n_1618), .CO(n_1657), .S(n_1656));
   FA_X1 i_1580 (.A(n_1611), .B(n_1604), .CI(n_1585), .CO(n_1659), .S(n_1658));
   FA_X1 i_1581 (.A(n_1652), .B(n_1646), .CI(n_1589), .CO(n_1661), .S(n_1660));
   FA_X1 i_1582 (.A(n_1587), .B(n_1654), .CI(n_1593), .CO(n_1663), .S(n_1662));
   FA_X1 i_1583 (.A(n_1591), .B(n_1658), .CI(n_1656), .CO(n_1665), .S(n_1664));
   FA_X1 i_1584 (.A(n_1660), .B(n_1595), .CI(n_1662), .CO(n_1667), .S(n_1666));
   FA_X1 i_1585 (.A(n_1597), .B(n_1664), .CI(n_1666), .CO(n_1669), .S(n_1668));
   HA_X1 i_1586 (.A(n_1599), .B(n_1668), .CO(n_1671), .S(n_1670));
   FA_X1 i_1637 (.A(n_1633), .B(n_1626), .CI(n_1619), .CO(n_1723), .S(n_1722));
   FA_X1 i_1638 (.A(n_1612), .B(n_1605), .CI(n_1653), .CO(n_1725), .S(n_1724));
   FA_X1 i_1639 (.A(n_1647), .B(n_1715), .CI(n_1709), .CO(n_1727), .S(n_1726));
   FA_X1 i_1640 (.A(n_1702), .B(n_1695), .CI(n_1688), .CO(n_1729), .S(n_1728));
   FA_X1 i_1641 (.A(n_1681), .B(n_1674), .CI(n_1724), .CO(n_1731), .S(n_1730));
   FA_X1 i_1642 (.A(n_1722), .B(n_1657), .CI(n_1655), .CO(n_1733), .S(n_1732));
   FA_X1 i_1643 (.A(n_1659), .B(n_1661), .CI(n_1730), .CO(n_1735), .S(n_1734));
   FA_X1 i_1644 (.A(n_1728), .B(n_1726), .CI(n_1663), .CO(n_1737), .S(n_1736));
   FA_X1 i_1645 (.A(n_1732), .B(n_1665), .CI(n_1734), .CO(n_1739), .S(n_1738));
   FA_X1 i_1646 (.A(n_1736), .B(n_1667), .CI(n_1738), .CO(n_1741), .S(n_1740));
   HA_X1 i_1647 (.A(n_1669), .B(n_1740), .CO(n_1743), .S(n_1742));
   FA_X1 i_1697 (.A(n_1710), .B(n_1703), .CI(n_1696), .CO(n_1794), .S(n_1793));
   FA_X1 i_1698 (.A(n_1689), .B(n_1682), .CI(n_1675), .CO(n_1796), .S(n_1795));
   FA_X1 i_1699 (.A(n_1723), .B(n_1716), .CI(n_1788), .CO(n_1798), .S(n_1797));
   FA_X1 i_1700 (.A(n_1781), .B(n_1774), .CI(n_1767), .CO(n_1800), .S(n_1799));
   FA_X1 i_1701 (.A(n_1760), .B(n_1753), .CI(n_1746), .CO(n_1802), .S(n_1801));
   FA_X1 i_1702 (.A(n_1725), .B(n_1795), .CI(n_1793), .CO(n_1804), .S(n_1803));
   FA_X1 i_1703 (.A(n_1729), .B(n_1727), .CI(n_1797), .CO(n_1806), .S(n_1805));
   FA_X1 i_1704 (.A(n_1733), .B(n_1731), .CI(n_1801), .CO(n_1808), .S(n_1807));
   FA_X1 i_1705 (.A(n_1799), .B(n_1805), .CI(n_1803), .CO(n_1810), .S(n_1809));
   FA_X1 i_1706 (.A(n_1735), .B(n_1737), .CI(n_1807), .CO(n_1812), .S(n_1811));
   FA_X1 i_1707 (.A(n_1739), .B(n_1809), .CI(n_1811), .CO(n_1814), .S(n_1813));
   HA_X1 i_1708 (.A(n_1741), .B(n_1743), .CO(n_1816), .S(n_1815));
   FA_X1 i_1766 (.A(n_1775), .B(n_1768), .CI(n_1761), .CO(n_1875), .S(n_1874));
   FA_X1 i_1767 (.A(n_1754), .B(n_1747), .CI(n_1796), .CO(n_1877), .S(n_1876));
   FA_X1 i_1768 (.A(n_1794), .B(n_1861), .CI(n_1854), .CO(n_1879), .S(n_1878));
   FA_X1 i_1769 (.A(n_1847), .B(n_1840), .CI(n_1833), .CO(n_1881), .S(n_1880));
   FA_X1 i_1770 (.A(n_1826), .B(n_1819), .CI(n_1876), .CO(n_1883), .S(n_1882));
   FA_X1 i_1771 (.A(n_1874), .B(n_1868), .CI(n_1802), .CO(n_1885), .S(n_1884));
   FA_X1 i_1772 (.A(n_1800), .B(n_1798), .CI(n_1804), .CO(n_1887), .S(n_1886));
   FA_X1 i_1773 (.A(n_1882), .B(n_1880), .CI(n_1878), .CO(n_1889), .S(n_1888));
   FA_X1 i_1774 (.A(n_1806), .B(n_1886), .CI(n_1884), .CO(n_1891), .S(n_1890));
   FA_X1 i_1775 (.A(n_1808), .B(n_1810), .CI(n_1888), .CO(n_1893), .S(n_1892));
   FA_X1 i_1776 (.A(n_1812), .B(n_1890), .CI(n_1892), .CO(n_1895), .S(n_1894));
   HA_X1 i_1777 (.A(n_1814), .B(n_1894), .CO(n_1897), .S(n_1896));
   FA_X1 i_1835 (.A(n_1855), .B(n_1848), .CI(n_1841), .CO(n_1956), .S(n_1955));
   FA_X1 i_1836 (.A(n_1834), .B(n_1827), .CI(n_1820), .CO(n_1958), .S(n_1957));
   FA_X1 i_1837 (.A(n_1875), .B(n_1869), .CI(n_1948), .CO(n_1960), .S(n_1959));
   FA_X1 i_1838 (.A(n_1942), .B(n_1935), .CI(n_1928), .CO(n_1962), .S(n_1961));
   FA_X1 i_1839 (.A(n_1921), .B(n_1914), .CI(n_1907), .CO(n_1964), .S(n_1963));
   FA_X1 i_1840 (.A(n_1900), .B(n_1877), .CI(n_1957), .CO(n_1966), .S(n_1965));
   FA_X1 i_1841 (.A(n_1955), .B(n_1881), .CI(n_1879), .CO(n_1968), .S(n_1967));
   FA_X1 i_1842 (.A(n_1959), .B(n_1885), .CI(n_1883), .CO(n_1970), .S(n_1969));
   FA_X1 i_1843 (.A(n_1963), .B(n_1961), .CI(n_1965), .CO(n_1972), .S(n_1971));
   FA_X1 i_1844 (.A(n_1887), .B(n_1967), .CI(n_1889), .CO(n_1974), .S(n_1973));
   FA_X1 i_1845 (.A(n_1969), .B(n_1891), .CI(n_1971), .CO(n_1976), .S(n_1975));
   FA_X1 i_1846 (.A(n_1973), .B(n_1893), .CI(n_1975), .CO(n_1978), .S(n_1977));
   HA_X1 i_1847 (.A(n_1895), .B(n_1977), .CO(n_1980), .S(n_1979));
   FA_X1 i_1904 (.A(n_1943), .B(n_1936), .CI(n_1929), .CO(n_2038), .S(n_2037));
   FA_X1 i_1905 (.A(n_1922), .B(n_1915), .CI(n_1908), .CO(n_2040), .S(n_2039));
   FA_X1 i_1906 (.A(n_1901), .B(n_1958), .CI(n_1956), .CO(n_2042), .S(n_2041));
   FA_X1 i_1907 (.A(n_1949), .B(n_2032), .CI(n_2025), .CO(n_2044), .S(n_2043));
   FA_X1 i_1908 (.A(n_2018), .B(n_2011), .CI(n_2004), .CO(n_2046), .S(n_2045));
   FA_X1 i_1909 (.A(n_1997), .B(n_1990), .CI(n_1983), .CO(n_2048), .S(n_2047));
   FA_X1 i_1910 (.A(n_2039), .B(n_2037), .CI(n_1964), .CO(n_2050), .S(n_2049));
   FA_X1 i_1911 (.A(n_1962), .B(n_1960), .CI(n_2041), .CO(n_2052), .S(n_2051));
   FA_X1 i_1912 (.A(n_1968), .B(n_1966), .CI(n_2047), .CO(n_2054), .S(n_2053));
   FA_X1 i_1913 (.A(n_2045), .B(n_2043), .CI(n_1970), .CO(n_2056), .S(n_2055));
   FA_X1 i_1914 (.A(n_2051), .B(n_2049), .CI(n_1972), .CO(n_2058), .S(n_2057));
   FA_X1 i_1915 (.A(n_2053), .B(n_1974), .CI(n_2055), .CO(n_2060), .S(n_2059));
   FA_X1 i_1916 (.A(n_2057), .B(n_1976), .CI(n_2059), .CO(n_2062), .S(n_2061));
   HA_X1 i_1917 (.A(n_1978), .B(n_2061), .CO(n_2064), .S(n_2063));
   FA_X1 i_1982 (.A(n_2019), .B(n_2012), .CI(n_2005), .CO(n_2130), .S(n_2129));
   FA_X1 i_1983 (.A(n_1998), .B(n_1991), .CI(n_1984), .CO(n_2132), .S(n_2131));
   FA_X1 i_1984 (.A(n_2040), .B(n_2038), .CI(n_2116), .CO(n_2134), .S(n_2133));
   FA_X1 i_1985 (.A(n_2109), .B(n_2102), .CI(n_2095), .CO(n_2136), .S(n_2135));
   FA_X1 i_1986 (.A(n_2088), .B(n_2081), .CI(n_2074), .CO(n_2138), .S(n_2137));
   FA_X1 i_1987 (.A(n_2067), .B(n_2042), .CI(n_2131), .CO(n_2140), .S(n_2139));
   FA_X1 i_1988 (.A(n_2129), .B(n_2123), .CI(n_2048), .CO(n_2142), .S(n_2141));
   FA_X1 i_1989 (.A(n_2046), .B(n_2044), .CI(n_2133), .CO(n_2144), .S(n_2143));
   FA_X1 i_1990 (.A(n_2050), .B(n_2137), .CI(n_2135), .CO(n_2146), .S(n_2145));
   FA_X1 i_1991 (.A(n_2139), .B(n_2052), .CI(n_2143), .CO(n_2148), .S(n_2147));
   FA_X1 i_1992 (.A(n_2141), .B(n_2054), .CI(n_2056), .CO(n_2150), .S(n_2149));
   FA_X1 i_1993 (.A(n_2058), .B(n_2145), .CI(n_2147), .CO(n_2152), .S(n_2151));
   FA_X1 i_1994 (.A(n_2149), .B(n_2060), .CI(n_2151), .CO(n_2154), .S(n_2153));
   HA_X1 i_1995 (.A(n_2062), .B(n_2153), .CO(n_2156), .S(n_2155));
   FA_X1 i_2060 (.A(n_2110), .B(n_2103), .CI(n_2096), .CO(n_2222), .S(n_2221));
   FA_X1 i_2061 (.A(n_2089), .B(n_2082), .CI(n_2075), .CO(n_2224), .S(n_2223));
   FA_X1 i_2062 (.A(n_2068), .B(n_2132), .CI(n_2130), .CO(n_2226), .S(n_2225));
   FA_X1 i_2063 (.A(n_2124), .B(n_2214), .CI(n_2208), .CO(n_2228), .S(n_2227));
   FA_X1 i_2064 (.A(n_2201), .B(n_2194), .CI(n_2187), .CO(n_2230), .S(n_2229));
   FA_X1 i_2065 (.A(n_2180), .B(n_2173), .CI(n_2166), .CO(n_2232), .S(n_2231));
   FA_X1 i_2066 (.A(n_2159), .B(n_2223), .CI(n_2221), .CO(n_2234), .S(n_2233));
   FA_X1 i_2067 (.A(n_2138), .B(n_2136), .CI(n_2134), .CO(n_2236), .S(n_2235));
   FA_X1 i_2068 (.A(n_2225), .B(n_2142), .CI(n_2140), .CO(n_2238), .S(n_2237));
   FA_X1 i_2069 (.A(n_2231), .B(n_2229), .CI(n_2227), .CO(n_2240), .S(n_2239));
   FA_X1 i_2070 (.A(n_2144), .B(n_2235), .CI(n_2233), .CO(n_2242), .S(n_2241));
   FA_X1 i_2071 (.A(n_2146), .B(n_2237), .CI(n_2148), .CO(n_2244), .S(n_2243));
   FA_X1 i_2072 (.A(n_2150), .B(n_2239), .CI(n_2241), .CO(n_2246), .S(n_2245));
   FA_X1 i_2073 (.A(n_2152), .B(n_2243), .CI(n_2245), .CO(n_2248), .S(n_2247));
   HA_X1 i_2074 (.A(n_2154), .B(n_2156), .CO(n_2250), .S(n_2249));
   FA_X1 i_2138 (.A(n_2209), .B(n_2202), .CI(n_2195), .CO(n_2315), .S(n_2314));
   FA_X1 i_2139 (.A(n_2188), .B(n_2181), .CI(n_2174), .CO(n_2317), .S(n_2316));
   FA_X1 i_2140 (.A(n_2167), .B(n_2160), .CI(n_2224), .CO(n_2319), .S(n_2318));
   FA_X1 i_2141 (.A(n_2222), .B(n_2215), .CI(n_2309), .CO(n_2321), .S(n_2320));
   FA_X1 i_2142 (.A(n_2302), .B(n_2295), .CI(n_2288), .CO(n_2323), .S(n_2322));
   FA_X1 i_2143 (.A(n_2281), .B(n_2274), .CI(n_2267), .CO(n_2325), .S(n_2324));
   FA_X1 i_2144 (.A(n_2260), .B(n_2253), .CI(n_2226), .CO(n_2327), .S(n_2326));
   FA_X1 i_2145 (.A(n_2318), .B(n_2316), .CI(n_2314), .CO(n_2329), .S(n_2328));
   FA_X1 i_2146 (.A(n_2232), .B(n_2230), .CI(n_2228), .CO(n_2331), .S(n_2330));
   FA_X1 i_2147 (.A(n_2320), .B(n_2236), .CI(n_2234), .CO(n_2333), .S(n_2332));
   FA_X1 i_2148 (.A(n_2326), .B(n_2324), .CI(n_2322), .CO(n_2335), .S(n_2334));
   FA_X1 i_2149 (.A(n_2238), .B(n_2330), .CI(n_2328), .CO(n_2337), .S(n_2336));
   FA_X1 i_2150 (.A(n_2240), .B(n_2332), .CI(n_2242), .CO(n_2339), .S(n_2338));
   FA_X1 i_2151 (.A(n_2334), .B(n_2244), .CI(n_2336), .CO(n_2341), .S(n_2340));
   FA_X1 i_2152 (.A(n_2338), .B(n_2246), .CI(n_2340), .CO(n_2343), .S(n_2342));
   HA_X1 i_2153 (.A(n_2248), .B(n_2342), .CO(n_2345), .S(n_2344));
   FA_X1 i_2225 (.A(n_2296), .B(n_2289), .CI(n_2282), .CO(n_2418), .S(n_2417));
   FA_X1 i_2226 (.A(n_2275), .B(n_2268), .CI(n_2261), .CO(n_2420), .S(n_2419));
   FA_X1 i_2227 (.A(n_2254), .B(n_2317), .CI(n_2315), .CO(n_2422), .S(n_2421));
   FA_X1 i_2228 (.A(n_2404), .B(n_2397), .CI(n_2390), .CO(n_2424), .S(n_2423));
   FA_X1 i_2229 (.A(n_2383), .B(n_2376), .CI(n_2369), .CO(n_2426), .S(n_2425));
   FA_X1 i_2230 (.A(n_2362), .B(n_2355), .CI(n_2348), .CO(n_2428), .S(n_2427));
   FA_X1 i_2231 (.A(n_2319), .B(n_2419), .CI(n_2417), .CO(n_2430), .S(n_2429));
   FA_X1 i_2232 (.A(n_2411), .B(n_2325), .CI(n_2323), .CO(n_2432), .S(n_2431));
   FA_X1 i_2233 (.A(n_2321), .B(n_2327), .CI(n_2421), .CO(n_2434), .S(n_2433));
   FA_X1 i_2234 (.A(n_2331), .B(n_2329), .CI(n_2427), .CO(n_2436), .S(n_2435));
   FA_X1 i_2235 (.A(n_2425), .B(n_2423), .CI(n_2333), .CO(n_2438), .S(n_2437));
   FA_X1 i_2236 (.A(n_2431), .B(n_2429), .CI(n_2335), .CO(n_2440), .S(n_2439));
   FA_X1 i_2237 (.A(n_2433), .B(n_2435), .CI(n_2337), .CO(n_2442), .S(n_2441));
   FA_X1 i_2238 (.A(n_2437), .B(n_2339), .CI(n_2439), .CO(n_2444), .S(n_2443));
   FA_X1 i_2239 (.A(n_2441), .B(n_2341), .CI(n_2443), .CO(n_2446), .S(n_2445));
   HA_X1 i_2240 (.A(n_2343), .B(n_2445), .CO(n_2448), .S(n_2447));
   FA_X1 i_2312 (.A(n_2398), .B(n_2391), .CI(n_2384), .CO(n_2521), .S(n_2520));
   FA_X1 i_2313 (.A(n_2377), .B(n_2370), .CI(n_2363), .CO(n_2523), .S(n_2522));
   FA_X1 i_2314 (.A(n_2356), .B(n_2349), .CI(n_2420), .CO(n_2525), .S(n_2524));
   FA_X1 i_2315 (.A(n_2418), .B(n_2412), .CI(n_2513), .CO(n_2527), .S(n_2526));
   FA_X1 i_2316 (.A(n_2507), .B(n_2500), .CI(n_2493), .CO(n_2529), .S(n_2528));
   FA_X1 i_2317 (.A(n_2486), .B(n_2479), .CI(n_2472), .CO(n_2531), .S(n_2530));
   FA_X1 i_2318 (.A(n_2465), .B(n_2458), .CI(n_2451), .CO(n_2533), .S(n_2532));
   FA_X1 i_2319 (.A(n_2422), .B(n_2524), .CI(n_2522), .CO(n_2535), .S(n_2534));
   FA_X1 i_2320 (.A(n_2520), .B(n_2428), .CI(n_2426), .CO(n_2537), .S(n_2536));
   FA_X1 i_2321 (.A(n_2424), .B(n_2526), .CI(n_2432), .CO(n_2539), .S(n_2538));
   FA_X1 i_2322 (.A(n_2430), .B(n_2532), .CI(n_2530), .CO(n_2541), .S(n_2540));
   FA_X1 i_2323 (.A(n_2528), .B(n_2434), .CI(n_2536), .CO(n_2543), .S(n_2542));
   FA_X1 i_2324 (.A(n_2534), .B(n_2436), .CI(n_2438), .CO(n_2545), .S(n_2544));
   FA_X1 i_2325 (.A(n_2538), .B(n_2440), .CI(n_2540), .CO(n_2547), .S(n_2546));
   FA_X1 i_2326 (.A(n_2542), .B(n_2442), .CI(n_2544), .CO(n_2549), .S(n_2548));
   FA_X1 i_2327 (.A(n_2546), .B(n_2444), .CI(n_2548), .CO(n_2551), .S(n_2550));
   HA_X1 i_2328 (.A(n_2446), .B(n_2550), .CO(n_2553), .S(n_2552));
   FA_X1 i_2399 (.A(n_2508), .B(n_2501), .CI(n_2494), .CO(n_2625), .S(n_2624));
   FA_X1 i_2400 (.A(n_2487), .B(n_2480), .CI(n_2473), .CO(n_2627), .S(n_2626));
   FA_X1 i_2401 (.A(n_2466), .B(n_2459), .CI(n_2452), .CO(n_2629), .S(n_2628));
   FA_X1 i_2402 (.A(n_2523), .B(n_2521), .CI(n_2514), .CO(n_2631), .S(n_2630));
   FA_X1 i_2403 (.A(n_2619), .B(n_2612), .CI(n_2605), .CO(n_2633), .S(n_2632));
   FA_X1 i_2404 (.A(n_2598), .B(n_2591), .CI(n_2584), .CO(n_2635), .S(n_2634));
   FA_X1 i_2405 (.A(n_2577), .B(n_2570), .CI(n_2563), .CO(n_2637), .S(n_2636));
   FA_X1 i_2406 (.A(n_2556), .B(n_2525), .CI(n_2628), .CO(n_2639), .S(n_2638));
   FA_X1 i_2407 (.A(n_2626), .B(n_2624), .CI(n_2533), .CO(n_2641), .S(n_2640));
   FA_X1 i_2408 (.A(n_2531), .B(n_2529), .CI(n_2527), .CO(n_2643), .S(n_2642));
   FA_X1 i_2409 (.A(n_2630), .B(n_2537), .CI(n_2535), .CO(n_2645), .S(n_2644));
   FA_X1 i_2410 (.A(n_2636), .B(n_2634), .CI(n_2632), .CO(n_2647), .S(n_2646));
   FA_X1 i_2411 (.A(n_2638), .B(n_2539), .CI(n_2642), .CO(n_2649), .S(n_2648));
   FA_X1 i_2412 (.A(n_2640), .B(n_2541), .CI(n_2644), .CO(n_2651), .S(n_2650));
   FA_X1 i_2413 (.A(n_2543), .B(n_2545), .CI(n_2646), .CO(n_2653), .S(n_2652));
   FA_X1 i_2414 (.A(n_2648), .B(n_2650), .CI(n_2547), .CO(n_2655), .S(n_2654));
   FA_X1 i_2415 (.A(n_2549), .B(n_2652), .CI(n_2654), .CO(n_2657), .S(n_2656));
   HA_X1 i_2416 (.A(n_2551), .B(n_2656), .CO(n_2659), .S(n_2658));
   FA_X1 i_2495 (.A(n_2606), .B(n_2599), .CI(n_2592), .CO(n_2739), .S(n_2738));
   FA_X1 i_2496 (.A(n_2585), .B(n_2578), .CI(n_2571), .CO(n_2741), .S(n_2740));
   FA_X1 i_2497 (.A(n_2564), .B(n_2557), .CI(n_2629), .CO(n_2743), .S(n_2742));
   FA_X1 i_2498 (.A(n_2627), .B(n_2625), .CI(n_2725), .CO(n_2745), .S(n_2744));
   FA_X1 i_2499 (.A(n_2718), .B(n_2711), .CI(n_2704), .CO(n_2747), .S(n_2746));
   FA_X1 i_2500 (.A(n_2697), .B(n_2690), .CI(n_2683), .CO(n_2749), .S(n_2748));
   FA_X1 i_2501 (.A(n_2676), .B(n_2669), .CI(n_2662), .CO(n_2751), .S(n_2750));
   FA_X1 i_2502 (.A(n_2631), .B(n_2742), .CI(n_2740), .CO(n_2753), .S(n_2752));
   FA_X1 i_2503 (.A(n_2738), .B(n_2732), .CI(n_2637), .CO(n_2755), .S(n_2754));
   FA_X1 i_2504 (.A(n_2635), .B(n_2633), .CI(n_2744), .CO(n_2757), .S(n_2756));
   FA_X1 i_2505 (.A(n_2643), .B(n_2641), .CI(n_2639), .CO(n_2759), .S(n_2758));
   FA_X1 i_2506 (.A(n_2750), .B(n_2748), .CI(n_2746), .CO(n_2761), .S(n_2760));
   FA_X1 i_2507 (.A(n_2645), .B(n_2756), .CI(n_2754), .CO(n_2763), .S(n_2762));
   FA_X1 i_2508 (.A(n_2752), .B(n_2647), .CI(n_2758), .CO(n_2765), .S(n_2764));
   FA_X1 i_2509 (.A(n_2649), .B(n_2760), .CI(n_2651), .CO(n_2767), .S(n_2766));
   FA_X1 i_2510 (.A(n_2764), .B(n_2762), .CI(n_2653), .CO(n_2769), .S(n_2768));
   FA_X1 i_2511 (.A(n_2655), .B(n_2766), .CI(n_2768), .CO(n_2771), .S(n_2770));
   HA_X1 i_2512 (.A(n_2657), .B(n_2770), .CO(n_2773), .S(n_2772));
   FA_X1 i_2591 (.A(n_2719), .B(n_2712), .CI(n_2705), .CO(n_2853), .S(n_2852));
   FA_X1 i_2592 (.A(n_2698), .B(n_2691), .CI(n_2684), .CO(n_2855), .S(n_2854));
   FA_X1 i_2593 (.A(n_2677), .B(n_2670), .CI(n_2663), .CO(n_2857), .S(n_2856));
   FA_X1 i_2594 (.A(n_2741), .B(n_2739), .CI(n_2733), .CO(n_2859), .S(n_2858));
   FA_X1 i_2595 (.A(n_2845), .B(n_2839), .CI(n_2832), .CO(n_2861), .S(n_2860));
   FA_X1 i_2596 (.A(n_2825), .B(n_2818), .CI(n_2811), .CO(n_2863), .S(n_2862));
   FA_X1 i_2597 (.A(n_2804), .B(n_2797), .CI(n_2790), .CO(n_2865), .S(n_2864));
   FA_X1 i_2598 (.A(n_2783), .B(n_2776), .CI(n_2743), .CO(n_2867), .S(n_2866));
   FA_X1 i_2599 (.A(n_2856), .B(n_2854), .CI(n_2852), .CO(n_2869), .S(n_2868));
   FA_X1 i_2600 (.A(n_2751), .B(n_2749), .CI(n_2747), .CO(n_2871), .S(n_2870));
   FA_X1 i_2601 (.A(n_2745), .B(n_2858), .CI(n_2755), .CO(n_2873), .S(n_2872));
   FA_X1 i_2602 (.A(n_2753), .B(n_2866), .CI(n_2864), .CO(n_2875), .S(n_2874));
   FA_X1 i_2603 (.A(n_2862), .B(n_2860), .CI(n_2759), .CO(n_2877), .S(n_2876));
   FA_X1 i_2604 (.A(n_2757), .B(n_2870), .CI(n_2868), .CO(n_2879), .S(n_2878));
   FA_X1 i_2605 (.A(n_2761), .B(n_2872), .CI(n_2763), .CO(n_2881), .S(n_2880));
   FA_X1 i_2606 (.A(n_2876), .B(n_2874), .CI(n_2765), .CO(n_2883), .S(n_2882));
   FA_X1 i_2607 (.A(n_2878), .B(n_2767), .CI(n_2880), .CO(n_2885), .S(n_2884));
   FA_X1 i_2608 (.A(n_2769), .B(n_2882), .CI(n_2884), .CO(n_2887), .S(n_2886));
   HA_X1 i_2609 (.A(n_2771), .B(n_2886), .CO(n_2889), .S(n_2888));
   FA_X1 i_2688 (.A(n_2826), .B(n_2819), .CI(n_2812), .CO(n_2969), .S(n_2968));
   FA_X1 i_2689 (.A(n_2805), .B(n_2798), .CI(n_2791), .CO(n_2971), .S(n_2970));
   FA_X1 i_2690 (.A(n_2784), .B(n_2777), .CI(n_2857), .CO(n_2973), .S(n_2972));
   FA_X1 i_2691 (.A(n_2855), .B(n_2853), .CI(n_2846), .CO(n_2975), .S(n_2974));
   FA_X1 i_2692 (.A(n_2955), .B(n_2948), .CI(n_2941), .CO(n_2977), .S(n_2976));
   FA_X1 i_2693 (.A(n_2934), .B(n_2927), .CI(n_2920), .CO(n_2979), .S(n_2978));
   FA_X1 i_2694 (.A(n_2913), .B(n_2906), .CI(n_2899), .CO(n_2981), .S(n_2980));
   FA_X1 i_2695 (.A(n_2892), .B(n_2859), .CI(n_2972), .CO(n_2983), .S(n_2982));
   FA_X1 i_2696 (.A(n_2970), .B(n_2968), .CI(n_2962), .CO(n_2985), .S(n_2984));
   FA_X1 i_2697 (.A(n_2865), .B(n_2863), .CI(n_2861), .CO(n_2987), .S(n_2986));
   FA_X1 i_2698 (.A(n_2867), .B(n_2974), .CI(n_2871), .CO(n_2989), .S(n_2988));
   FA_X1 i_2699 (.A(n_2869), .B(n_2980), .CI(n_2978), .CO(n_2991), .S(n_2990));
   FA_X1 i_2700 (.A(n_2976), .B(n_2982), .CI(n_2873), .CO(n_2993), .S(n_2992));
   FA_X1 i_2701 (.A(n_2986), .B(n_2984), .CI(n_2875), .CO(n_2995), .S(n_2994));
   FA_X1 i_2702 (.A(n_2877), .B(n_2988), .CI(n_2879), .CO(n_2997), .S(n_2996));
   FA_X1 i_2703 (.A(n_2990), .B(n_2992), .CI(n_2881), .CO(n_2999), .S(n_2998));
   FA_X1 i_2704 (.A(n_2994), .B(n_2883), .CI(n_2996), .CO(n_3001), .S(n_3000));
   FA_X1 i_2705 (.A(n_2998), .B(n_2885), .CI(n_3000), .CO(n_3003), .S(n_3002));
   HA_X1 i_2706 (.A(n_2887), .B(n_3002), .CO(n_3005), .S(n_3004));
   FA_X1 i_2777 (.A(n_2956), .B(n_2949), .CI(n_2942), .CO(n_3077), .S(n_3076));
   FA_X1 i_2778 (.A(n_2935), .B(n_2928), .CI(n_2921), .CO(n_3079), .S(n_3078));
   FA_X1 i_2779 (.A(n_2914), .B(n_2907), .CI(n_2900), .CO(n_3081), .S(n_3080));
   FA_X1 i_2780 (.A(n_2893), .B(n_2971), .CI(n_2969), .CO(n_3083), .S(n_3082));
   FA_X1 i_2781 (.A(n_2963), .B(n_3071), .CI(n_3064), .CO(n_3085), .S(n_3084));
   FA_X1 i_2782 (.A(n_3057), .B(n_3050), .CI(n_3043), .CO(n_3087), .S(n_3086));
   FA_X1 i_2783 (.A(n_3036), .B(n_3029), .CI(n_3022), .CO(n_3089), .S(n_3088));
   FA_X1 i_2784 (.A(n_3015), .B(n_3008), .CI(n_2975), .CO(n_3091), .S(n_3090));
   FA_X1 i_2785 (.A(n_2973), .B(n_3080), .CI(n_3078), .CO(n_3093), .S(n_3092));
   FA_X1 i_2786 (.A(n_3076), .B(n_2981), .CI(n_2979), .CO(n_3095), .S(n_3094));
   FA_X1 i_2787 (.A(n_2977), .B(n_3082), .CI(n_2987), .CO(n_3097), .S(n_3096));
   FA_X1 i_2788 (.A(n_2985), .B(n_2983), .CI(n_3090), .CO(n_3099), .S(n_3098));
   FA_X1 i_2789 (.A(n_3088), .B(n_3086), .CI(n_3084), .CO(n_3101), .S(n_3100));
   FA_X1 i_2790 (.A(n_2989), .B(n_3094), .CI(n_3092), .CO(n_3103), .S(n_3102));
   FA_X1 i_2791 (.A(n_2991), .B(n_2993), .CI(n_3098), .CO(n_3105), .S(n_3104));
   FA_X1 i_2792 (.A(n_3096), .B(n_2995), .CI(n_3100), .CO(n_3107), .S(n_3106));
   FA_X1 i_2793 (.A(n_2997), .B(n_3102), .CI(n_3104), .CO(n_3109), .S(n_3108));
   FA_X1 i_2794 (.A(n_2999), .B(n_3106), .CI(n_3001), .CO(n_3111), .S(n_3110));
   FA_X1 i_2795 (.A(n_3108), .B(n_3110), .CI(n_3003), .CO(n_3113), .S(n_3112));
   FA_X1 i_2867 (.A(n_3065), .B(n_3058), .CI(n_3051), .CO(n_3186), .S(n_3185));
   FA_X1 i_2868 (.A(n_3044), .B(n_3037), .CI(n_3030), .CO(n_3188), .S(n_3187));
   FA_X1 i_2869 (.A(n_3023), .B(n_3016), .CI(n_3009), .CO(n_3190), .S(n_3189));
   FA_X1 i_2870 (.A(n_3081), .B(n_3079), .CI(n_3077), .CO(n_3192), .S(n_3191));
   FA_X1 i_2871 (.A(n_3178), .B(n_3172), .CI(n_3165), .CO(n_3194), .S(n_3193));
   FA_X1 i_2872 (.A(n_3158), .B(n_3151), .CI(n_3144), .CO(n_3196), .S(n_3195));
   FA_X1 i_2873 (.A(n_3137), .B(n_3130), .CI(n_3123), .CO(n_3198), .S(n_3197));
   FA_X1 i_2874 (.A(n_3116), .B(n_3083), .CI(n_3189), .CO(n_3200), .S(n_3199));
   FA_X1 i_2875 (.A(n_3187), .B(n_3185), .CI(n_3089), .CO(n_3202), .S(n_3201));
   FA_X1 i_2876 (.A(n_3087), .B(n_3085), .CI(n_3091), .CO(n_3204), .S(n_3203));
   FA_X1 i_2877 (.A(n_3191), .B(n_3095), .CI(n_3093), .CO(n_3206), .S(n_3205));
   FA_X1 i_2878 (.A(n_3197), .B(n_3195), .CI(n_3193), .CO(n_3208), .S(n_3207));
   FA_X1 i_2879 (.A(n_3199), .B(n_3097), .CI(n_3203), .CO(n_3210), .S(n_3209));
   FA_X1 i_2880 (.A(n_3201), .B(n_3101), .CI(n_3099), .CO(n_3212), .S(n_3211));
   FA_X1 i_2881 (.A(n_3205), .B(n_3103), .CI(n_3207), .CO(n_3214), .S(n_3213));
   FA_X1 i_2882 (.A(n_3209), .B(n_3105), .CI(n_3211), .CO(n_3216), .S(n_3215));
   FA_X1 i_2883 (.A(n_3107), .B(n_3213), .CI(n_3109), .CO(n_3218), .S(n_3217));
   FA_X1 i_2884 (.A(n_3215), .B(n_3111), .CI(n_3217), .CO(n_3220), .S(n_3219));
   FA_X1 i_2956 (.A(n_3159), .B(n_3152), .CI(n_3145), .CO(n_3293), .S(n_3292));
   FA_X1 i_2957 (.A(n_3138), .B(n_3131), .CI(n_3124), .CO(n_3295), .S(n_3294));
   FA_X1 i_2958 (.A(n_3117), .B(n_3190), .CI(n_3188), .CO(n_3297), .S(n_3296));
   FA_X1 i_2959 (.A(n_3186), .B(n_3179), .CI(n_3279), .CO(n_3299), .S(n_3298));
   FA_X1 i_2960 (.A(n_3272), .B(n_3265), .CI(n_3258), .CO(n_3301), .S(n_3300));
   FA_X1 i_2961 (.A(n_3251), .B(n_3244), .CI(n_3237), .CO(n_3303), .S(n_3302));
   FA_X1 i_2962 (.A(n_3230), .B(n_3223), .CI(n_3192), .CO(n_3305), .S(n_3304));
   FA_X1 i_2963 (.A(n_3294), .B(n_3292), .CI(n_3286), .CO(n_3307), .S(n_3306));
   FA_X1 i_2964 (.A(n_3198), .B(n_3196), .CI(n_3194), .CO(n_3309), .S(n_3308));
   FA_X1 i_2965 (.A(n_3298), .B(n_3296), .CI(n_3202), .CO(n_3311), .S(n_3310));
   FA_X1 i_2966 (.A(n_3200), .B(n_3204), .CI(n_3304), .CO(n_3313), .S(n_3312));
   FA_X1 i_2967 (.A(n_3302), .B(n_3300), .CI(n_3206), .CO(n_3315), .S(n_3314));
   FA_X1 i_2968 (.A(n_3308), .B(n_3306), .CI(n_3208), .CO(n_3317), .S(n_3316));
   FA_X1 i_2969 (.A(n_3310), .B(n_3212), .CI(n_3210), .CO(n_3319), .S(n_3318));
   FA_X1 i_2970 (.A(n_3312), .B(n_3314), .CI(n_3316), .CO(n_3321), .S(n_3320));
   FA_X1 i_2971 (.A(n_3214), .B(n_3318), .CI(n_3216), .CO(n_3323), .S(n_3322));
   FA_X1 i_2972 (.A(n_3320), .B(n_3218), .CI(n_3322), .CO(n_3325), .S(n_3324));
   FA_X1 i_3036 (.A(n_3280), .B(n_3273), .CI(n_3266), .CO(n_3390), .S(n_3389));
   FA_X1 i_3037 (.A(n_3259), .B(n_3252), .CI(n_3245), .CO(n_3392), .S(n_3391));
   FA_X1 i_3038 (.A(n_3238), .B(n_3231), .CI(n_3224), .CO(n_3394), .S(n_3393));
   FA_X1 i_3039 (.A(n_3295), .B(n_3293), .CI(n_3287), .CO(n_3396), .S(n_3395));
   FA_X1 i_3040 (.A(n_3384), .B(n_3377), .CI(n_3370), .CO(n_3398), .S(n_3397));
   FA_X1 i_3041 (.A(n_3363), .B(n_3356), .CI(n_3349), .CO(n_3400), .S(n_3399));
   FA_X1 i_3042 (.A(n_3342), .B(n_3335), .CI(n_3328), .CO(n_3402), .S(n_3401));
   FA_X1 i_3043 (.A(n_3297), .B(n_3393), .CI(n_3391), .CO(n_3404), .S(n_3403));
   FA_X1 i_3044 (.A(n_3389), .B(n_3303), .CI(n_3301), .CO(n_3406), .S(n_3405));
   FA_X1 i_3045 (.A(n_3299), .B(n_3305), .CI(n_3395), .CO(n_3408), .S(n_3407));
   FA_X1 i_3046 (.A(n_3309), .B(n_3307), .CI(n_3401), .CO(n_3410), .S(n_3409));
   FA_X1 i_3047 (.A(n_3399), .B(n_3397), .CI(n_3311), .CO(n_3412), .S(n_3411));
   FA_X1 i_3048 (.A(n_3405), .B(n_3403), .CI(n_3313), .CO(n_3414), .S(n_3413));
   FA_X1 i_3049 (.A(n_3407), .B(n_3315), .CI(n_3409), .CO(n_3416), .S(n_3415));
   FA_X1 i_3050 (.A(n_3317), .B(n_3411), .CI(n_3319), .CO(n_3418), .S(n_3417));
   FA_X1 i_3051 (.A(n_3413), .B(n_3415), .CI(n_3321), .CO(n_3420), .S(n_3419));
   FA_X1 i_3052 (.A(n_3417), .B(n_3323), .CI(n_3419), .CO(n_3422), .S(n_3421));
   FA_X1 i_3117 (.A(n_3378), .B(n_3371), .CI(n_3364), .CO(n_3488), .S(n_3487));
   FA_X1 i_3118 (.A(n_3357), .B(n_3350), .CI(n_3343), .CO(n_3490), .S(n_3489));
   FA_X1 i_3119 (.A(n_3336), .B(n_3329), .CI(n_3394), .CO(n_3492), .S(n_3491));
   FA_X1 i_3120 (.A(n_3392), .B(n_3390), .CI(n_3480), .CO(n_3494), .S(n_3493));
   FA_X1 i_3121 (.A(n_3474), .B(n_3467), .CI(n_3460), .CO(n_3496), .S(n_3495));
   FA_X1 i_3122 (.A(n_3453), .B(n_3446), .CI(n_3439), .CO(n_3498), .S(n_3497));
   FA_X1 i_3123 (.A(n_3432), .B(n_3425), .CI(n_3396), .CO(n_3500), .S(n_3499));
   FA_X1 i_3124 (.A(n_3491), .B(n_3489), .CI(n_3487), .CO(n_3502), .S(n_3501));
   FA_X1 i_3125 (.A(n_3402), .B(n_3400), .CI(n_3398), .CO(n_3504), .S(n_3503));
   FA_X1 i_3126 (.A(n_3493), .B(n_3406), .CI(n_3404), .CO(n_3506), .S(n_3505));
   FA_X1 i_3127 (.A(n_3499), .B(n_3497), .CI(n_3495), .CO(n_3508), .S(n_3507));
   FA_X1 i_3128 (.A(n_3408), .B(n_3503), .CI(n_3501), .CO(n_3510), .S(n_3509));
   FA_X1 i_3129 (.A(n_3410), .B(n_3412), .CI(n_3505), .CO(n_3512), .S(n_3511));
   FA_X1 i_3130 (.A(n_3414), .B(n_3507), .CI(n_3416), .CO(n_3514), .S(n_3513));
   FA_X1 i_3131 (.A(n_3509), .B(n_3511), .CI(n_3418), .CO(n_3516), .S(n_3515));
   FA_X1 i_3132 (.A(n_3513), .B(n_3420), .CI(n_3515), .CO(n_3518), .S(n_3517));
   FA_X1 i_3197 (.A(n_3461), .B(n_3454), .CI(n_3447), .CO(n_3584), .S(n_3583));
   FA_X1 i_3198 (.A(n_3440), .B(n_3433), .CI(n_3426), .CO(n_3586), .S(n_3585));
   FA_X1 i_3199 (.A(n_3490), .B(n_3488), .CI(n_3481), .CO(n_3588), .S(n_3587));
   FA_X1 i_3200 (.A(n_3570), .B(n_3563), .CI(n_3556), .CO(n_3590), .S(n_3589));
   FA_X1 i_3201 (.A(n_3549), .B(n_3542), .CI(n_3535), .CO(n_3592), .S(n_3591));
   FA_X1 i_3202 (.A(n_3528), .B(n_3521), .CI(n_3492), .CO(n_3594), .S(n_3593));
   FA_X1 i_3203 (.A(n_3585), .B(n_3583), .CI(n_3577), .CO(n_3596), .S(n_3595));
   FA_X1 i_3204 (.A(n_3498), .B(n_3496), .CI(n_3494), .CO(n_3598), .S(n_3597));
   FA_X1 i_3205 (.A(n_3500), .B(n_3587), .CI(n_3504), .CO(n_3600), .S(n_3599));
   FA_X1 i_3206 (.A(n_3502), .B(n_3593), .CI(n_3591), .CO(n_3602), .S(n_3601));
   FA_X1 i_3207 (.A(n_3589), .B(n_3506), .CI(n_3597), .CO(n_3604), .S(n_3603));
   FA_X1 i_3208 (.A(n_3595), .B(n_3508), .CI(n_3599), .CO(n_3606), .S(n_3605));
   FA_X1 i_3209 (.A(n_3510), .B(n_3601), .CI(n_3603), .CO(n_3608), .S(n_3607));
   FA_X1 i_3210 (.A(n_3512), .B(n_3605), .CI(n_3514), .CO(n_3610), .S(n_3609));
   FA_X1 i_3211 (.A(n_3516), .B(n_3607), .CI(n_3609), .CO(n_3612), .S(n_3611));
   FA_X1 i_3268 (.A(n_3571), .B(n_3564), .CI(n_3557), .CO(n_3670), .S(n_3669));
   FA_X1 i_3269 (.A(n_3550), .B(n_3543), .CI(n_3536), .CO(n_3672), .S(n_3671));
   FA_X1 i_3270 (.A(n_3529), .B(n_3522), .CI(n_3586), .CO(n_3674), .S(n_3673));
   FA_X1 i_3271 (.A(n_3584), .B(n_3578), .CI(n_3664), .CO(n_3676), .S(n_3675));
   FA_X1 i_3272 (.A(n_3657), .B(n_3650), .CI(n_3643), .CO(n_3678), .S(n_3677));
   FA_X1 i_3273 (.A(n_3636), .B(n_3629), .CI(n_3622), .CO(n_3680), .S(n_3679));
   FA_X1 i_3274 (.A(n_3615), .B(n_3588), .CI(n_3673), .CO(n_3682), .S(n_3681));
   FA_X1 i_3275 (.A(n_3671), .B(n_3669), .CI(n_3592), .CO(n_3684), .S(n_3683));
   FA_X1 i_3276 (.A(n_3590), .B(n_3594), .CI(n_3675), .CO(n_3686), .S(n_3685));
   FA_X1 i_3277 (.A(n_3598), .B(n_3596), .CI(n_3679), .CO(n_3688), .S(n_3687));
   FA_X1 i_3278 (.A(n_3677), .B(n_3681), .CI(n_3600), .CO(n_3690), .S(n_3689));
   FA_X1 i_3279 (.A(n_3683), .B(n_3602), .CI(n_3685), .CO(n_3692), .S(n_3691));
   FA_X1 i_3280 (.A(n_3687), .B(n_3604), .CI(n_3689), .CO(n_3694), .S(n_3693));
   FA_X1 i_3281 (.A(n_3606), .B(n_3691), .CI(n_3608), .CO(n_3696), .S(n_3695));
   FA_X1 i_3282 (.A(n_3693), .B(n_3610), .CI(n_3695), .CO(n_3698), .S(n_3697));
   FA_X1 i_3340 (.A(n_3658), .B(n_3651), .CI(n_3644), .CO(n_3757), .S(n_3756));
   FA_X1 i_3341 (.A(n_3637), .B(n_3630), .CI(n_3623), .CO(n_3759), .S(n_3758));
   FA_X1 i_3342 (.A(n_3616), .B(n_3672), .CI(n_3670), .CO(n_3761), .S(n_3760));
   FA_X1 i_3343 (.A(n_3749), .B(n_3743), .CI(n_3736), .CO(n_3763), .S(n_3762));
   FA_X1 i_3344 (.A(n_3729), .B(n_3722), .CI(n_3715), .CO(n_3765), .S(n_3764));
   FA_X1 i_3345 (.A(n_3708), .B(n_3701), .CI(n_3674), .CO(n_3767), .S(n_3766));
   FA_X1 i_3346 (.A(n_3758), .B(n_3756), .CI(n_3680), .CO(n_3769), .S(n_3768));
   FA_X1 i_3347 (.A(n_3678), .B(n_3676), .CI(n_3760), .CO(n_3771), .S(n_3770));
   FA_X1 i_3348 (.A(n_3684), .B(n_3682), .CI(n_3766), .CO(n_3773), .S(n_3772));
   FA_X1 i_3349 (.A(n_3764), .B(n_3762), .CI(n_3686), .CO(n_3775), .S(n_3774));
   FA_X1 i_3350 (.A(n_3770), .B(n_3768), .CI(n_3688), .CO(n_3777), .S(n_3776));
   FA_X1 i_3351 (.A(n_3690), .B(n_3772), .CI(n_3692), .CO(n_3779), .S(n_3778));
   FA_X1 i_3352 (.A(n_3774), .B(n_3776), .CI(n_3694), .CO(n_3781), .S(n_3780));
   FA_X1 i_3353 (.A(n_3778), .B(n_3696), .CI(n_3780), .CO(n_3783), .S(n_3782));
   FA_X1 i_3411 (.A(n_3730), .B(n_3723), .CI(n_3716), .CO(n_1), .S(n_0));
   FA_X1 i_3412 (.A(n_3709), .B(n_3702), .CI(n_3759), .CO(n_3), .S(n_2));
   FA_X1 i_3413 (.A(n_3757), .B(n_3750), .CI(n_491), .CO(n_5), .S(n_4));
   FA_X1 i_3414 (.A(n_490), .B(n_3814), .CI(n_3807), .CO(n_7), .S(n_6));
   FA_X1 i_3415 (.A(n_3800), .B(n_3793), .CI(n_3786), .CO(n_9), .S(n_8));
   FA_X1 i_3416 (.A(n_3761), .B(n_2), .CI(n_0), .CO(n_11), .S(n_10));
   FA_X1 i_3417 (.A(n_489), .B(n_3765), .CI(n_3763), .CO(n_13), .S(n_12));
   FA_X1 i_3418 (.A(n_3767), .B(n_4), .CI(n_3769), .CO(n_15), .S(n_14));
   FA_X1 i_3419 (.A(n_8), .B(n_6), .CI(n_3771), .CO(n_17), .S(n_16));
   FA_X1 i_3420 (.A(n_12), .B(n_10), .CI(n_3773), .CO(n_19), .S(n_18));
   FA_X1 i_3421 (.A(n_3775), .B(n_14), .CI(n_3777), .CO(n_21), .S(n_20));
   FA_X1 i_3422 (.A(n_16), .B(n_3779), .CI(n_18), .CO(n_23), .S(n_22));
   FA_X1 i_3423 (.A(n_20), .B(n_3781), .CI(n_22), .CO(n_25), .S(n_24));
   FA_X1 i_3473 (.A(n_488), .B(n_487), .CI(n_3815), .CO(n_27), .S(n_26));
   FA_X1 i_3474 (.A(n_3808), .B(n_3801), .CI(n_3794), .CO(n_29), .S(n_28));
   FA_X1 i_3475 (.A(n_3787), .B(n_1), .CI(n_486), .CO(n_31), .S(n_30));
   FA_X1 i_3476 (.A(n_485), .B(n_484), .CI(n_483), .CO(n_33), .S(n_32));
   FA_X1 i_3477 (.A(n_482), .B(n_481), .CI(n_480), .CO(n_35), .S(n_34));
   FA_X1 i_3478 (.A(n_479), .B(n_3), .CI(n_28), .CO(n_37), .S(n_36));
   FA_X1 i_3479 (.A(n_26), .B(n_9), .CI(n_7), .CO(n_39), .S(n_38));
   FA_X1 i_3480 (.A(n_5), .B(n_30), .CI(n_13), .CO(n_41), .S(n_40));
   FA_X1 i_3481 (.A(n_11), .B(n_34), .CI(n_32), .CO(n_43), .S(n_42));
   FA_X1 i_3482 (.A(n_36), .B(n_15), .CI(n_38), .CO(n_45), .S(n_44));
   FA_X1 i_3483 (.A(n_17), .B(n_40), .CI(n_19), .CO(n_47), .S(n_46));
   FA_X1 i_3484 (.A(n_42), .B(n_44), .CI(n_21), .CO(n_49), .S(n_48));
   FA_X1 i_3485 (.A(n_46), .B(n_23), .CI(n_48), .CO(n_51), .S(n_50));
   FA_X1 i_3536 (.A(n_478), .B(n_477), .CI(n_476), .CO(n_53), .S(n_52));
   FA_X1 i_3537 (.A(n_475), .B(n_474), .CI(n_473), .CO(n_55), .S(n_54));
   FA_X1 i_3538 (.A(n_29), .B(n_27), .CI(n_472), .CO(n_57), .S(n_56));
   FA_X1 i_3539 (.A(n_471), .B(n_470), .CI(n_469), .CO(n_59), .S(n_58));
   FA_X1 i_3540 (.A(n_468), .B(n_467), .CI(n_466), .CO(n_61), .S(n_60));
   FA_X1 i_3541 (.A(n_31), .B(n_54), .CI(n_52), .CO(n_63), .S(n_62));
   FA_X1 i_3542 (.A(n_35), .B(n_33), .CI(n_56), .CO(n_65), .S(n_64));
   FA_X1 i_3543 (.A(n_39), .B(n_37), .CI(n_60), .CO(n_67), .S(n_66));
   FA_X1 i_3544 (.A(n_58), .B(n_41), .CI(n_64), .CO(n_69), .S(n_68));
   FA_X1 i_3545 (.A(n_62), .B(n_43), .CI(n_66), .CO(n_71), .S(n_70));
   FA_X1 i_3546 (.A(n_45), .B(n_68), .CI(n_47), .CO(n_73), .S(n_72));
   FA_X1 i_3547 (.A(n_70), .B(n_49), .CI(n_72), .CO(n_75), .S(n_74));
   FA_X1 i_3598 (.A(n_465), .B(n_464), .CI(n_463), .CO(n_77), .S(n_76));
   FA_X1 i_3599 (.A(n_462), .B(n_55), .CI(n_53), .CO(n_79), .S(n_78));
   FA_X1 i_3600 (.A(n_461), .B(n_460), .CI(n_459), .CO(n_81), .S(n_80));
   FA_X1 i_3601 (.A(n_458), .B(n_457), .CI(n_456), .CO(n_83), .S(n_82));
   FA_X1 i_3602 (.A(n_455), .B(n_76), .CI(n_454), .CO(n_85), .S(n_84));
   FA_X1 i_3603 (.A(n_61), .B(n_59), .CI(n_57), .CO(n_87), .S(n_86));
   FA_X1 i_3604 (.A(n_78), .B(n_63), .CI(n_82), .CO(n_89), .S(n_88));
   FA_X1 i_3605 (.A(n_80), .B(n_65), .CI(n_86), .CO(n_91), .S(n_90));
   FA_X1 i_3606 (.A(n_84), .B(n_67), .CI(n_88), .CO(n_93), .S(n_92));
   FA_X1 i_3607 (.A(n_69), .B(n_90), .CI(n_71), .CO(n_95), .S(n_94));
   FA_X1 i_3608 (.A(n_92), .B(n_73), .CI(n_94), .CO(n_97), .S(n_96));
   FA_X1 i_3651 (.A(n_453), .B(n_452), .CI(n_451), .CO(n_99), .S(n_98));
   FA_X1 i_3652 (.A(n_450), .B(n_449), .CI(n_448), .CO(n_101), .S(n_100));
   FA_X1 i_3653 (.A(n_77), .B(n_447), .CI(n_446), .CO(n_103), .S(n_102));
   FA_X1 i_3654 (.A(n_445), .B(n_444), .CI(n_443), .CO(n_105), .S(n_104));
   FA_X1 i_3655 (.A(n_442), .B(n_441), .CI(n_79), .CO(n_107), .S(n_106));
   FA_X1 i_3656 (.A(n_100), .B(n_98), .CI(n_83), .CO(n_109), .S(n_108));
   FA_X1 i_3657 (.A(n_81), .B(n_102), .CI(n_87), .CO(n_111), .S(n_110));
   FA_X1 i_3658 (.A(n_85), .B(n_106), .CI(n_104), .CO(n_113), .S(n_112));
   FA_X1 i_3659 (.A(n_108), .B(n_89), .CI(n_110), .CO(n_115), .S(n_114));
   FA_X1 i_3660 (.A(n_91), .B(n_112), .CI(n_93), .CO(n_117), .S(n_116));
   FA_X1 i_3661 (.A(n_114), .B(n_95), .CI(n_116), .CO(n_119), .S(n_118));
   FA_X1 i_3705 (.A(n_440), .B(n_439), .CI(n_438), .CO(n_121), .S(n_120));
   FA_X1 i_3706 (.A(n_437), .B(n_436), .CI(n_101), .CO(n_123), .S(n_122));
   FA_X1 i_3707 (.A(n_99), .B(n_435), .CI(n_434), .CO(n_125), .S(n_124));
   FA_X1 i_3708 (.A(n_433), .B(n_432), .CI(n_431), .CO(n_127), .S(n_126));
   FA_X1 i_3709 (.A(n_430), .B(n_122), .CI(n_120), .CO(n_129), .S(n_128));
   FA_X1 i_3710 (.A(n_105), .B(n_103), .CI(n_107), .CO(n_131), .S(n_130));
   FA_X1 i_3711 (.A(n_109), .B(n_126), .CI(n_124), .CO(n_133), .S(n_132));
   FA_X1 i_3712 (.A(n_111), .B(n_130), .CI(n_128), .CO(n_135), .S(n_134));
   FA_X1 i_3713 (.A(n_113), .B(n_132), .CI(n_115), .CO(n_137), .S(n_136));
   FA_X1 i_3714 (.A(n_134), .B(n_117), .CI(n_136), .CO(n_139), .S(n_138));
   FA_X1 i_3758 (.A(n_429), .B(n_428), .CI(n_427), .CO(n_141), .S(n_140));
   FA_X1 i_3759 (.A(n_121), .B(n_426), .CI(n_425), .CO(n_143), .S(n_142));
   FA_X1 i_3760 (.A(n_424), .B(n_423), .CI(n_422), .CO(n_145), .S(n_144));
   FA_X1 i_3761 (.A(n_421), .B(n_123), .CI(n_140), .CO(n_147), .S(n_146));
   FA_X1 i_3762 (.A(n_420), .B(n_127), .CI(n_125), .CO(n_149), .S(n_148));
   FA_X1 i_3763 (.A(n_142), .B(n_129), .CI(n_131), .CO(n_151), .S(n_150));
   FA_X1 i_3764 (.A(n_144), .B(n_146), .CI(n_148), .CO(n_153), .S(n_152));
   FA_X1 i_3765 (.A(n_133), .B(n_150), .CI(n_135), .CO(n_155), .S(n_154));
   FA_X1 i_3766 (.A(n_152), .B(n_137), .CI(n_154), .CO(n_157), .S(n_156));
   FA_X1 i_3802 (.A(n_419), .B(n_418), .CI(n_417), .CO(n_159), .S(n_158));
   FA_X1 i_3803 (.A(n_416), .B(n_415), .CI(n_141), .CO(n_161), .S(n_160));
   FA_X1 i_3804 (.A(n_414), .B(n_413), .CI(n_412), .CO(n_163), .S(n_162));
   FA_X1 i_3805 (.A(n_411), .B(n_410), .CI(n_409), .CO(n_165), .S(n_164));
   FA_X1 i_3806 (.A(n_160), .B(n_158), .CI(n_145), .CO(n_167), .S(n_166));
   FA_X1 i_3807 (.A(n_143), .B(n_149), .CI(n_147), .CO(n_169), .S(n_168));
   FA_X1 i_3808 (.A(n_164), .B(n_162), .CI(n_151), .CO(n_171), .S(n_170));
   FA_X1 i_3809 (.A(n_166), .B(n_168), .CI(n_153), .CO(n_173), .S(n_172));
   FA_X1 i_3810 (.A(n_170), .B(n_155), .CI(n_172), .CO(n_175), .S(n_174));
   FA_X1 i_3847 (.A(n_408), .B(n_407), .CI(n_406), .CO(n_177), .S(n_176));
   FA_X1 i_3848 (.A(n_405), .B(n_159), .CI(n_404), .CO(n_179), .S(n_178));
   FA_X1 i_3849 (.A(n_403), .B(n_402), .CI(n_401), .CO(n_181), .S(n_180));
   FA_X1 i_3850 (.A(n_400), .B(n_161), .CI(n_176), .CO(n_183), .S(n_182));
   FA_X1 i_3851 (.A(n_165), .B(n_163), .CI(n_178), .CO(n_185), .S(n_184));
   FA_X1 i_3852 (.A(n_167), .B(n_180), .CI(n_182), .CO(n_187), .S(n_186));
   FA_X1 i_3853 (.A(n_169), .B(n_184), .CI(n_171), .CO(n_189), .S(n_188));
   FA_X1 i_3854 (.A(n_186), .B(n_173), .CI(n_188), .CO(n_191), .S(n_190));
   FA_X1 i_3891 (.A(n_399), .B(n_398), .CI(n_177), .CO(n_193), .S(n_192));
   FA_X1 i_3892 (.A(n_397), .B(n_396), .CI(n_395), .CO(n_195), .S(n_194));
   FA_X1 i_3893 (.A(n_394), .B(n_393), .CI(n_192), .CO(n_197), .S(n_196));
   FA_X1 i_3894 (.A(n_392), .B(n_181), .CI(n_179), .CO(n_199), .S(n_198));
   FA_X1 i_3895 (.A(n_183), .B(n_196), .CI(n_194), .CO(n_201), .S(n_200));
   FA_X1 i_3896 (.A(n_185), .B(n_198), .CI(n_187), .CO(n_203), .S(n_202));
   FA_X1 i_3897 (.A(n_189), .B(n_200), .CI(n_202), .CO(n_205), .S(n_204));
   FA_X1 i_3926 (.A(n_391), .B(n_390), .CI(n_389), .CO(n_207), .S(n_206));
   FA_X1 i_3927 (.A(n_388), .B(n_387), .CI(n_386), .CO(n_209), .S(n_208));
   FA_X1 i_3928 (.A(n_385), .B(n_384), .CI(n_383), .CO(n_211), .S(n_210));
   FA_X1 i_3929 (.A(n_193), .B(n_206), .CI(n_195), .CO(n_213), .S(n_212));
   FA_X1 i_3930 (.A(n_208), .B(n_199), .CI(n_197), .CO(n_215), .S(n_214));
   FA_X1 i_3931 (.A(n_210), .B(n_212), .CI(n_201), .CO(n_217), .S(n_216));
   FA_X1 i_3932 (.A(n_214), .B(n_203), .CI(n_216), .CO(n_219), .S(n_218));
   FA_X1 i_3962 (.A(n_382), .B(n_381), .CI(n_380), .CO(n_221), .S(n_220));
   FA_X1 i_3963 (.A(n_207), .B(n_379), .CI(n_377), .CO(n_223), .S(n_222));
   FA_X1 i_3964 (.A(n_376), .B(n_375), .CI(n_220), .CO(n_225), .S(n_224));
   FA_X1 i_3965 (.A(n_211), .B(n_209), .CI(n_213), .CO(n_227), .S(n_226));
   FA_X1 i_3966 (.A(n_224), .B(n_222), .CI(n_215), .CO(n_229), .S(n_228));
   FA_X1 i_3967 (.A(n_226), .B(n_217), .CI(n_228), .CO(n_231), .S(n_230));
   FA_X1 i_3997 (.A(n_374), .B(n_221), .CI(n_378), .CO(n_233), .S(n_232));
   FA_X1 i_3998 (.A(n_373), .B(n_372), .CI(n_371), .CO(n_235), .S(n_234));
   FA_X1 i_3999 (.A(n_370), .B(n_223), .CI(n_232), .CO(n_237), .S(n_236));
   FA_X1 i_4000 (.A(n_225), .B(n_234), .CI(n_227), .CO(n_239), .S(n_238));
   FA_X1 i_4001 (.A(n_236), .B(n_229), .CI(n_238), .CO(n_241), .S(n_240));
   FA_X1 i_4023 (.A(n_369), .B(n_368), .CI(n_367), .CO(n_243), .S(n_242));
   FA_X1 i_4024 (.A(n_366), .B(n_365), .CI(n_364), .CO(n_245), .S(n_244));
   FA_X1 i_4025 (.A(n_363), .B(n_233), .CI(n_242), .CO(n_247), .S(n_246));
   FA_X1 i_4026 (.A(n_235), .B(n_244), .CI(n_246), .CO(n_249), .S(n_248));
   FA_X1 i_4027 (.A(n_237), .B(n_239), .CI(n_248), .CO(n_251), .S(n_250));
   FA_X1 i_4050 (.A(n_362), .B(n_361), .CI(n_243), .CO(n_253), .S(n_252));
   FA_X1 i_4051 (.A(n_360), .B(n_359), .CI(n_358), .CO(n_255), .S(n_254));
   FA_X1 i_4052 (.A(n_252), .B(n_245), .CI(n_247), .CO(n_257), .S(n_256));
   FA_X1 i_4053 (.A(n_254), .B(n_256), .CI(n_249), .CO(n_259), .S(n_258));
   FA_X1 i_4076 (.A(n_357), .B(n_356), .CI(n_355), .CO(n_261), .S(n_260));
   FA_X1 i_4077 (.A(n_253), .B(n_354), .CI(n_255), .CO(n_263), .S(n_262));
   FA_X1 i_4078 (.A(n_260), .B(n_257), .CI(n_262), .CO(n_265), .S(n_264));
   FA_X1 i_4093 (.A(n_353), .B(n_352), .CI(n_351), .CO(n_267), .S(n_266));
   FA_X1 i_4094 (.A(n_350), .B(n_349), .CI(n_266), .CO(n_269), .S(n_268));
   FA_X1 i_4095 (.A(n_261), .B(n_263), .CI(n_268), .CO(n_271), .S(n_270));
   FA_X1 i_4111 (.A(n_348), .B(n_347), .CI(n_346), .CO(n_273), .S(n_272));
   FA_X1 i_4112 (.A(n_267), .B(n_269), .CI(n_272), .CO(n_275), .S(n_274));
   FA_X1 i_4128 (.A(n_345), .B(n_344), .CI(n_273), .CO(n_277), .S(n_276));
   FA_X1 i_4136 (.A(n_343), .B(n_342), .CI(n_341), .CO(n_279), .S(n_278));
   FA_X1 i_4157 (.A(n_1034), .B(n_1029), .CI(n_340), .CO(n_280), .S(p_0[3]));
   FA_X1 i_4158 (.A(n_1039), .B(n_1052), .CI(n_280), .CO(n_281), .S(p_0[4]));
   FA_X1 i_4159 (.A(n_1070), .B(n_1068), .CI(n_281), .CO(n_282), .S(p_0[5]));
   FA_X1 i_4160 (.A(n_1096), .B(n_1094), .CI(n_282), .CO(n_283), .S(p_0[6]));
   FA_X1 i_4161 (.A(n_1122), .B(n_1124), .CI(n_283), .CO(n_284), .S(p_0[7]));
   FA_X1 i_4162 (.A(n_1151), .B(n_1153), .CI(n_284), .CO(n_285), .S(p_0[8]));
   FA_X1 i_4163 (.A(n_1190), .B(n_1188), .CI(n_285), .CO(n_286), .S(p_0[9]));
   FA_X1 i_4164 (.A(n_1229), .B(n_1227), .CI(n_286), .CO(n_287), .S(p_0[10]));
   FA_X1 i_4165 (.A(n_1267), .B(n_1269), .CI(n_287), .CO(n_288), .S(p_0[11]));
   FA_X1 i_4166 (.A(n_1315), .B(n_1317), .CI(n_288), .CO(n_289), .S(p_0[12]));
   FA_X1 i_4167 (.A(n_1365), .B(n_1367), .CI(n_289), .CO(n_290), .S(p_0[13]));
   FA_X1 i_4168 (.A(n_1416), .B(n_1418), .CI(n_290), .CO(n_291), .S(p_0[14]));
   FA_X1 i_4169 (.A(n_1475), .B(n_1477), .CI(n_291), .CO(n_292), .S(p_0[15]));
   FA_X1 i_4170 (.A(n_1536), .B(n_1538), .CI(n_292), .CO(n_293), .S(p_0[16]));
   FA_X1 i_4171 (.A(n_1598), .B(n_1600), .CI(n_293), .CO(n_294), .S(p_0[17]));
   FA_X1 i_4172 (.A(n_1601), .B(n_1670), .CI(n_294), .CO(n_295), .S(p_0[18]));
   FA_X1 i_4173 (.A(n_1671), .B(n_1742), .CI(n_295), .CO(n_296), .S(p_0[19]));
   FA_X1 i_4174 (.A(n_1813), .B(n_1815), .CI(n_296), .CO(n_297), .S(p_0[20]));
   FA_X1 i_4175 (.A(n_1816), .B(n_1896), .CI(n_297), .CO(n_298), .S(p_0[21]));
   FA_X1 i_4176 (.A(n_1897), .B(n_1979), .CI(n_298), .CO(n_299), .S(p_0[22]));
   FA_X1 i_4177 (.A(n_1980), .B(n_2063), .CI(n_299), .CO(n_300), .S(p_0[23]));
   FA_X1 i_4178 (.A(n_2064), .B(n_2155), .CI(n_300), .CO(n_301), .S(p_0[24]));
   FA_X1 i_4179 (.A(n_2247), .B(n_2249), .CI(n_301), .CO(n_302), .S(p_0[25]));
   FA_X1 i_4180 (.A(n_2250), .B(n_2344), .CI(n_302), .CO(n_303), .S(p_0[26]));
   FA_X1 i_4181 (.A(n_2345), .B(n_2447), .CI(n_303), .CO(n_304), .S(p_0[27]));
   FA_X1 i_4182 (.A(n_2448), .B(n_2552), .CI(n_304), .CO(n_305), .S(p_0[28]));
   FA_X1 i_4183 (.A(n_2553), .B(n_2658), .CI(n_305), .CO(n_306), .S(p_0[29]));
   FA_X1 i_4184 (.A(n_2659), .B(n_2772), .CI(n_306), .CO(n_307), .S(p_0[30]));
   FA_X1 i_4185 (.A(n_2773), .B(n_2888), .CI(n_307), .CO(n_308), .S(p_0[31]));
   FA_X1 i_4186 (.A(n_2889), .B(n_3004), .CI(n_308), .CO(n_309), .S(p_0[32]));
   FA_X1 i_4187 (.A(n_3005), .B(n_3112), .CI(n_309), .CO(n_310), .S(p_0[33]));
   FA_X1 i_4188 (.A(n_3113), .B(n_3219), .CI(n_310), .CO(n_311), .S(p_0[34]));
   FA_X1 i_4189 (.A(n_3220), .B(n_3324), .CI(n_311), .CO(n_312), .S(p_0[35]));
   FA_X1 i_4190 (.A(n_3421), .B(n_3325), .CI(n_312), .CO(n_313), .S(p_0[36]));
   FA_X1 i_4191 (.A(n_3422), .B(n_3517), .CI(n_313), .CO(n_314), .S(p_0[37]));
   FA_X1 i_4192 (.A(n_3518), .B(n_3611), .CI(n_314), .CO(n_315), .S(p_0[38]));
   FA_X1 i_4193 (.A(n_3612), .B(n_3697), .CI(n_315), .CO(n_316), .S(p_0[39]));
   FA_X1 i_4194 (.A(n_3698), .B(n_3782), .CI(n_316), .CO(n_317), .S(p_0[40]));
   FA_X1 i_4195 (.A(n_3783), .B(n_24), .CI(n_317), .CO(n_318), .S(p_0[41]));
   FA_X1 i_4196 (.A(n_25), .B(n_50), .CI(n_318), .CO(n_319), .S(p_0[42]));
   FA_X1 i_4197 (.A(n_51), .B(n_74), .CI(n_319), .CO(n_320), .S(p_0[43]));
   FA_X1 i_4198 (.A(n_75), .B(n_96), .CI(n_320), .CO(n_321), .S(p_0[44]));
   FA_X1 i_4199 (.A(n_97), .B(n_118), .CI(n_321), .CO(n_322), .S(p_0[45]));
   FA_X1 i_4200 (.A(n_119), .B(n_138), .CI(n_322), .CO(n_323), .S(p_0[46]));
   FA_X1 i_4201 (.A(n_139), .B(n_156), .CI(n_323), .CO(n_324), .S(p_0[47]));
   FA_X1 i_4202 (.A(n_157), .B(n_174), .CI(n_324), .CO(n_325), .S(p_0[48]));
   FA_X1 i_4203 (.A(n_190), .B(n_175), .CI(n_325), .CO(n_326), .S(p_0[49]));
   FA_X1 i_4204 (.A(n_191), .B(n_204), .CI(n_326), .CO(n_327), .S(p_0[50]));
   FA_X1 i_4205 (.A(n_205), .B(n_218), .CI(n_327), .CO(n_328), .S(p_0[51]));
   FA_X1 i_4206 (.A(n_230), .B(n_219), .CI(n_328), .CO(n_329), .S(p_0[52]));
   FA_X1 i_4207 (.A(n_231), .B(n_240), .CI(n_329), .CO(n_330), .S(p_0[53]));
   FA_X1 i_4208 (.A(n_241), .B(n_250), .CI(n_330), .CO(n_331), .S(p_0[54]));
   FA_X1 i_4209 (.A(n_258), .B(n_251), .CI(n_331), .CO(n_332), .S(p_0[55]));
   FA_X1 i_4210 (.A(n_259), .B(n_264), .CI(n_332), .CO(n_333), .S(p_0[56]));
   FA_X1 i_4211 (.A(n_270), .B(n_265), .CI(n_333), .CO(n_334), .S(p_0[57]));
   FA_X1 i_4212 (.A(n_271), .B(n_274), .CI(n_334), .CO(n_335), .S(p_0[58]));
   FA_X1 i_4213 (.A(n_276), .B(n_275), .CI(n_335), .CO(n_336), .S(p_0[59]));
   FA_X1 i_4214 (.A(n_277), .B(n_278), .CI(n_336), .CO(n_337), .S(p_0[60]));
   FA_X1 i_4215 (.A(n_339), .B(n_279), .CI(n_337), .CO(n_338), .S(p_0[61]));
   NAND2_X1 i_0 (.A1(a[30]), .A2(b[30]), .ZN(n_492));
   INV_X1 i_1 (.A(n_492), .ZN(n_493));
   NAND3_X1 i_2 (.A1(n_493), .A2(b[31]), .A3(a[29]), .ZN(n_494));
   INV_X1 i_3 (.A(n_494), .ZN(n_495));
   INV_X1 i_4 (.A(b[31]), .ZN(n_496));
   INV_X1 i_5 (.A(a[29]), .ZN(n_497));
   OAI21_X1 i_6 (.A(n_492), .B1(n_496), .B2(n_497), .ZN(n_498));
   INV_X1 i_7 (.A(a[31]), .ZN(n_499));
   INV_X1 i_8 (.A(b[29]), .ZN(n_500));
   NOR2_X1 i_9 (.A1(n_499), .A2(n_500), .ZN(n_501));
   AOI21_X1 i_10 (.A(n_495), .B1(n_498), .B2(n_501), .ZN(n_502));
   NAND2_X1 i_11 (.A1(a[31]), .A2(b[31]), .ZN(n_503));
   NOR2_X1 i_12 (.A1(n_492), .A2(n_503), .ZN(n_504));
   AOI22_X1 i_13 (.A1(a[31]), .A2(b[30]), .B1(b[31]), .B2(a[30]), .ZN(n_505));
   NOR2_X1 i_14 (.A1(n_504), .A2(n_505), .ZN(n_506));
   XNOR2_X1 i_15 (.A(n_502), .B(n_506), .ZN(n_339));
   NAND2_X1 i_16 (.A1(b[2]), .A2(a[1]), .ZN(n_507));
   NAND2_X1 i_17 (.A1(b[3]), .A2(a[2]), .ZN(n_508));
   NOR2_X1 i_18 (.A1(n_507), .A2(n_508), .ZN(n_509));
   AOI22_X1 i_19 (.A1(b[2]), .A2(a[2]), .B1(b[3]), .B2(a[1]), .ZN(n_510));
   NOR2_X1 i_20 (.A1(n_509), .A2(n_510), .ZN(n_511));
   NAND2_X1 i_21 (.A1(b[4]), .A2(a[0]), .ZN(n_512));
   XNOR2_X1 i_22 (.A(n_511), .B(n_512), .ZN(n_1039));
   INV_X1 i_23 (.A(a[0]), .ZN(n_513));
   INV_X1 i_24 (.A(b[0]), .ZN(n_514));
   NOR2_X1 i_25 (.A1(n_513), .A2(n_514), .ZN(p_0[0]));
   INV_X1 i_26 (.A(n_507), .ZN(n_515));
   NAND3_X1 i_27 (.A1(n_515), .A2(b[1]), .A3(a[0]), .ZN(n_516));
   INV_X1 i_28 (.A(n_516), .ZN(n_517));
   AOI22_X1 i_29 (.A1(b[1]), .A2(a[1]), .B1(b[2]), .B2(a[0]), .ZN(n_518));
   NOR2_X1 i_30 (.A1(n_517), .A2(n_518), .ZN(n_519));
   AOI21_X1 i_31 (.A(n_519), .B1(a[2]), .B2(b[0]), .ZN(n_520));
   NAND3_X1 i_32 (.A1(p_0[0]), .A2(b[1]), .A3(a[1]), .ZN(n_521));
   NAND3_X1 i_33 (.A1(n_519), .A2(a[2]), .A3(b[0]), .ZN(n_522));
   AOI21_X1 i_34 (.A(n_520), .B1(n_521), .B2(n_522), .ZN(n_340));
   NAND3_X1 i_35 (.A1(n_515), .A2(a[2]), .A3(b[1]), .ZN(n_523));
   AOI21_X1 i_36 (.A(n_515), .B1(a[2]), .B2(b[1]), .ZN(n_524));
   INV_X1 i_37 (.A(n_524), .ZN(n_525));
   NAND2_X1 i_38 (.A1(n_523), .A2(n_525), .ZN(n_526));
   NAND2_X1 i_39 (.A1(b[3]), .A2(a[0]), .ZN(n_527));
   XOR2_X1 i_40 (.A(n_526), .B(n_527), .Z(n_1029));
   NAND2_X1 i_41 (.A1(a[3]), .A2(b[0]), .ZN(n_528));
   XOR2_X1 i_42 (.A(n_516), .B(n_528), .Z(n_1034));
   AOI22_X1 i_43 (.A1(a[31]), .A2(b[27]), .B1(a[30]), .B2(b[28]), .ZN(n_529));
   NAND2_X1 i_44 (.A1(a[30]), .A2(b[27]), .ZN(n_530));
   INV_X1 i_45 (.A(b[26]), .ZN(n_531));
   OR3_X1 i_46 (.A1(n_530), .A2(n_499), .A3(n_531), .ZN(n_532));
   INV_X1 i_47 (.A(n_532), .ZN(n_533));
   AND2_X1 i_48 (.A1(a[29]), .A2(b[28]), .ZN(n_534));
   OAI21_X1 i_49 (.A(n_530), .B1(n_499), .B2(n_531), .ZN(n_535));
   AOI21_X1 i_50 (.A(n_533), .B1(n_534), .B2(n_535), .ZN(n_536));
   NAND2_X1 i_51 (.A1(a[31]), .A2(b[28]), .ZN(n_537));
   NOR2_X1 i_52 (.A1(n_530), .A2(n_537), .ZN(n_538));
   INV_X1 i_53 (.A(n_538), .ZN(n_539));
   AOI21_X1 i_54 (.A(n_529), .B1(n_536), .B2(n_539), .ZN(n_540));
   INV_X1 i_55 (.A(a[28]), .ZN(n_541));
   NOR2_X1 i_56 (.A1(n_500), .A2(n_541), .ZN(n_542));
   NAND3_X1 i_57 (.A1(n_542), .A2(a[29]), .A3(b[30]), .ZN(n_543));
   AOI22_X1 i_58 (.A1(b[30]), .A2(a[28]), .B1(a[29]), .B2(b[29]), .ZN(n_544));
   NAND2_X1 i_59 (.A1(b[31]), .A2(a[27]), .ZN(n_545));
   OAI21_X1 i_60 (.A(n_543), .B1(n_544), .B2(n_545), .ZN(n_546));
   NOR2_X1 i_61 (.A1(n_540), .A2(n_546), .ZN(n_547));
   NAND2_X1 i_62 (.A1(n_540), .A2(n_546), .ZN(n_548));
   AOI21_X1 i_63 (.A(n_547), .B1(n_537), .B2(n_548), .ZN(n_341));
   NAND2_X1 i_64 (.A1(n_494), .A2(n_498), .ZN(n_549));
   XNOR2_X1 i_65 (.A(n_549), .B(n_501), .ZN(n_342));
   NAND3_X1 i_66 (.A1(n_493), .A2(a[29]), .A3(b[29]), .ZN(n_550));
   AOI22_X1 i_67 (.A1(a[29]), .A2(b[30]), .B1(a[30]), .B2(b[29]), .ZN(n_551));
   NAND2_X1 i_68 (.A1(b[31]), .A2(a[28]), .ZN(n_552));
   OAI21_X1 i_69 (.A(n_550), .B1(n_551), .B2(n_552), .ZN(n_343));
   INV_X1 i_70 (.A(n_547), .ZN(n_553));
   NAND2_X1 i_71 (.A1(n_553), .A2(n_548), .ZN(n_554));
   XOR2_X1 i_72 (.A(n_554), .B(n_537), .Z(n_344));
   INV_X1 i_73 (.A(n_551), .ZN(n_555));
   NAND2_X1 i_74 (.A1(n_550), .A2(n_555), .ZN(n_556));
   XOR2_X1 i_75 (.A(n_556), .B(n_552), .Z(n_345));
   INV_X1 i_76 (.A(n_544), .ZN(n_557));
   NAND2_X1 i_77 (.A1(n_543), .A2(n_557), .ZN(n_558));
   XOR2_X1 i_78 (.A(n_558), .B(n_545), .Z(n_346));
   NOR2_X1 i_79 (.A1(n_538), .A2(n_529), .ZN(n_559));
   XNOR2_X1 i_80 (.A(n_536), .B(n_559), .ZN(n_347));
   NAND3_X1 i_81 (.A1(n_542), .A2(b[30]), .A3(a[27]), .ZN(n_560));
   AOI21_X1 i_82 (.A(n_542), .B1(b[30]), .B2(a[27]), .ZN(n_561));
   NAND2_X1 i_83 (.A1(b[31]), .A2(a[26]), .ZN(n_562));
   OAI21_X1 i_84 (.A(n_560), .B1(n_561), .B2(n_562), .ZN(n_348));
   INV_X1 i_85 (.A(n_561), .ZN(n_563));
   NAND2_X1 i_86 (.A1(n_560), .A2(n_563), .ZN(n_564));
   XOR2_X1 i_87 (.A(n_564), .B(n_562), .Z(n_349));
   NAND2_X1 i_88 (.A1(n_532), .A2(n_535), .ZN(n_565));
   XNOR2_X1 i_89 (.A(n_565), .B(n_534), .ZN(n_350));
   NAND2_X1 i_90 (.A1(a[29]), .A2(b[26]), .ZN(n_566));
   INV_X1 i_91 (.A(n_566), .ZN(n_567));
   NAND3_X1 i_92 (.A1(n_567), .A2(a[28]), .A3(b[27]), .ZN(n_568));
   AOI21_X1 i_93 (.A(n_567), .B1(a[28]), .B2(b[27]), .ZN(n_569));
   NAND2_X1 i_94 (.A1(b[28]), .A2(a[27]), .ZN(n_570));
   OAI21_X1 i_95 (.A(n_568), .B1(n_569), .B2(n_570), .ZN(n_571));
   NAND4_X1 i_96 (.A1(b[30]), .A2(b[29]), .A3(a[26]), .A4(a[25]), .ZN(n_572));
   AOI22_X1 i_97 (.A1(b[30]), .A2(a[25]), .B1(b[29]), .B2(a[26]), .ZN(n_573));
   NAND2_X1 i_98 (.A1(b[31]), .A2(a[24]), .ZN(n_574));
   OAI21_X1 i_99 (.A(n_572), .B1(n_573), .B2(n_574), .ZN(n_575));
   NOR2_X1 i_100 (.A1(n_571), .A2(n_575), .ZN(n_576));
   NAND2_X1 i_101 (.A1(a[31]), .A2(b[25]), .ZN(n_577));
   NAND2_X1 i_102 (.A1(n_571), .A2(n_575), .ZN(n_578));
   AOI21_X1 i_103 (.A(n_576), .B1(n_577), .B2(n_578), .ZN(n_351));
   NAND4_X1 i_104 (.A1(b[30]), .A2(b[29]), .A3(a[26]), .A4(a[27]), .ZN(n_579));
   AOI22_X1 i_105 (.A1(b[30]), .A2(a[26]), .B1(b[29]), .B2(a[27]), .ZN(n_580));
   NAND2_X1 i_106 (.A1(b[31]), .A2(a[25]), .ZN(n_581));
   OAI21_X1 i_107 (.A(n_579), .B1(n_580), .B2(n_581), .ZN(n_352));
   NOR2_X1 i_108 (.A1(n_530), .A2(n_566), .ZN(n_582));
   INV_X1 i_109 (.A(n_582), .ZN(n_583));
   AOI22_X1 i_110 (.A1(a[29]), .A2(b[27]), .B1(a[30]), .B2(b[26]), .ZN(n_584));
   NAND2_X1 i_111 (.A1(a[28]), .A2(b[28]), .ZN(n_585));
   OAI21_X1 i_112 (.A(n_583), .B1(n_584), .B2(n_585), .ZN(n_353));
   INV_X1 i_113 (.A(n_576), .ZN(n_586));
   NAND2_X1 i_114 (.A1(n_578), .A2(n_586), .ZN(n_587));
   XOR2_X1 i_115 (.A(n_587), .B(n_577), .Z(n_354));
   INV_X1 i_116 (.A(n_580), .ZN(n_588));
   NAND2_X1 i_117 (.A1(n_588), .A2(n_579), .ZN(n_589));
   XOR2_X1 i_118 (.A(n_589), .B(n_581), .Z(n_355));
   NOR2_X1 i_119 (.A1(n_582), .A2(n_584), .ZN(n_590));
   XNOR2_X1 i_120 (.A(n_590), .B(n_585), .ZN(n_356));
   INV_X1 i_121 (.A(b[25]), .ZN(n_591));
   NAND2_X1 i_122 (.A1(a[30]), .A2(b[24]), .ZN(n_592));
   NAND2_X1 i_123 (.A1(a[31]), .A2(b[23]), .ZN(n_593));
   AOI211_X1 i_124 (.A(n_497), .B(n_591), .C1(n_592), .C2(n_593), .ZN(n_594));
   AOI21_X1 i_125 (.A(n_594), .B1(a[31]), .B2(b[24]), .ZN(n_595));
   AND2_X1 i_126 (.A1(a[30]), .A2(b[23]), .ZN(n_596));
   OAI211_X1 i_127 (.A(a[31]), .B(b[24]), .C1(n_594), .C2(n_596), .ZN(n_597));
   NAND2_X1 i_128 (.A1(a[30]), .A2(b[25]), .ZN(n_598));
   AOI21_X1 i_129 (.A(n_595), .B1(n_597), .B2(n_598), .ZN(n_357));
   INV_X1 i_130 (.A(n_573), .ZN(n_599));
   NAND2_X1 i_131 (.A1(n_599), .A2(n_572), .ZN(n_600));
   XOR2_X1 i_132 (.A(n_600), .B(n_574), .Z(n_358));
   INV_X1 i_133 (.A(n_569), .ZN(n_601));
   NAND2_X1 i_134 (.A1(n_568), .A2(n_601), .ZN(n_602));
   XOR2_X1 i_135 (.A(n_602), .B(n_570), .Z(n_359));
   INV_X1 i_136 (.A(n_595), .ZN(n_603));
   NAND2_X1 i_137 (.A1(n_597), .A2(n_603), .ZN(n_604));
   XOR2_X1 i_138 (.A(n_604), .B(n_598), .Z(n_360));
   NAND4_X1 i_139 (.A1(b[30]), .A2(b[29]), .A3(a[25]), .A4(a[24]), .ZN(n_605));
   AOI22_X1 i_140 (.A1(b[30]), .A2(a[24]), .B1(b[29]), .B2(a[25]), .ZN(n_606));
   NAND2_X1 i_141 (.A1(b[31]), .A2(a[23]), .ZN(n_607));
   OAI21_X1 i_142 (.A(n_605), .B1(n_606), .B2(n_607), .ZN(n_361));
   NAND4_X1 i_143 (.A1(a[28]), .A2(a[27]), .A3(b[27]), .A4(b[26]), .ZN(n_608));
   AOI22_X1 i_144 (.A1(a[27]), .A2(b[27]), .B1(a[28]), .B2(b[26]), .ZN(n_609));
   NAND2_X1 i_145 (.A1(b[28]), .A2(a[26]), .ZN(n_610));
   OAI21_X1 i_146 (.A(n_608), .B1(n_609), .B2(n_610), .ZN(n_362));
   INV_X1 i_147 (.A(n_606), .ZN(n_611));
   NAND2_X1 i_148 (.A1(n_611), .A2(n_605), .ZN(n_612));
   XOR2_X1 i_149 (.A(n_612), .B(n_607), .Z(n_363));
   INV_X1 i_150 (.A(n_609), .ZN(n_613));
   NAND2_X1 i_151 (.A1(n_613), .A2(n_608), .ZN(n_614));
   XOR2_X1 i_152 (.A(n_614), .B(n_610), .Z(n_364));
   XOR2_X1 i_153 (.A(n_592), .B(n_593), .Z(n_615));
   NAND2_X1 i_154 (.A1(a[29]), .A2(b[25]), .ZN(n_616));
   XNOR2_X1 i_155 (.A(n_615), .B(n_616), .ZN(n_365));
   NAND4_X1 i_156 (.A1(a[26]), .A2(b[27]), .A3(b[26]), .A4(a[25]), .ZN(n_617));
   AOI22_X1 i_157 (.A1(b[27]), .A2(a[25]), .B1(a[26]), .B2(b[26]), .ZN(n_618));
   NAND2_X1 i_158 (.A1(b[28]), .A2(a[24]), .ZN(n_619));
   OAI21_X1 i_159 (.A(n_617), .B1(n_618), .B2(n_619), .ZN(n_620));
   NAND4_X1 i_160 (.A1(a[29]), .A2(a[28]), .A3(b[24]), .A4(b[23]), .ZN(n_621));
   AOI22_X1 i_161 (.A1(a[28]), .A2(b[24]), .B1(a[29]), .B2(b[23]), .ZN(n_622));
   NAND2_X1 i_162 (.A1(a[27]), .A2(b[25]), .ZN(n_623));
   OAI21_X1 i_163 (.A(n_621), .B1(n_622), .B2(n_623), .ZN(n_624));
   NOR2_X1 i_164 (.A1(n_620), .A2(n_624), .ZN(n_625));
   NAND2_X1 i_165 (.A1(a[31]), .A2(b[22]), .ZN(n_626));
   NAND2_X1 i_166 (.A1(n_620), .A2(n_624), .ZN(n_627));
   AOI21_X1 i_167 (.A(n_625), .B1(n_626), .B2(n_627), .ZN(n_366));
   NAND4_X1 i_168 (.A1(b[30]), .A2(b[29]), .A3(a[23]), .A4(a[24]), .ZN(n_628));
   AOI22_X1 i_169 (.A1(b[30]), .A2(a[23]), .B1(b[29]), .B2(a[24]), .ZN(n_629));
   NAND2_X1 i_170 (.A1(b[31]), .A2(a[22]), .ZN(n_630));
   OAI21_X1 i_171 (.A(n_628), .B1(n_629), .B2(n_630), .ZN(n_367));
   NAND4_X1 i_172 (.A1(a[26]), .A2(a[27]), .A3(b[27]), .A4(b[26]), .ZN(n_631));
   AOI22_X1 i_173 (.A1(a[26]), .A2(b[27]), .B1(a[27]), .B2(b[26]), .ZN(n_632));
   NAND2_X1 i_174 (.A1(b[28]), .A2(a[25]), .ZN(n_633));
   OAI21_X1 i_175 (.A(n_631), .B1(n_632), .B2(n_633), .ZN(n_368));
   INV_X1 i_176 (.A(n_592), .ZN(n_634));
   NAND3_X1 i_177 (.A1(n_634), .A2(a[29]), .A3(b[23]), .ZN(n_635));
   AOI21_X1 i_178 (.A(n_596), .B1(a[29]), .B2(b[24]), .ZN(n_636));
   NAND2_X1 i_179 (.A1(a[28]), .A2(b[25]), .ZN(n_637));
   OAI21_X1 i_180 (.A(n_635), .B1(n_636), .B2(n_637), .ZN(n_369));
   INV_X1 i_181 (.A(n_625), .ZN(n_638));
   NAND2_X1 i_182 (.A1(n_638), .A2(n_627), .ZN(n_639));
   XOR2_X1 i_183 (.A(n_639), .B(n_626), .Z(n_370));
   INV_X1 i_184 (.A(n_629), .ZN(n_640));
   NAND2_X1 i_185 (.A1(n_640), .A2(n_628), .ZN(n_641));
   XOR2_X1 i_186 (.A(n_641), .B(n_630), .Z(n_371));
   INV_X1 i_187 (.A(n_632), .ZN(n_642));
   NAND2_X1 i_188 (.A1(n_642), .A2(n_631), .ZN(n_643));
   XOR2_X1 i_189 (.A(n_643), .B(n_633), .Z(n_372));
   INV_X1 i_190 (.A(n_636), .ZN(n_644));
   NAND2_X1 i_191 (.A1(n_635), .A2(n_644), .ZN(n_645));
   XOR2_X1 i_192 (.A(n_645), .B(n_637), .Z(n_373));
   NAND4_X1 i_193 (.A1(b[30]), .A2(b[29]), .A3(a[23]), .A4(a[22]), .ZN(n_646));
   AOI22_X1 i_194 (.A1(b[30]), .A2(a[22]), .B1(b[29]), .B2(a[23]), .ZN(n_647));
   NAND2_X1 i_195 (.A1(b[31]), .A2(a[21]), .ZN(n_648));
   OAI21_X1 i_196 (.A(n_646), .B1(n_647), .B2(n_648), .ZN(n_374));
   INV_X1 i_197 (.A(n_647), .ZN(n_649));
   NAND2_X1 i_198 (.A1(n_649), .A2(n_646), .ZN(n_650));
   XOR2_X1 i_199 (.A(n_650), .B(n_648), .Z(n_375));
   INV_X1 i_200 (.A(n_618), .ZN(n_651));
   NAND2_X1 i_201 (.A1(n_651), .A2(n_617), .ZN(n_652));
   XOR2_X1 i_202 (.A(n_652), .B(n_619), .Z(n_376));
   INV_X1 i_203 (.A(n_622), .ZN(n_653));
   NAND2_X1 i_204 (.A1(n_653), .A2(n_621), .ZN(n_654));
   XOR2_X1 i_205 (.A(n_654), .B(n_623), .Z(n_377));
   INV_X1 i_206 (.A(b[22]), .ZN(n_655));
   NAND2_X1 i_207 (.A1(a[30]), .A2(b[21]), .ZN(n_656));
   NAND2_X1 i_208 (.A1(a[31]), .A2(b[20]), .ZN(n_657));
   AOI211_X1 i_209 (.A(n_497), .B(n_655), .C1(n_656), .C2(n_657), .ZN(n_658));
   INV_X1 i_210 (.A(a[30]), .ZN(n_659));
   INV_X1 i_211 (.A(b[20]), .ZN(n_660));
   NOR2_X1 i_212 (.A1(n_659), .A2(n_660), .ZN(n_661));
   OAI211_X1 i_213 (.A(a[31]), .B(b[21]), .C1(n_658), .C2(n_661), .ZN(n_662));
   AOI21_X1 i_214 (.A(n_658), .B1(a[31]), .B2(b[21]), .ZN(n_663));
   NAND2_X1 i_215 (.A1(a[30]), .A2(b[22]), .ZN(n_664));
   OAI21_X1 i_216 (.A(n_662), .B1(n_663), .B2(n_664), .ZN(n_378));
   AND2_X1 i_217 (.A1(n_663), .A2(n_664), .ZN(n_665));
   OAI22_X1 i_218 (.A1(n_662), .A2(n_664), .B1(n_378), .B2(n_665), .ZN(n_379));
   NAND4_X1 i_219 (.A1(b[30]), .A2(b[29]), .A3(a[22]), .A4(a[21]), .ZN(n_666));
   AOI22_X1 i_220 (.A1(b[30]), .A2(a[21]), .B1(b[29]), .B2(a[22]), .ZN(n_667));
   NAND2_X1 i_221 (.A1(b[31]), .A2(a[20]), .ZN(n_668));
   OAI21_X1 i_222 (.A(n_666), .B1(n_667), .B2(n_668), .ZN(n_380));
   NAND4_X1 i_223 (.A1(b[27]), .A2(b[26]), .A3(a[25]), .A4(a[24]), .ZN(n_669));
   AOI22_X1 i_224 (.A1(b[27]), .A2(a[24]), .B1(b[26]), .B2(a[25]), .ZN(n_670));
   NAND2_X1 i_225 (.A1(b[28]), .A2(a[23]), .ZN(n_671));
   OAI21_X1 i_226 (.A(n_669), .B1(n_670), .B2(n_671), .ZN(n_381));
   NAND4_X1 i_227 (.A1(a[28]), .A2(a[27]), .A3(b[24]), .A4(b[23]), .ZN(n_672));
   AOI22_X1 i_228 (.A1(a[27]), .A2(b[24]), .B1(a[28]), .B2(b[23]), .ZN(n_673));
   NAND2_X1 i_229 (.A1(a[26]), .A2(b[25]), .ZN(n_674));
   OAI21_X1 i_230 (.A(n_672), .B1(n_673), .B2(n_674), .ZN(n_382));
   INV_X1 i_231 (.A(n_667), .ZN(n_675));
   NAND2_X1 i_232 (.A1(n_675), .A2(n_666), .ZN(n_676));
   XOR2_X1 i_233 (.A(n_676), .B(n_668), .Z(n_383));
   INV_X1 i_234 (.A(n_670), .ZN(n_677));
   NAND2_X1 i_235 (.A1(n_677), .A2(n_669), .ZN(n_678));
   XOR2_X1 i_236 (.A(n_678), .B(n_671), .Z(n_384));
   INV_X1 i_237 (.A(n_673), .ZN(n_679));
   NAND2_X1 i_238 (.A1(n_679), .A2(n_672), .ZN(n_680));
   XOR2_X1 i_239 (.A(n_680), .B(n_674), .Z(n_385));
   XOR2_X1 i_240 (.A(n_656), .B(n_657), .Z(n_681));
   NAND2_X1 i_241 (.A1(a[29]), .A2(b[22]), .ZN(n_682));
   XNOR2_X1 i_242 (.A(n_681), .B(n_682), .ZN(n_386));
   NOR2_X1 i_243 (.A1(n_497), .A2(n_660), .ZN(n_683));
   NAND3_X1 i_244 (.A1(n_683), .A2(a[28]), .A3(b[21]), .ZN(n_684));
   AOI21_X1 i_245 (.A(n_683), .B1(a[28]), .B2(b[21]), .ZN(n_685));
   NAND2_X1 i_246 (.A1(a[27]), .A2(b[22]), .ZN(n_686));
   OAI21_X1 i_247 (.A(n_684), .B1(n_685), .B2(n_686), .ZN(n_687));
   NAND4_X1 i_248 (.A1(a[26]), .A2(a[25]), .A3(b[24]), .A4(b[23]), .ZN(n_688));
   AOI22_X1 i_249 (.A1(a[25]), .A2(b[24]), .B1(a[26]), .B2(b[23]), .ZN(n_689));
   NAND2_X1 i_250 (.A1(b[25]), .A2(a[24]), .ZN(n_690));
   OAI21_X1 i_251 (.A(n_688), .B1(n_689), .B2(n_690), .ZN(n_691));
   NOR2_X1 i_252 (.A1(n_687), .A2(n_691), .ZN(n_692));
   NAND2_X1 i_253 (.A1(a[31]), .A2(b[19]), .ZN(n_693));
   NAND2_X1 i_254 (.A1(n_687), .A2(n_691), .ZN(n_694));
   AOI21_X1 i_255 (.A(n_692), .B1(n_693), .B2(n_694), .ZN(n_387));
   NAND4_X1 i_256 (.A1(b[30]), .A2(b[29]), .A3(a[20]), .A4(a[21]), .ZN(n_695));
   AOI22_X1 i_257 (.A1(b[30]), .A2(a[20]), .B1(b[29]), .B2(a[21]), .ZN(n_696));
   NAND2_X1 i_258 (.A1(b[31]), .A2(a[19]), .ZN(n_697));
   OAI21_X1 i_259 (.A(n_695), .B1(n_696), .B2(n_697), .ZN(n_388));
   NAND4_X1 i_260 (.A1(b[27]), .A2(b[26]), .A3(a[23]), .A4(a[24]), .ZN(n_698));
   AOI22_X1 i_261 (.A1(b[27]), .A2(a[23]), .B1(b[26]), .B2(a[24]), .ZN(n_699));
   NAND2_X1 i_262 (.A1(b[28]), .A2(a[22]), .ZN(n_700));
   OAI21_X1 i_263 (.A(n_698), .B1(n_699), .B2(n_700), .ZN(n_389));
   NAND4_X1 i_264 (.A1(a[26]), .A2(a[27]), .A3(b[24]), .A4(b[23]), .ZN(n_701));
   AOI22_X1 i_265 (.A1(a[26]), .A2(b[24]), .B1(a[27]), .B2(b[23]), .ZN(n_702));
   NAND2_X1 i_266 (.A1(a[25]), .A2(b[25]), .ZN(n_703));
   OAI21_X1 i_267 (.A(n_701), .B1(n_702), .B2(n_703), .ZN(n_390));
   INV_X1 i_268 (.A(n_656), .ZN(n_704));
   NAND2_X1 i_269 (.A1(n_704), .A2(n_683), .ZN(n_705));
   AOI21_X1 i_270 (.A(n_661), .B1(a[29]), .B2(b[21]), .ZN(n_706));
   NAND2_X1 i_271 (.A1(a[28]), .A2(b[22]), .ZN(n_707));
   OAI21_X1 i_272 (.A(n_705), .B1(n_706), .B2(n_707), .ZN(n_391));
   INV_X1 i_273 (.A(n_692), .ZN(n_708));
   NAND2_X1 i_274 (.A1(n_694), .A2(n_708), .ZN(n_709));
   XOR2_X1 i_275 (.A(n_709), .B(n_693), .Z(n_392));
   INV_X1 i_276 (.A(n_696), .ZN(n_710));
   NAND2_X1 i_277 (.A1(n_710), .A2(n_695), .ZN(n_711));
   XOR2_X1 i_278 (.A(n_711), .B(n_697), .Z(n_393));
   INV_X1 i_279 (.A(n_699), .ZN(n_712));
   NAND2_X1 i_280 (.A1(n_712), .A2(n_698), .ZN(n_713));
   XOR2_X1 i_281 (.A(n_713), .B(n_700), .Z(n_394));
   INV_X1 i_282 (.A(n_702), .ZN(n_714));
   NAND2_X1 i_283 (.A1(n_714), .A2(n_701), .ZN(n_715));
   XOR2_X1 i_284 (.A(n_715), .B(n_703), .Z(n_395));
   INV_X1 i_285 (.A(n_706), .ZN(n_716));
   NAND2_X1 i_286 (.A1(n_705), .A2(n_716), .ZN(n_717));
   XOR2_X1 i_287 (.A(n_717), .B(n_707), .Z(n_396));
   NAND2_X1 i_288 (.A1(a[29]), .A2(b[19]), .ZN(n_718));
   NAND2_X1 i_289 (.A1(a[30]), .A2(b[18]), .ZN(n_719));
   NAND2_X1 i_290 (.A1(a[31]), .A2(b[17]), .ZN(n_720));
   AOI21_X1 i_291 (.A(n_718), .B1(n_719), .B2(n_720), .ZN(n_721));
   AND2_X1 i_292 (.A1(a[30]), .A2(b[17]), .ZN(n_722));
   OAI211_X1 i_293 (.A(a[31]), .B(b[18]), .C1(n_721), .C2(n_722), .ZN(n_723));
   AOI21_X1 i_294 (.A(n_721), .B1(a[31]), .B2(b[18]), .ZN(n_724));
   NAND2_X1 i_295 (.A1(a[30]), .A2(b[19]), .ZN(n_725));
   OAI21_X1 i_296 (.A(n_723), .B1(n_724), .B2(n_725), .ZN(n_397));
   NAND4_X1 i_297 (.A1(b[30]), .A2(b[29]), .A3(a[20]), .A4(a[19]), .ZN(n_726));
   AOI22_X1 i_298 (.A1(b[30]), .A2(a[19]), .B1(b[29]), .B2(a[20]), .ZN(n_727));
   NAND2_X1 i_299 (.A1(b[31]), .A2(a[18]), .ZN(n_728));
   OAI21_X1 i_300 (.A(n_726), .B1(n_727), .B2(n_728), .ZN(n_398));
   NAND4_X1 i_301 (.A1(b[27]), .A2(b[26]), .A3(a[23]), .A4(a[22]), .ZN(n_729));
   AOI22_X1 i_302 (.A1(b[27]), .A2(a[22]), .B1(b[26]), .B2(a[23]), .ZN(n_730));
   NAND2_X1 i_303 (.A1(b[28]), .A2(a[21]), .ZN(n_731));
   OAI21_X1 i_304 (.A(n_729), .B1(n_730), .B2(n_731), .ZN(n_399));
   INV_X1 i_305 (.A(n_727), .ZN(n_732));
   NAND2_X1 i_306 (.A1(n_732), .A2(n_726), .ZN(n_733));
   XOR2_X1 i_307 (.A(n_733), .B(n_728), .Z(n_400));
   INV_X1 i_308 (.A(n_730), .ZN(n_734));
   NAND2_X1 i_309 (.A1(n_734), .A2(n_729), .ZN(n_735));
   XOR2_X1 i_310 (.A(n_735), .B(n_731), .Z(n_401));
   INV_X1 i_311 (.A(n_689), .ZN(n_736));
   NAND2_X1 i_312 (.A1(n_736), .A2(n_688), .ZN(n_737));
   XOR2_X1 i_313 (.A(n_737), .B(n_690), .Z(n_402));
   INV_X1 i_314 (.A(n_685), .ZN(n_738));
   NAND2_X1 i_315 (.A1(n_684), .A2(n_738), .ZN(n_739));
   XOR2_X1 i_316 (.A(n_739), .B(n_686), .Z(n_403));
   INV_X1 i_317 (.A(n_724), .ZN(n_740));
   NAND2_X1 i_318 (.A1(n_723), .A2(n_740), .ZN(n_741));
   XOR2_X1 i_319 (.A(n_741), .B(n_725), .Z(n_404));
   NAND4_X1 i_320 (.A1(b[30]), .A2(b[29]), .A3(a[19]), .A4(a[18]), .ZN(n_742));
   AOI22_X1 i_321 (.A1(b[30]), .A2(a[18]), .B1(b[29]), .B2(a[19]), .ZN(n_743));
   NAND2_X1 i_322 (.A1(b[31]), .A2(a[17]), .ZN(n_744));
   OAI21_X1 i_323 (.A(n_742), .B1(n_743), .B2(n_744), .ZN(n_405));
   NAND4_X1 i_324 (.A1(b[27]), .A2(b[26]), .A3(a[22]), .A4(a[21]), .ZN(n_745));
   AOI22_X1 i_325 (.A1(b[27]), .A2(a[21]), .B1(b[26]), .B2(a[22]), .ZN(n_746));
   NAND2_X1 i_326 (.A1(b[28]), .A2(a[20]), .ZN(n_747));
   OAI21_X1 i_327 (.A(n_745), .B1(n_746), .B2(n_747), .ZN(n_406));
   NAND4_X1 i_328 (.A1(a[25]), .A2(a[24]), .A3(b[24]), .A4(b[23]), .ZN(n_748));
   AOI22_X1 i_329 (.A1(a[24]), .A2(b[24]), .B1(a[25]), .B2(b[23]), .ZN(n_749));
   NAND2_X1 i_330 (.A1(b[25]), .A2(a[23]), .ZN(n_750));
   OAI21_X1 i_331 (.A(n_748), .B1(n_749), .B2(n_750), .ZN(n_407));
   NAND4_X1 i_332 (.A1(a[28]), .A2(a[27]), .A3(b[21]), .A4(b[20]), .ZN(n_751));
   AOI22_X1 i_333 (.A1(a[27]), .A2(b[21]), .B1(a[28]), .B2(b[20]), .ZN(n_752));
   NAND2_X1 i_334 (.A1(a[26]), .A2(b[22]), .ZN(n_753));
   OAI21_X1 i_335 (.A(n_751), .B1(n_752), .B2(n_753), .ZN(n_408));
   INV_X1 i_336 (.A(n_743), .ZN(n_754));
   NAND2_X1 i_337 (.A1(n_754), .A2(n_742), .ZN(n_755));
   XOR2_X1 i_338 (.A(n_755), .B(n_744), .Z(n_409));
   INV_X1 i_339 (.A(n_746), .ZN(n_756));
   NAND2_X1 i_340 (.A1(n_756), .A2(n_745), .ZN(n_757));
   XOR2_X1 i_341 (.A(n_757), .B(n_747), .Z(n_410));
   INV_X1 i_342 (.A(n_749), .ZN(n_758));
   NAND2_X1 i_343 (.A1(n_758), .A2(n_748), .ZN(n_759));
   XOR2_X1 i_344 (.A(n_759), .B(n_750), .Z(n_411));
   INV_X1 i_345 (.A(n_752), .ZN(n_760));
   NAND2_X1 i_346 (.A1(n_760), .A2(n_751), .ZN(n_761));
   XOR2_X1 i_347 (.A(n_761), .B(n_753), .Z(n_412));
   XNOR2_X1 i_348 (.A(n_719), .B(n_720), .ZN(n_762));
   XOR2_X1 i_349 (.A(n_762), .B(n_718), .Z(n_413));
   NAND4_X1 i_350 (.A1(a[26]), .A2(a[25]), .A3(b[21]), .A4(b[20]), .ZN(n_763));
   AOI22_X1 i_351 (.A1(a[25]), .A2(b[21]), .B1(a[26]), .B2(b[20]), .ZN(n_764));
   NAND2_X1 i_352 (.A1(a[24]), .A2(b[22]), .ZN(n_765));
   OAI21_X1 i_353 (.A(n_763), .B1(n_764), .B2(n_765), .ZN(n_766));
   NAND4_X1 i_354 (.A1(a[29]), .A2(a[28]), .A3(b[18]), .A4(b[17]), .ZN(n_767));
   AOI22_X1 i_355 (.A1(a[28]), .A2(b[18]), .B1(a[29]), .B2(b[17]), .ZN(n_768));
   NAND2_X1 i_356 (.A1(a[27]), .A2(b[19]), .ZN(n_769));
   OAI21_X1 i_357 (.A(n_767), .B1(n_768), .B2(n_769), .ZN(n_770));
   NOR2_X1 i_358 (.A1(n_766), .A2(n_770), .ZN(n_771));
   NAND2_X1 i_359 (.A1(a[31]), .A2(b[16]), .ZN(n_772));
   NAND2_X1 i_360 (.A1(n_766), .A2(n_770), .ZN(n_773));
   AOI21_X1 i_361 (.A(n_771), .B1(n_772), .B2(n_773), .ZN(n_414));
   NAND4_X1 i_362 (.A1(b[30]), .A2(b[29]), .A3(a[17]), .A4(a[18]), .ZN(n_774));
   AOI22_X1 i_363 (.A1(b[30]), .A2(a[17]), .B1(b[29]), .B2(a[18]), .ZN(n_775));
   NAND2_X1 i_364 (.A1(b[31]), .A2(a[16]), .ZN(n_776));
   OAI21_X1 i_365 (.A(n_774), .B1(n_775), .B2(n_776), .ZN(n_415));
   NAND4_X1 i_366 (.A1(b[27]), .A2(b[26]), .A3(a[20]), .A4(a[21]), .ZN(n_777));
   AOI22_X1 i_367 (.A1(b[27]), .A2(a[20]), .B1(b[26]), .B2(a[21]), .ZN(n_778));
   NAND2_X1 i_368 (.A1(b[28]), .A2(a[19]), .ZN(n_779));
   OAI21_X1 i_369 (.A(n_777), .B1(n_778), .B2(n_779), .ZN(n_416));
   NAND4_X1 i_370 (.A1(a[23]), .A2(a[24]), .A3(b[24]), .A4(b[23]), .ZN(n_780));
   AOI22_X1 i_371 (.A1(a[23]), .A2(b[24]), .B1(a[24]), .B2(b[23]), .ZN(n_781));
   NAND2_X1 i_372 (.A1(b[25]), .A2(a[22]), .ZN(n_782));
   OAI21_X1 i_373 (.A(n_780), .B1(n_781), .B2(n_782), .ZN(n_417));
   NAND4_X1 i_374 (.A1(a[26]), .A2(a[27]), .A3(b[21]), .A4(b[20]), .ZN(n_783));
   AOI22_X1 i_375 (.A1(a[26]), .A2(b[21]), .B1(a[27]), .B2(b[20]), .ZN(n_784));
   NAND2_X1 i_376 (.A1(a[25]), .A2(b[22]), .ZN(n_785));
   OAI21_X1 i_377 (.A(n_783), .B1(n_784), .B2(n_785), .ZN(n_418));
   INV_X1 i_378 (.A(n_719), .ZN(n_786));
   NAND3_X1 i_379 (.A1(n_786), .A2(a[29]), .A3(b[17]), .ZN(n_787));
   AOI21_X1 i_380 (.A(n_722), .B1(a[29]), .B2(b[18]), .ZN(n_788));
   NAND2_X1 i_381 (.A1(a[28]), .A2(b[19]), .ZN(n_789));
   OAI21_X1 i_382 (.A(n_787), .B1(n_788), .B2(n_789), .ZN(n_419));
   INV_X1 i_383 (.A(n_771), .ZN(n_790));
   NAND2_X1 i_384 (.A1(n_790), .A2(n_773), .ZN(n_791));
   XOR2_X1 i_385 (.A(n_791), .B(n_772), .Z(n_420));
   INV_X1 i_386 (.A(n_775), .ZN(n_792));
   NAND2_X1 i_387 (.A1(n_792), .A2(n_774), .ZN(n_793));
   XOR2_X1 i_388 (.A(n_793), .B(n_776), .Z(n_421));
   INV_X1 i_389 (.A(n_778), .ZN(n_794));
   NAND2_X1 i_390 (.A1(n_794), .A2(n_777), .ZN(n_795));
   XOR2_X1 i_391 (.A(n_795), .B(n_779), .Z(n_422));
   INV_X1 i_392 (.A(n_781), .ZN(n_796));
   NAND2_X1 i_393 (.A1(n_796), .A2(n_780), .ZN(n_797));
   XOR2_X1 i_394 (.A(n_797), .B(n_782), .Z(n_423));
   INV_X1 i_395 (.A(n_784), .ZN(n_798));
   NAND2_X1 i_396 (.A1(n_798), .A2(n_783), .ZN(n_799));
   XOR2_X1 i_397 (.A(n_799), .B(n_785), .Z(n_424));
   INV_X1 i_398 (.A(n_788), .ZN(n_800));
   NAND2_X1 i_399 (.A1(n_787), .A2(n_800), .ZN(n_801));
   XOR2_X1 i_400 (.A(n_801), .B(n_789), .Z(n_425));
   INV_X1 i_401 (.A(b[16]), .ZN(n_802));
   NAND2_X1 i_402 (.A1(a[30]), .A2(b[15]), .ZN(n_803));
   NAND2_X1 i_403 (.A1(a[31]), .A2(b[14]), .ZN(n_804));
   AOI211_X1 i_404 (.A(n_497), .B(n_802), .C1(n_803), .C2(n_804), .ZN(n_805));
   AOI21_X1 i_405 (.A(n_805), .B1(a[31]), .B2(b[15]), .ZN(n_806));
   AND2_X1 i_406 (.A1(a[30]), .A2(b[14]), .ZN(n_807));
   OAI211_X1 i_407 (.A(a[31]), .B(b[15]), .C1(n_805), .C2(n_807), .ZN(n_808));
   NAND2_X1 i_408 (.A1(a[30]), .A2(b[16]), .ZN(n_809));
   AOI21_X1 i_409 (.A(n_806), .B1(n_808), .B2(n_809), .ZN(n_426));
   NAND4_X1 i_410 (.A1(b[30]), .A2(b[29]), .A3(a[17]), .A4(a[16]), .ZN(n_810));
   AOI22_X1 i_411 (.A1(b[30]), .A2(a[16]), .B1(b[29]), .B2(a[17]), .ZN(n_811));
   NAND2_X1 i_412 (.A1(b[31]), .A2(a[15]), .ZN(n_812));
   OAI21_X1 i_413 (.A(n_810), .B1(n_811), .B2(n_812), .ZN(n_427));
   NAND4_X1 i_414 (.A1(b[27]), .A2(b[26]), .A3(a[20]), .A4(a[19]), .ZN(n_813));
   AOI22_X1 i_415 (.A1(b[27]), .A2(a[19]), .B1(b[26]), .B2(a[20]), .ZN(n_814));
   NAND2_X1 i_416 (.A1(b[28]), .A2(a[18]), .ZN(n_815));
   OAI21_X1 i_417 (.A(n_813), .B1(n_814), .B2(n_815), .ZN(n_428));
   NAND4_X1 i_418 (.A1(a[23]), .A2(b[24]), .A3(b[23]), .A4(a[22]), .ZN(n_816));
   AOI22_X1 i_419 (.A1(b[24]), .A2(a[22]), .B1(a[23]), .B2(b[23]), .ZN(n_817));
   NAND2_X1 i_420 (.A1(b[25]), .A2(a[21]), .ZN(n_818));
   OAI21_X1 i_421 (.A(n_816), .B1(n_817), .B2(n_818), .ZN(n_429));
   INV_X1 i_422 (.A(n_811), .ZN(n_819));
   NAND2_X1 i_423 (.A1(n_819), .A2(n_810), .ZN(n_820));
   XOR2_X1 i_424 (.A(n_820), .B(n_812), .Z(n_430));
   INV_X1 i_425 (.A(n_814), .ZN(n_821));
   NAND2_X1 i_426 (.A1(n_821), .A2(n_813), .ZN(n_822));
   XOR2_X1 i_427 (.A(n_822), .B(n_815), .Z(n_431));
   INV_X1 i_428 (.A(n_817), .ZN(n_823));
   NAND2_X1 i_429 (.A1(n_823), .A2(n_816), .ZN(n_824));
   XOR2_X1 i_430 (.A(n_824), .B(n_818), .Z(n_432));
   INV_X1 i_431 (.A(n_764), .ZN(n_825));
   NAND2_X1 i_432 (.A1(n_825), .A2(n_763), .ZN(n_826));
   XOR2_X1 i_433 (.A(n_826), .B(n_765), .Z(n_433));
   INV_X1 i_434 (.A(n_768), .ZN(n_827));
   NAND2_X1 i_435 (.A1(n_827), .A2(n_767), .ZN(n_828));
   XOR2_X1 i_436 (.A(n_828), .B(n_769), .Z(n_434));
   INV_X1 i_437 (.A(n_806), .ZN(n_829));
   NAND2_X1 i_438 (.A1(n_808), .A2(n_829), .ZN(n_830));
   XOR2_X1 i_439 (.A(n_830), .B(n_809), .Z(n_435));
   NAND4_X1 i_440 (.A1(b[30]), .A2(b[29]), .A3(a[16]), .A4(a[15]), .ZN(n_831));
   AOI22_X1 i_441 (.A1(b[30]), .A2(a[15]), .B1(b[29]), .B2(a[16]), .ZN(n_832));
   NAND2_X1 i_442 (.A1(b[31]), .A2(a[14]), .ZN(n_833));
   OAI21_X1 i_443 (.A(n_831), .B1(n_832), .B2(n_833), .ZN(n_436));
   NAND4_X1 i_444 (.A1(b[27]), .A2(b[26]), .A3(a[19]), .A4(a[18]), .ZN(n_834));
   AOI22_X1 i_445 (.A1(b[27]), .A2(a[18]), .B1(b[26]), .B2(a[19]), .ZN(n_835));
   NAND2_X1 i_446 (.A1(b[28]), .A2(a[17]), .ZN(n_836));
   OAI21_X1 i_447 (.A(n_834), .B1(n_835), .B2(n_836), .ZN(n_437));
   NAND4_X1 i_448 (.A1(b[24]), .A2(b[23]), .A3(a[22]), .A4(a[21]), .ZN(n_837));
   AOI22_X1 i_449 (.A1(b[24]), .A2(a[21]), .B1(b[23]), .B2(a[22]), .ZN(n_838));
   NAND2_X1 i_450 (.A1(b[25]), .A2(a[20]), .ZN(n_839));
   OAI21_X1 i_451 (.A(n_837), .B1(n_838), .B2(n_839), .ZN(n_438));
   NAND4_X1 i_452 (.A1(a[25]), .A2(a[24]), .A3(b[21]), .A4(b[20]), .ZN(n_840));
   AOI22_X1 i_453 (.A1(a[24]), .A2(b[21]), .B1(a[25]), .B2(b[20]), .ZN(n_841));
   NAND2_X1 i_454 (.A1(a[23]), .A2(b[22]), .ZN(n_842));
   OAI21_X1 i_455 (.A(n_840), .B1(n_841), .B2(n_842), .ZN(n_439));
   NAND4_X1 i_456 (.A1(a[28]), .A2(a[27]), .A3(b[18]), .A4(b[17]), .ZN(n_843));
   AOI22_X1 i_457 (.A1(a[27]), .A2(b[18]), .B1(a[28]), .B2(b[17]), .ZN(n_844));
   NAND2_X1 i_458 (.A1(a[26]), .A2(b[19]), .ZN(n_845));
   OAI21_X1 i_459 (.A(n_843), .B1(n_844), .B2(n_845), .ZN(n_440));
   INV_X1 i_460 (.A(n_832), .ZN(n_846));
   NAND2_X1 i_461 (.A1(n_846), .A2(n_831), .ZN(n_847));
   XOR2_X1 i_462 (.A(n_847), .B(n_833), .Z(n_441));
   INV_X1 i_463 (.A(n_835), .ZN(n_848));
   NAND2_X1 i_464 (.A1(n_848), .A2(n_834), .ZN(n_849));
   XOR2_X1 i_465 (.A(n_849), .B(n_836), .Z(n_442));
   INV_X1 i_466 (.A(n_838), .ZN(n_850));
   NAND2_X1 i_467 (.A1(n_850), .A2(n_837), .ZN(n_851));
   XOR2_X1 i_468 (.A(n_851), .B(n_839), .Z(n_443));
   INV_X1 i_469 (.A(n_841), .ZN(n_852));
   NAND2_X1 i_470 (.A1(n_852), .A2(n_840), .ZN(n_853));
   XOR2_X1 i_471 (.A(n_853), .B(n_842), .Z(n_444));
   INV_X1 i_472 (.A(n_844), .ZN(n_854));
   NAND2_X1 i_473 (.A1(n_854), .A2(n_843), .ZN(n_855));
   XOR2_X1 i_474 (.A(n_855), .B(n_845), .Z(n_445));
   XOR2_X1 i_475 (.A(n_803), .B(n_804), .Z(n_856));
   NAND2_X1 i_476 (.A1(a[29]), .A2(b[16]), .ZN(n_857));
   XNOR2_X1 i_477 (.A(n_856), .B(n_857), .ZN(n_446));
   NAND4_X1 i_478 (.A1(a[26]), .A2(a[25]), .A3(b[18]), .A4(b[17]), .ZN(n_858));
   AOI22_X1 i_479 (.A1(a[25]), .A2(b[18]), .B1(a[26]), .B2(b[17]), .ZN(n_859));
   NAND2_X1 i_480 (.A1(a[24]), .A2(b[19]), .ZN(n_860));
   OAI21_X1 i_481 (.A(n_858), .B1(n_859), .B2(n_860), .ZN(n_861));
   NAND4_X1 i_482 (.A1(a[29]), .A2(a[28]), .A3(b[15]), .A4(b[14]), .ZN(n_862));
   AOI22_X1 i_483 (.A1(a[28]), .A2(b[15]), .B1(a[29]), .B2(b[14]), .ZN(n_863));
   NAND2_X1 i_484 (.A1(a[27]), .A2(b[16]), .ZN(n_864));
   OAI21_X1 i_485 (.A(n_862), .B1(n_863), .B2(n_864), .ZN(n_865));
   NOR2_X1 i_486 (.A1(n_861), .A2(n_865), .ZN(n_866));
   NAND2_X1 i_487 (.A1(a[31]), .A2(b[13]), .ZN(n_867));
   NAND2_X1 i_488 (.A1(n_861), .A2(n_865), .ZN(n_868));
   AOI21_X1 i_489 (.A(n_866), .B1(n_867), .B2(n_868), .ZN(n_447));
   NAND4_X1 i_490 (.A1(b[30]), .A2(b[29]), .A3(a[14]), .A4(a[15]), .ZN(n_869));
   AOI22_X1 i_491 (.A1(b[30]), .A2(a[14]), .B1(b[29]), .B2(a[15]), .ZN(n_870));
   NAND2_X1 i_492 (.A1(b[31]), .A2(a[13]), .ZN(n_871));
   OAI21_X1 i_493 (.A(n_869), .B1(n_870), .B2(n_871), .ZN(n_448));
   NAND4_X1 i_494 (.A1(b[27]), .A2(b[26]), .A3(a[17]), .A4(a[18]), .ZN(n_872));
   AOI22_X1 i_495 (.A1(b[27]), .A2(a[17]), .B1(b[26]), .B2(a[18]), .ZN(n_873));
   NAND2_X1 i_496 (.A1(b[28]), .A2(a[16]), .ZN(n_874));
   OAI21_X1 i_497 (.A(n_872), .B1(n_873), .B2(n_874), .ZN(n_449));
   NAND4_X1 i_498 (.A1(b[24]), .A2(b[23]), .A3(a[20]), .A4(a[21]), .ZN(n_875));
   AOI22_X1 i_499 (.A1(b[24]), .A2(a[20]), .B1(b[23]), .B2(a[21]), .ZN(n_876));
   NAND2_X1 i_500 (.A1(b[25]), .A2(a[19]), .ZN(n_877));
   OAI21_X1 i_501 (.A(n_875), .B1(n_876), .B2(n_877), .ZN(n_450));
   NAND4_X1 i_502 (.A1(a[23]), .A2(a[24]), .A3(b[21]), .A4(b[20]), .ZN(n_878));
   AOI22_X1 i_503 (.A1(a[23]), .A2(b[21]), .B1(a[24]), .B2(b[20]), .ZN(n_879));
   NAND2_X1 i_504 (.A1(a[22]), .A2(b[22]), .ZN(n_880));
   OAI21_X1 i_505 (.A(n_878), .B1(n_879), .B2(n_880), .ZN(n_451));
   NAND4_X1 i_506 (.A1(a[26]), .A2(a[27]), .A3(b[18]), .A4(b[17]), .ZN(n_881));
   AOI22_X1 i_507 (.A1(a[26]), .A2(b[18]), .B1(a[27]), .B2(b[17]), .ZN(n_882));
   NAND2_X1 i_508 (.A1(a[25]), .A2(b[19]), .ZN(n_883));
   OAI21_X1 i_509 (.A(n_881), .B1(n_882), .B2(n_883), .ZN(n_452));
   INV_X1 i_510 (.A(n_803), .ZN(n_884));
   NAND3_X1 i_511 (.A1(n_884), .A2(a[29]), .A3(b[14]), .ZN(n_885));
   AOI21_X1 i_512 (.A(n_807), .B1(a[29]), .B2(b[15]), .ZN(n_886));
   NAND2_X1 i_513 (.A1(a[28]), .A2(b[16]), .ZN(n_887));
   OAI21_X1 i_514 (.A(n_885), .B1(n_886), .B2(n_887), .ZN(n_453));
   INV_X1 i_515 (.A(n_866), .ZN(n_888));
   NAND2_X1 i_516 (.A1(n_888), .A2(n_868), .ZN(n_889));
   XOR2_X1 i_517 (.A(n_889), .B(n_867), .Z(n_454));
   INV_X1 i_518 (.A(n_870), .ZN(n_890));
   NAND2_X1 i_519 (.A1(n_890), .A2(n_869), .ZN(n_891));
   XOR2_X1 i_520 (.A(n_891), .B(n_871), .Z(n_455));
   INV_X1 i_521 (.A(n_873), .ZN(n_892));
   NAND2_X1 i_522 (.A1(n_892), .A2(n_872), .ZN(n_893));
   XOR2_X1 i_523 (.A(n_893), .B(n_874), .Z(n_456));
   INV_X1 i_524 (.A(n_876), .ZN(n_894));
   NAND2_X1 i_525 (.A1(n_894), .A2(n_875), .ZN(n_895));
   XOR2_X1 i_526 (.A(n_895), .B(n_877), .Z(n_457));
   INV_X1 i_527 (.A(n_879), .ZN(n_896));
   NAND2_X1 i_528 (.A1(n_896), .A2(n_878), .ZN(n_897));
   XOR2_X1 i_529 (.A(n_897), .B(n_880), .Z(n_458));
   INV_X1 i_530 (.A(n_882), .ZN(n_898));
   NAND2_X1 i_531 (.A1(n_898), .A2(n_881), .ZN(n_899));
   XOR2_X1 i_532 (.A(n_899), .B(n_883), .Z(n_459));
   INV_X1 i_533 (.A(n_886), .ZN(n_900));
   NAND2_X1 i_534 (.A1(n_885), .A2(n_900), .ZN(n_901));
   XOR2_X1 i_535 (.A(n_901), .B(n_887), .Z(n_460));
   NAND2_X1 i_536 (.A1(a[29]), .A2(b[13]), .ZN(n_902));
   NAND2_X1 i_537 (.A1(a[30]), .A2(b[12]), .ZN(n_903));
   NAND2_X1 i_538 (.A1(a[31]), .A2(b[11]), .ZN(n_904));
   AOI21_X1 i_539 (.A(n_902), .B1(n_903), .B2(n_904), .ZN(n_905));
   AND2_X1 i_540 (.A1(a[30]), .A2(b[11]), .ZN(n_906));
   OAI211_X1 i_541 (.A(a[31]), .B(b[12]), .C1(n_905), .C2(n_906), .ZN(n_907));
   AOI21_X1 i_542 (.A(n_905), .B1(a[31]), .B2(b[12]), .ZN(n_908));
   NAND2_X1 i_543 (.A1(a[30]), .A2(b[13]), .ZN(n_909));
   OAI21_X1 i_544 (.A(n_907), .B1(n_908), .B2(n_909), .ZN(n_461));
   NAND4_X1 i_545 (.A1(b[30]), .A2(b[29]), .A3(a[14]), .A4(a[13]), .ZN(n_910));
   AOI22_X1 i_546 (.A1(b[30]), .A2(a[13]), .B1(b[29]), .B2(a[14]), .ZN(n_911));
   NAND2_X1 i_547 (.A1(b[31]), .A2(a[12]), .ZN(n_912));
   OAI21_X1 i_548 (.A(n_910), .B1(n_911), .B2(n_912), .ZN(n_462));
   NAND4_X1 i_549 (.A1(b[27]), .A2(b[26]), .A3(a[17]), .A4(a[16]), .ZN(n_913));
   AOI22_X1 i_550 (.A1(b[27]), .A2(a[16]), .B1(b[26]), .B2(a[17]), .ZN(n_914));
   NAND2_X1 i_551 (.A1(b[28]), .A2(a[15]), .ZN(n_915));
   OAI21_X1 i_552 (.A(n_913), .B1(n_914), .B2(n_915), .ZN(n_463));
   NAND4_X1 i_553 (.A1(b[24]), .A2(b[23]), .A3(a[20]), .A4(a[19]), .ZN(n_916));
   AOI22_X1 i_554 (.A1(b[24]), .A2(a[19]), .B1(b[23]), .B2(a[20]), .ZN(n_917));
   NAND2_X1 i_555 (.A1(b[25]), .A2(a[18]), .ZN(n_918));
   OAI21_X1 i_556 (.A(n_916), .B1(n_917), .B2(n_918), .ZN(n_464));
   NAND4_X1 i_557 (.A1(a[23]), .A2(a[22]), .A3(b[21]), .A4(b[20]), .ZN(n_919));
   AOI22_X1 i_558 (.A1(a[22]), .A2(b[21]), .B1(a[23]), .B2(b[20]), .ZN(n_920));
   NAND2_X1 i_559 (.A1(b[22]), .A2(a[21]), .ZN(n_921));
   OAI21_X1 i_560 (.A(n_919), .B1(n_920), .B2(n_921), .ZN(n_465));
   INV_X1 i_561 (.A(n_911), .ZN(n_922));
   NAND2_X1 i_562 (.A1(n_922), .A2(n_910), .ZN(n_923));
   XOR2_X1 i_563 (.A(n_923), .B(n_912), .Z(n_466));
   INV_X1 i_564 (.A(n_914), .ZN(n_924));
   NAND2_X1 i_565 (.A1(n_924), .A2(n_913), .ZN(n_925));
   XOR2_X1 i_566 (.A(n_925), .B(n_915), .Z(n_467));
   INV_X1 i_567 (.A(n_917), .ZN(n_926));
   NAND2_X1 i_568 (.A1(n_926), .A2(n_916), .ZN(n_927));
   XOR2_X1 i_569 (.A(n_927), .B(n_918), .Z(n_468));
   INV_X1 i_570 (.A(n_920), .ZN(n_928));
   NAND2_X1 i_571 (.A1(n_928), .A2(n_919), .ZN(n_929));
   XOR2_X1 i_572 (.A(n_929), .B(n_921), .Z(n_469));
   INV_X1 i_573 (.A(n_859), .ZN(n_930));
   NAND2_X1 i_574 (.A1(n_930), .A2(n_858), .ZN(n_931));
   XOR2_X1 i_575 (.A(n_931), .B(n_860), .Z(n_470));
   INV_X1 i_576 (.A(n_863), .ZN(n_932));
   NAND2_X1 i_577 (.A1(n_932), .A2(n_862), .ZN(n_933));
   XOR2_X1 i_578 (.A(n_933), .B(n_864), .Z(n_471));
   INV_X1 i_579 (.A(n_908), .ZN(n_934));
   NAND2_X1 i_580 (.A1(n_907), .A2(n_934), .ZN(n_935));
   XOR2_X1 i_581 (.A(n_935), .B(n_909), .Z(n_472));
   NAND4_X1 i_582 (.A1(b[30]), .A2(b[29]), .A3(a[13]), .A4(a[12]), .ZN(n_936));
   AOI22_X1 i_583 (.A1(b[30]), .A2(a[12]), .B1(b[29]), .B2(a[13]), .ZN(n_937));
   NAND2_X1 i_584 (.A1(b[31]), .A2(a[11]), .ZN(n_938));
   OAI21_X1 i_585 (.A(n_936), .B1(n_937), .B2(n_938), .ZN(n_473));
   NAND4_X1 i_586 (.A1(b[27]), .A2(b[26]), .A3(a[16]), .A4(a[15]), .ZN(n_939));
   AOI22_X1 i_587 (.A1(b[27]), .A2(a[15]), .B1(b[26]), .B2(a[16]), .ZN(n_940));
   NAND2_X1 i_588 (.A1(b[28]), .A2(a[14]), .ZN(n_941));
   OAI21_X1 i_589 (.A(n_939), .B1(n_940), .B2(n_941), .ZN(n_474));
   NAND4_X1 i_590 (.A1(b[24]), .A2(b[23]), .A3(a[19]), .A4(a[18]), .ZN(n_942));
   AOI22_X1 i_591 (.A1(b[24]), .A2(a[18]), .B1(b[23]), .B2(a[19]), .ZN(n_943));
   NAND2_X1 i_592 (.A1(b[25]), .A2(a[17]), .ZN(n_944));
   OAI21_X1 i_593 (.A(n_942), .B1(n_943), .B2(n_944), .ZN(n_475));
   NAND4_X1 i_594 (.A1(a[22]), .A2(a[21]), .A3(b[21]), .A4(b[20]), .ZN(n_945));
   AOI22_X1 i_595 (.A1(a[21]), .A2(b[21]), .B1(a[22]), .B2(b[20]), .ZN(n_946));
   NAND2_X1 i_596 (.A1(b[22]), .A2(a[20]), .ZN(n_947));
   OAI21_X1 i_597 (.A(n_945), .B1(n_946), .B2(n_947), .ZN(n_476));
   NAND4_X1 i_598 (.A1(a[25]), .A2(a[24]), .A3(b[18]), .A4(b[17]), .ZN(n_948));
   AOI22_X1 i_599 (.A1(a[24]), .A2(b[18]), .B1(a[25]), .B2(b[17]), .ZN(n_949));
   NAND2_X1 i_600 (.A1(a[23]), .A2(b[19]), .ZN(n_950));
   OAI21_X1 i_601 (.A(n_948), .B1(n_949), .B2(n_950), .ZN(n_477));
   NAND4_X1 i_602 (.A1(a[28]), .A2(a[27]), .A3(b[15]), .A4(b[14]), .ZN(n_951));
   AOI22_X1 i_603 (.A1(a[27]), .A2(b[15]), .B1(a[28]), .B2(b[14]), .ZN(n_952));
   NAND2_X1 i_604 (.A1(a[26]), .A2(b[16]), .ZN(n_953));
   OAI21_X1 i_605 (.A(n_951), .B1(n_952), .B2(n_953), .ZN(n_478));
   INV_X1 i_606 (.A(n_937), .ZN(n_954));
   NAND2_X1 i_607 (.A1(n_954), .A2(n_936), .ZN(n_955));
   XOR2_X1 i_608 (.A(n_955), .B(n_938), .Z(n_479));
   INV_X1 i_609 (.A(n_940), .ZN(n_956));
   NAND2_X1 i_610 (.A1(n_956), .A2(n_939), .ZN(n_957));
   XOR2_X1 i_611 (.A(n_957), .B(n_941), .Z(n_480));
   INV_X1 i_612 (.A(n_943), .ZN(n_958));
   NAND2_X1 i_613 (.A1(n_958), .A2(n_942), .ZN(n_959));
   XOR2_X1 i_614 (.A(n_959), .B(n_944), .Z(n_481));
   INV_X1 i_615 (.A(n_946), .ZN(n_960));
   NAND2_X1 i_616 (.A1(n_960), .A2(n_945), .ZN(n_961));
   XOR2_X1 i_617 (.A(n_961), .B(n_947), .Z(n_482));
   INV_X1 i_618 (.A(n_949), .ZN(n_962));
   NAND2_X1 i_619 (.A1(n_962), .A2(n_948), .ZN(n_963));
   XOR2_X1 i_620 (.A(n_963), .B(n_950), .Z(n_483));
   INV_X1 i_621 (.A(n_952), .ZN(n_964));
   NAND2_X1 i_622 (.A1(n_964), .A2(n_951), .ZN(n_965));
   XOR2_X1 i_623 (.A(n_965), .B(n_953), .Z(n_484));
   XNOR2_X1 i_624 (.A(n_903), .B(n_904), .ZN(n_966));
   XOR2_X1 i_625 (.A(n_966), .B(n_902), .Z(n_485));
   NAND4_X1 i_626 (.A1(a[26]), .A2(a[25]), .A3(b[15]), .A4(b[14]), .ZN(n_967));
   AOI22_X1 i_627 (.A1(a[25]), .A2(b[15]), .B1(a[26]), .B2(b[14]), .ZN(n_968));
   NAND2_X1 i_628 (.A1(a[24]), .A2(b[16]), .ZN(n_969));
   OAI21_X1 i_629 (.A(n_967), .B1(n_968), .B2(n_969), .ZN(n_970));
   NAND4_X1 i_630 (.A1(a[29]), .A2(a[28]), .A3(b[12]), .A4(b[11]), .ZN(n_971));
   AOI22_X1 i_631 (.A1(a[28]), .A2(b[12]), .B1(a[29]), .B2(b[11]), .ZN(n_972));
   NAND2_X1 i_632 (.A1(a[27]), .A2(b[13]), .ZN(n_973));
   OAI21_X1 i_633 (.A(n_971), .B1(n_972), .B2(n_973), .ZN(n_974));
   NOR2_X1 i_634 (.A1(n_970), .A2(n_974), .ZN(n_975));
   NAND2_X1 i_635 (.A1(a[31]), .A2(b[10]), .ZN(n_976));
   NAND2_X1 i_636 (.A1(n_970), .A2(n_974), .ZN(n_977));
   AOI21_X1 i_637 (.A(n_975), .B1(n_976), .B2(n_977), .ZN(n_486));
   NAND4_X1 i_638 (.A1(b[30]), .A2(b[29]), .A3(a[11]), .A4(a[12]), .ZN(n_978));
   AOI22_X1 i_639 (.A1(b[30]), .A2(a[11]), .B1(b[29]), .B2(a[12]), .ZN(n_979));
   NAND2_X1 i_640 (.A1(b[31]), .A2(a[10]), .ZN(n_980));
   OAI21_X1 i_641 (.A(n_978), .B1(n_979), .B2(n_980), .ZN(n_3787));
   NAND4_X1 i_642 (.A1(b[27]), .A2(b[26]), .A3(a[14]), .A4(a[15]), .ZN(n_981));
   AOI22_X1 i_643 (.A1(b[27]), .A2(a[14]), .B1(b[26]), .B2(a[15]), .ZN(n_982));
   NAND2_X1 i_644 (.A1(b[28]), .A2(a[13]), .ZN(n_983));
   OAI21_X1 i_645 (.A(n_981), .B1(n_982), .B2(n_983), .ZN(n_3794));
   NAND4_X1 i_646 (.A1(b[24]), .A2(b[23]), .A3(a[17]), .A4(a[18]), .ZN(n_984));
   AOI22_X1 i_647 (.A1(b[24]), .A2(a[17]), .B1(b[23]), .B2(a[18]), .ZN(n_985));
   NAND2_X1 i_648 (.A1(b[25]), .A2(a[16]), .ZN(n_986));
   OAI21_X1 i_649 (.A(n_984), .B1(n_985), .B2(n_986), .ZN(n_3801));
   NAND4_X1 i_650 (.A1(a[20]), .A2(a[21]), .A3(b[21]), .A4(b[20]), .ZN(n_987));
   AOI22_X1 i_651 (.A1(a[20]), .A2(b[21]), .B1(a[21]), .B2(b[20]), .ZN(n_988));
   NAND2_X1 i_652 (.A1(b[22]), .A2(a[19]), .ZN(n_989));
   OAI21_X1 i_653 (.A(n_987), .B1(n_988), .B2(n_989), .ZN(n_3808));
   NAND4_X1 i_654 (.A1(a[23]), .A2(a[24]), .A3(b[18]), .A4(b[17]), .ZN(n_990));
   AOI22_X1 i_655 (.A1(a[23]), .A2(b[18]), .B1(a[24]), .B2(b[17]), .ZN(n_991));
   NAND2_X1 i_656 (.A1(a[22]), .A2(b[19]), .ZN(n_992));
   OAI21_X1 i_657 (.A(n_990), .B1(n_991), .B2(n_992), .ZN(n_3815));
   NAND4_X1 i_658 (.A1(a[26]), .A2(a[27]), .A3(b[15]), .A4(b[14]), .ZN(n_993));
   AOI22_X1 i_659 (.A1(a[26]), .A2(b[15]), .B1(a[27]), .B2(b[14]), .ZN(n_994));
   NAND2_X1 i_660 (.A1(a[25]), .A2(b[16]), .ZN(n_995));
   OAI21_X1 i_661 (.A(n_993), .B1(n_994), .B2(n_995), .ZN(n_487));
   INV_X1 i_662 (.A(n_903), .ZN(n_996));
   NAND3_X1 i_663 (.A1(n_996), .A2(a[29]), .A3(b[11]), .ZN(n_997));
   AOI21_X1 i_664 (.A(n_906), .B1(a[29]), .B2(b[12]), .ZN(n_998));
   NAND2_X1 i_665 (.A1(a[28]), .A2(b[13]), .ZN(n_999));
   OAI21_X1 i_666 (.A(n_997), .B1(n_998), .B2(n_999), .ZN(n_488));
   INV_X1 i_667 (.A(n_975), .ZN(n_1000));
   NAND2_X1 i_668 (.A1(n_1000), .A2(n_977), .ZN(n_1001));
   XOR2_X1 i_669 (.A(n_1001), .B(n_976), .Z(n_489));
   INV_X1 i_670 (.A(n_979), .ZN(n_1002));
   NAND2_X1 i_671 (.A1(n_1002), .A2(n_978), .ZN(n_1003));
   XOR2_X1 i_672 (.A(n_1003), .B(n_980), .Z(n_3786));
   INV_X1 i_673 (.A(n_982), .ZN(n_1004));
   NAND2_X1 i_674 (.A1(n_1004), .A2(n_981), .ZN(n_1005));
   XOR2_X1 i_675 (.A(n_1005), .B(n_983), .Z(n_3793));
   INV_X1 i_676 (.A(n_985), .ZN(n_1006));
   NAND2_X1 i_677 (.A1(n_1006), .A2(n_984), .ZN(n_1007));
   XOR2_X1 i_678 (.A(n_1007), .B(n_986), .Z(n_3800));
   INV_X1 i_679 (.A(n_988), .ZN(n_1008));
   NAND2_X1 i_680 (.A1(n_1008), .A2(n_987), .ZN(n_1009));
   XOR2_X1 i_681 (.A(n_1009), .B(n_989), .Z(n_3807));
   INV_X1 i_682 (.A(n_991), .ZN(n_1010));
   NAND2_X1 i_683 (.A1(n_1010), .A2(n_990), .ZN(n_1011));
   XOR2_X1 i_684 (.A(n_1011), .B(n_992), .Z(n_3814));
   INV_X1 i_685 (.A(n_994), .ZN(n_1012));
   NAND2_X1 i_686 (.A1(n_1012), .A2(n_993), .ZN(n_1013));
   XOR2_X1 i_687 (.A(n_1013), .B(n_995), .Z(n_490));
   INV_X1 i_688 (.A(n_998), .ZN(n_1014));
   NAND2_X1 i_689 (.A1(n_997), .A2(n_1014), .ZN(n_1015));
   XOR2_X1 i_690 (.A(n_1015), .B(n_999), .Z(n_491));
   NAND4_X1 i_691 (.A1(b[30]), .A2(b[29]), .A3(a[11]), .A4(a[10]), .ZN(n_1016));
   AOI22_X1 i_692 (.A1(b[30]), .A2(a[10]), .B1(b[29]), .B2(a[11]), .ZN(n_1017));
   NAND2_X1 i_693 (.A1(b[31]), .A2(a[9]), .ZN(n_1018));
   OAI21_X1 i_694 (.A(n_1016), .B1(n_1017), .B2(n_1018), .ZN(n_3702));
   NAND4_X1 i_695 (.A1(b[27]), .A2(b[26]), .A3(a[14]), .A4(a[13]), .ZN(n_1019));
   AOI22_X1 i_696 (.A1(b[27]), .A2(a[13]), .B1(b[26]), .B2(a[14]), .ZN(n_1020));
   NAND2_X1 i_697 (.A1(b[28]), .A2(a[12]), .ZN(n_1021));
   OAI21_X1 i_698 (.A(n_1019), .B1(n_1020), .B2(n_1021), .ZN(n_3709));
   NAND4_X1 i_699 (.A1(b[24]), .A2(b[23]), .A3(a[17]), .A4(a[16]), .ZN(n_1022));
   AOI22_X1 i_700 (.A1(b[24]), .A2(a[16]), .B1(b[23]), .B2(a[17]), .ZN(n_1023));
   NAND2_X1 i_701 (.A1(b[25]), .A2(a[15]), .ZN(n_1024));
   OAI21_X1 i_702 (.A(n_1022), .B1(n_1023), .B2(n_1024), .ZN(n_3716));
   NAND4_X1 i_703 (.A1(a[20]), .A2(b[21]), .A3(b[20]), .A4(a[19]), .ZN(n_1025));
   AOI22_X1 i_704 (.A1(b[21]), .A2(a[19]), .B1(a[20]), .B2(b[20]), .ZN(n_1026));
   NAND2_X1 i_705 (.A1(b[22]), .A2(a[18]), .ZN(n_1027));
   OAI21_X1 i_706 (.A(n_1025), .B1(n_1026), .B2(n_1027), .ZN(n_3723));
   NAND4_X1 i_707 (.A1(a[23]), .A2(a[22]), .A3(b[18]), .A4(b[17]), .ZN(n_1028));
   AOI22_X1 i_708 (.A1(a[22]), .A2(b[18]), .B1(a[23]), .B2(b[17]), .ZN(n_1031));
   NAND2_X1 i_709 (.A1(a[21]), .A2(b[19]), .ZN(n_1032));
   OAI21_X1 i_710 (.A(n_1028), .B1(n_1031), .B2(n_1032), .ZN(n_3730));
   INV_X1 i_711 (.A(n_1017), .ZN(n_1033));
   NAND2_X1 i_712 (.A1(n_1033), .A2(n_1016), .ZN(n_1035));
   XOR2_X1 i_713 (.A(n_1035), .B(n_1018), .Z(n_3701));
   INV_X1 i_714 (.A(n_1020), .ZN(n_1036));
   NAND2_X1 i_715 (.A1(n_1036), .A2(n_1019), .ZN(n_1037));
   XOR2_X1 i_716 (.A(n_1037), .B(n_1021), .Z(n_3708));
   INV_X1 i_717 (.A(n_1023), .ZN(n_1038));
   NAND2_X1 i_718 (.A1(n_1038), .A2(n_1022), .ZN(n_1041));
   XOR2_X1 i_719 (.A(n_1041), .B(n_1024), .Z(n_3715));
   INV_X1 i_720 (.A(n_1026), .ZN(n_1042));
   NAND2_X1 i_721 (.A1(n_1042), .A2(n_1025), .ZN(n_1043));
   XOR2_X1 i_722 (.A(n_1043), .B(n_1027), .Z(n_3722));
   INV_X1 i_723 (.A(n_1031), .ZN(n_1044));
   NAND2_X1 i_724 (.A1(n_1044), .A2(n_1028), .ZN(n_1047));
   XOR2_X1 i_725 (.A(n_1047), .B(n_1032), .Z(n_3729));
   INV_X1 i_726 (.A(n_968), .ZN(n_1048));
   NAND2_X1 i_727 (.A1(n_1048), .A2(n_967), .ZN(n_1049));
   XOR2_X1 i_728 (.A(n_1049), .B(n_969), .Z(n_3736));
   INV_X1 i_729 (.A(n_972), .ZN(n_1050));
   NAND2_X1 i_730 (.A1(n_1050), .A2(n_971), .ZN(n_1051));
   XOR2_X1 i_731 (.A(n_1051), .B(n_973), .Z(n_3743));
   INV_X1 i_732 (.A(b[10]), .ZN(n_1054));
   NAND2_X1 i_733 (.A1(a[30]), .A2(b[9]), .ZN(n_1055));
   NAND2_X1 i_734 (.A1(a[31]), .A2(b[8]), .ZN(n_1057));
   AOI211_X1 i_735 (.A(n_497), .B(n_1054), .C1(n_1055), .C2(n_1057), .ZN(n_1058));
   INV_X1 i_736 (.A(b[8]), .ZN(n_1059));
   NOR2_X1 i_737 (.A1(n_659), .A2(n_1059), .ZN(n_1060));
   OAI211_X1 i_738 (.A(a[31]), .B(b[9]), .C1(n_1058), .C2(n_1060), .ZN(n_1061));
   AOI21_X1 i_739 (.A(n_1058), .B1(a[31]), .B2(b[9]), .ZN(n_1062));
   NAND2_X1 i_740 (.A1(a[30]), .A2(b[10]), .ZN(n_1064));
   OAI21_X1 i_741 (.A(n_1061), .B1(n_1062), .B2(n_1064), .ZN(n_3750));
   AND2_X1 i_742 (.A1(n_1062), .A2(n_1064), .ZN(n_1065));
   OAI22_X1 i_743 (.A1(n_1061), .A2(n_1064), .B1(n_3750), .B2(n_1065), .ZN(
      n_3749));
   NAND4_X1 i_744 (.A1(b[30]), .A2(b[29]), .A3(a[10]), .A4(a[9]), .ZN(n_1066));
   AOI22_X1 i_745 (.A1(b[30]), .A2(a[9]), .B1(b[29]), .B2(a[10]), .ZN(n_1067));
   NAND2_X1 i_746 (.A1(b[31]), .A2(a[8]), .ZN(n_1072));
   OAI21_X1 i_747 (.A(n_1066), .B1(n_1067), .B2(n_1072), .ZN(n_3616));
   NAND4_X1 i_748 (.A1(b[27]), .A2(b[26]), .A3(a[13]), .A4(a[12]), .ZN(n_1073));
   AOI22_X1 i_749 (.A1(b[27]), .A2(a[12]), .B1(b[26]), .B2(a[13]), .ZN(n_1076));
   NAND2_X1 i_750 (.A1(b[28]), .A2(a[11]), .ZN(n_1077));
   OAI21_X1 i_751 (.A(n_1073), .B1(n_1076), .B2(n_1077), .ZN(n_3623));
   NAND4_X1 i_752 (.A1(b[24]), .A2(b[23]), .A3(a[16]), .A4(a[15]), .ZN(n_1078));
   AOI22_X1 i_753 (.A1(b[24]), .A2(a[15]), .B1(b[23]), .B2(a[16]), .ZN(n_1079));
   NAND2_X1 i_754 (.A1(b[25]), .A2(a[14]), .ZN(n_1080));
   OAI21_X1 i_755 (.A(n_1078), .B1(n_1079), .B2(n_1080), .ZN(n_3630));
   NAND4_X1 i_756 (.A1(b[21]), .A2(b[20]), .A3(a[19]), .A4(a[18]), .ZN(n_1082));
   AOI22_X1 i_757 (.A1(b[21]), .A2(a[18]), .B1(b[20]), .B2(a[19]), .ZN(n_1083));
   NAND2_X1 i_758 (.A1(b[22]), .A2(a[17]), .ZN(n_1084));
   OAI21_X1 i_759 (.A(n_1082), .B1(n_1083), .B2(n_1084), .ZN(n_3637));
   NAND4_X1 i_760 (.A1(a[22]), .A2(a[21]), .A3(b[18]), .A4(b[17]), .ZN(n_1085));
   AOI22_X1 i_761 (.A1(a[21]), .A2(b[18]), .B1(a[22]), .B2(b[17]), .ZN(n_1086));
   NAND2_X1 i_762 (.A1(a[20]), .A2(b[19]), .ZN(n_1087));
   OAI21_X1 i_763 (.A(n_1085), .B1(n_1086), .B2(n_1087), .ZN(n_3644));
   NAND4_X1 i_764 (.A1(a[25]), .A2(a[24]), .A3(b[15]), .A4(b[14]), .ZN(n_1090));
   AOI22_X1 i_765 (.A1(a[24]), .A2(b[15]), .B1(a[25]), .B2(b[14]), .ZN(n_1091));
   NAND2_X1 i_766 (.A1(a[23]), .A2(b[16]), .ZN(n_1092));
   OAI21_X1 i_767 (.A(n_1090), .B1(n_1091), .B2(n_1092), .ZN(n_3651));
   NAND4_X1 i_768 (.A1(a[28]), .A2(a[27]), .A3(b[12]), .A4(b[11]), .ZN(n_1093));
   AOI22_X1 i_769 (.A1(a[27]), .A2(b[12]), .B1(a[28]), .B2(b[11]), .ZN(n_1098));
   NAND2_X1 i_770 (.A1(a[26]), .A2(b[13]), .ZN(n_1099));
   OAI21_X1 i_771 (.A(n_1093), .B1(n_1098), .B2(n_1099), .ZN(n_3658));
   INV_X1 i_772 (.A(n_1067), .ZN(n_1102));
   NAND2_X1 i_773 (.A1(n_1102), .A2(n_1066), .ZN(n_1103));
   XOR2_X1 i_774 (.A(n_1103), .B(n_1072), .Z(n_3615));
   INV_X1 i_775 (.A(n_1076), .ZN(n_1104));
   NAND2_X1 i_776 (.A1(n_1104), .A2(n_1073), .ZN(n_1105));
   XOR2_X1 i_777 (.A(n_1105), .B(n_1077), .Z(n_3622));
   INV_X1 i_778 (.A(n_1079), .ZN(n_1106));
   NAND2_X1 i_779 (.A1(n_1106), .A2(n_1078), .ZN(n_1109));
   XOR2_X1 i_780 (.A(n_1109), .B(n_1080), .Z(n_3629));
   INV_X1 i_781 (.A(n_1083), .ZN(n_1110));
   NAND2_X1 i_782 (.A1(n_1110), .A2(n_1082), .ZN(n_1111));
   XOR2_X1 i_783 (.A(n_1111), .B(n_1084), .Z(n_3636));
   INV_X1 i_784 (.A(n_1086), .ZN(n_1112));
   NAND2_X1 i_785 (.A1(n_1112), .A2(n_1085), .ZN(n_1115));
   XOR2_X1 i_786 (.A(n_1115), .B(n_1087), .Z(n_3643));
   INV_X1 i_787 (.A(n_1091), .ZN(n_1116));
   NAND2_X1 i_788 (.A1(n_1116), .A2(n_1090), .ZN(n_1117));
   XOR2_X1 i_789 (.A(n_1117), .B(n_1092), .Z(n_3650));
   INV_X1 i_790 (.A(n_1098), .ZN(n_1118));
   NAND2_X1 i_791 (.A1(n_1118), .A2(n_1093), .ZN(n_1119));
   XOR2_X1 i_792 (.A(n_1119), .B(n_1099), .Z(n_3657));
   XOR2_X1 i_793 (.A(n_1055), .B(n_1057), .Z(n_1126));
   NAND2_X1 i_794 (.A1(a[29]), .A2(b[10]), .ZN(n_1127));
   XNOR2_X1 i_795 (.A(n_1126), .B(n_1127), .ZN(n_3664));
   NOR2_X1 i_796 (.A1(n_497), .A2(n_1059), .ZN(n_1130));
   NAND3_X1 i_797 (.A1(n_1130), .A2(a[28]), .A3(b[9]), .ZN(n_1131));
   AOI21_X1 i_798 (.A(n_1130), .B1(a[28]), .B2(b[9]), .ZN(n_1132));
   NAND2_X1 i_799 (.A1(a[27]), .A2(b[10]), .ZN(n_1133));
   OAI21_X1 i_800 (.A(n_1131), .B1(n_1132), .B2(n_1133), .ZN(n_1134));
   NAND4_X1 i_801 (.A1(a[26]), .A2(a[25]), .A3(b[12]), .A4(b[11]), .ZN(n_1136));
   AOI22_X1 i_802 (.A1(a[25]), .A2(b[12]), .B1(a[26]), .B2(b[11]), .ZN(n_1137));
   NAND2_X1 i_803 (.A1(a[24]), .A2(b[13]), .ZN(n_1138));
   OAI21_X1 i_804 (.A(n_1136), .B1(n_1137), .B2(n_1138), .ZN(n_1139));
   NOR2_X1 i_805 (.A1(n_1134), .A2(n_1139), .ZN(n_1140));
   NAND2_X1 i_806 (.A1(a[31]), .A2(b[7]), .ZN(n_1141));
   NAND2_X1 i_807 (.A1(n_1134), .A2(n_1139), .ZN(n_1143));
   AOI21_X1 i_808 (.A(n_1140), .B1(n_1141), .B2(n_1143), .ZN(n_3578));
   NAND4_X1 i_809 (.A1(b[30]), .A2(b[29]), .A3(a[8]), .A4(a[9]), .ZN(n_1144));
   AOI22_X1 i_810 (.A1(b[30]), .A2(a[8]), .B1(b[29]), .B2(a[9]), .ZN(n_1145));
   NAND2_X1 i_811 (.A1(b[31]), .A2(a[7]), .ZN(n_1146));
   OAI21_X1 i_812 (.A(n_1144), .B1(n_1145), .B2(n_1146), .ZN(n_3522));
   NAND4_X1 i_813 (.A1(b[27]), .A2(b[26]), .A3(a[11]), .A4(a[12]), .ZN(n_1155));
   AOI22_X1 i_814 (.A1(b[27]), .A2(a[11]), .B1(b[26]), .B2(a[12]), .ZN(n_1156));
   NAND2_X1 i_815 (.A1(b[28]), .A2(a[10]), .ZN(n_1159));
   OAI21_X1 i_816 (.A(n_1155), .B1(n_1156), .B2(n_1159), .ZN(n_3529));
   NAND4_X1 i_817 (.A1(b[24]), .A2(b[23]), .A3(a[14]), .A4(a[15]), .ZN(n_1160));
   AOI22_X1 i_818 (.A1(b[24]), .A2(a[14]), .B1(b[23]), .B2(a[15]), .ZN(n_1161));
   NAND2_X1 i_819 (.A1(b[25]), .A2(a[13]), .ZN(n_1162));
   OAI21_X1 i_820 (.A(n_1160), .B1(n_1161), .B2(n_1162), .ZN(n_3536));
   NAND4_X1 i_821 (.A1(b[21]), .A2(b[20]), .A3(a[17]), .A4(a[18]), .ZN(n_1163));
   AOI22_X1 i_822 (.A1(b[21]), .A2(a[17]), .B1(b[20]), .B2(a[18]), .ZN(n_1166));
   NAND2_X1 i_823 (.A1(b[22]), .A2(a[16]), .ZN(n_1167));
   OAI21_X1 i_824 (.A(n_1163), .B1(n_1166), .B2(n_1167), .ZN(n_3543));
   NAND4_X1 i_825 (.A1(a[20]), .A2(a[21]), .A3(b[18]), .A4(b[17]), .ZN(n_1168));
   AOI22_X1 i_826 (.A1(a[20]), .A2(b[18]), .B1(a[21]), .B2(b[17]), .ZN(n_1169));
   NAND2_X1 i_827 (.A1(a[19]), .A2(b[19]), .ZN(n_1170));
   OAI21_X1 i_828 (.A(n_1168), .B1(n_1169), .B2(n_1170), .ZN(n_3550));
   NAND4_X1 i_829 (.A1(a[23]), .A2(a[24]), .A3(b[15]), .A4(b[14]), .ZN(n_1172));
   AOI22_X1 i_830 (.A1(a[23]), .A2(b[15]), .B1(a[24]), .B2(b[14]), .ZN(n_1173));
   NAND2_X1 i_831 (.A1(a[22]), .A2(b[16]), .ZN(n_1174));
   OAI21_X1 i_832 (.A(n_1172), .B1(n_1173), .B2(n_1174), .ZN(n_3557));
   NAND4_X1 i_833 (.A1(a[26]), .A2(a[27]), .A3(b[12]), .A4(b[11]), .ZN(n_1175));
   AOI22_X1 i_834 (.A1(a[26]), .A2(b[12]), .B1(a[27]), .B2(b[11]), .ZN(n_1176));
   NAND2_X1 i_835 (.A1(a[25]), .A2(b[13]), .ZN(n_1177));
   OAI21_X1 i_836 (.A(n_1175), .B1(n_1176), .B2(n_1177), .ZN(n_3564));
   INV_X1 i_837 (.A(n_1055), .ZN(n_1180));
   NAND2_X1 i_838 (.A1(n_1180), .A2(n_1130), .ZN(n_1181));
   AOI21_X1 i_839 (.A(n_1060), .B1(a[29]), .B2(b[9]), .ZN(n_1182));
   NAND2_X1 i_840 (.A1(a[28]), .A2(b[10]), .ZN(n_1183));
   OAI21_X1 i_841 (.A(n_1181), .B1(n_1182), .B2(n_1183), .ZN(n_3571));
   INV_X1 i_842 (.A(n_1140), .ZN(n_1192));
   NAND2_X1 i_843 (.A1(n_1143), .A2(n_1192), .ZN(n_1193));
   XOR2_X1 i_844 (.A(n_1193), .B(n_1141), .Z(n_3577));
   INV_X1 i_845 (.A(n_1145), .ZN(n_1196));
   NAND2_X1 i_846 (.A1(n_1196), .A2(n_1144), .ZN(n_1197));
   XOR2_X1 i_847 (.A(n_1197), .B(n_1146), .Z(n_3521));
   INV_X1 i_848 (.A(n_1156), .ZN(n_1198));
   NAND2_X1 i_849 (.A1(n_1198), .A2(n_1155), .ZN(n_1199));
   XOR2_X1 i_850 (.A(n_1199), .B(n_1159), .Z(n_3528));
   INV_X1 i_851 (.A(n_1161), .ZN(n_1200));
   NAND2_X1 i_852 (.A1(n_1200), .A2(n_1160), .ZN(n_1203));
   XOR2_X1 i_853 (.A(n_1203), .B(n_1162), .Z(n_3535));
   INV_X1 i_854 (.A(n_1166), .ZN(n_1204));
   NAND2_X1 i_855 (.A1(n_1204), .A2(n_1163), .ZN(n_1205));
   XOR2_X1 i_856 (.A(n_1205), .B(n_1167), .Z(n_3542));
   INV_X1 i_857 (.A(n_1169), .ZN(n_1206));
   NAND2_X1 i_858 (.A1(n_1206), .A2(n_1168), .ZN(n_1207));
   XOR2_X1 i_859 (.A(n_1207), .B(n_1170), .Z(n_3549));
   INV_X1 i_860 (.A(n_1173), .ZN(n_1210));
   NAND2_X1 i_861 (.A1(n_1210), .A2(n_1172), .ZN(n_1211));
   XOR2_X1 i_862 (.A(n_1211), .B(n_1174), .Z(n_3556));
   INV_X1 i_863 (.A(n_1176), .ZN(n_1212));
   NAND2_X1 i_864 (.A1(n_1212), .A2(n_1175), .ZN(n_1213));
   XOR2_X1 i_865 (.A(n_1213), .B(n_1177), .Z(n_3563));
   INV_X1 i_866 (.A(n_1182), .ZN(n_1216));
   NAND2_X1 i_867 (.A1(n_1181), .A2(n_1216), .ZN(n_1217));
   XOR2_X1 i_868 (.A(n_1217), .B(n_1183), .Z(n_3570));
   NAND2_X1 i_869 (.A1(a[29]), .A2(b[7]), .ZN(n_1218));
   NAND2_X1 i_870 (.A1(a[30]), .A2(b[6]), .ZN(n_1219));
   NAND2_X1 i_871 (.A1(a[31]), .A2(b[5]), .ZN(n_1220));
   AOI21_X1 i_872 (.A(n_1218), .B1(n_1219), .B2(n_1220), .ZN(n_1231));
   INV_X1 i_873 (.A(b[5]), .ZN(n_1232));
   NOR2_X1 i_874 (.A1(n_659), .A2(n_1232), .ZN(n_1235));
   OAI211_X1 i_875 (.A(a[31]), .B(b[6]), .C1(n_1231), .C2(n_1235), .ZN(n_1236));
   AOI21_X1 i_876 (.A(n_1231), .B1(a[31]), .B2(b[6]), .ZN(n_1237));
   NAND2_X1 i_877 (.A1(a[30]), .A2(b[7]), .ZN(n_1238));
   OAI21_X1 i_878 (.A(n_1236), .B1(n_1237), .B2(n_1238), .ZN(n_3481));
   NAND4_X1 i_879 (.A1(b[30]), .A2(b[29]), .A3(a[8]), .A4(a[7]), .ZN(n_1239));
   AOI22_X1 i_880 (.A1(b[30]), .A2(a[7]), .B1(b[29]), .B2(a[8]), .ZN(n_1242));
   NAND2_X1 i_881 (.A1(b[31]), .A2(a[6]), .ZN(n_1243));
   OAI21_X1 i_882 (.A(n_1239), .B1(n_1242), .B2(n_1243), .ZN(n_3426));
   NAND4_X1 i_883 (.A1(b[27]), .A2(b[26]), .A3(a[11]), .A4(a[10]), .ZN(n_1244));
   AOI22_X1 i_884 (.A1(b[27]), .A2(a[10]), .B1(b[26]), .B2(a[11]), .ZN(n_1245));
   NAND2_X1 i_885 (.A1(b[28]), .A2(a[9]), .ZN(n_1246));
   OAI21_X1 i_886 (.A(n_1244), .B1(n_1245), .B2(n_1246), .ZN(n_3433));
   NAND4_X1 i_887 (.A1(b[24]), .A2(b[23]), .A3(a[14]), .A4(a[13]), .ZN(n_1248));
   AOI22_X1 i_888 (.A1(b[24]), .A2(a[13]), .B1(b[23]), .B2(a[14]), .ZN(n_1249));
   NAND2_X1 i_889 (.A1(b[25]), .A2(a[12]), .ZN(n_1250));
   OAI21_X1 i_890 (.A(n_1248), .B1(n_1249), .B2(n_1250), .ZN(n_3440));
   NAND4_X1 i_891 (.A1(b[21]), .A2(b[20]), .A3(a[17]), .A4(a[16]), .ZN(n_1251));
   AOI22_X1 i_892 (.A1(b[21]), .A2(a[16]), .B1(b[20]), .B2(a[17]), .ZN(n_1252));
   NAND2_X1 i_893 (.A1(b[22]), .A2(a[15]), .ZN(n_1253));
   OAI21_X1 i_894 (.A(n_1251), .B1(n_1252), .B2(n_1253), .ZN(n_3447));
   NAND4_X1 i_895 (.A1(a[20]), .A2(a[19]), .A3(b[18]), .A4(b[17]), .ZN(n_1255));
   AOI22_X1 i_896 (.A1(a[19]), .A2(b[18]), .B1(a[20]), .B2(b[17]), .ZN(n_1256));
   NAND2_X1 i_897 (.A1(b[19]), .A2(a[18]), .ZN(n_1257));
   OAI21_X1 i_898 (.A(n_1255), .B1(n_1256), .B2(n_1257), .ZN(n_3454));
   NAND4_X1 i_899 (.A1(a[23]), .A2(a[22]), .A3(b[15]), .A4(b[14]), .ZN(n_1258));
   AOI22_X1 i_900 (.A1(a[22]), .A2(b[15]), .B1(a[23]), .B2(b[14]), .ZN(n_1271));
   NAND2_X1 i_901 (.A1(a[21]), .A2(b[16]), .ZN(n_1272));
   OAI21_X1 i_902 (.A(n_1258), .B1(n_1271), .B2(n_1272), .ZN(n_3461));
   INV_X1 i_903 (.A(n_1242), .ZN(n_1275));
   NAND2_X1 i_904 (.A1(n_1275), .A2(n_1239), .ZN(n_1276));
   XOR2_X1 i_905 (.A(n_1276), .B(n_1243), .Z(n_3425));
   INV_X1 i_906 (.A(n_1245), .ZN(n_1277));
   NAND2_X1 i_907 (.A1(n_1277), .A2(n_1244), .ZN(n_1278));
   XOR2_X1 i_908 (.A(n_1278), .B(n_1246), .Z(n_3432));
   INV_X1 i_909 (.A(n_1249), .ZN(n_1279));
   NAND2_X1 i_910 (.A1(n_1279), .A2(n_1248), .ZN(n_1282));
   XOR2_X1 i_911 (.A(n_1282), .B(n_1250), .Z(n_3439));
   INV_X1 i_912 (.A(n_1252), .ZN(n_1283));
   NAND2_X1 i_913 (.A1(n_1283), .A2(n_1251), .ZN(n_1284));
   XOR2_X1 i_914 (.A(n_1284), .B(n_1253), .Z(n_3446));
   INV_X1 i_915 (.A(n_1256), .ZN(n_1285));
   NAND2_X1 i_916 (.A1(n_1285), .A2(n_1255), .ZN(n_1286));
   XOR2_X1 i_917 (.A(n_1286), .B(n_1257), .Z(n_3453));
   INV_X1 i_918 (.A(n_1271), .ZN(n_1289));
   NAND2_X1 i_919 (.A1(n_1289), .A2(n_1258), .ZN(n_1290));
   XOR2_X1 i_920 (.A(n_1290), .B(n_1272), .Z(n_3460));
   INV_X1 i_921 (.A(n_1137), .ZN(n_1291));
   NAND2_X1 i_922 (.A1(n_1291), .A2(n_1136), .ZN(n_1292));
   XOR2_X1 i_923 (.A(n_1292), .B(n_1138), .Z(n_3467));
   INV_X1 i_924 (.A(n_1132), .ZN(n_1293));
   NAND2_X1 i_925 (.A1(n_1131), .A2(n_1293), .ZN(n_1295));
   XOR2_X1 i_926 (.A(n_1295), .B(n_1133), .Z(n_3474));
   INV_X1 i_927 (.A(n_1237), .ZN(n_1296));
   NAND2_X1 i_928 (.A1(n_1236), .A2(n_1296), .ZN(n_1297));
   XOR2_X1 i_929 (.A(n_1297), .B(n_1238), .Z(n_3480));
   NAND4_X1 i_930 (.A1(b[30]), .A2(b[29]), .A3(a[7]), .A4(a[6]), .ZN(n_1298));
   AOI22_X1 i_931 (.A1(b[30]), .A2(a[6]), .B1(b[29]), .B2(a[7]), .ZN(n_1299));
   NAND2_X1 i_932 (.A1(b[31]), .A2(a[5]), .ZN(n_1300));
   OAI21_X1 i_933 (.A(n_1298), .B1(n_1299), .B2(n_1300), .ZN(n_3329));
   NAND4_X1 i_934 (.A1(b[27]), .A2(b[26]), .A3(a[10]), .A4(a[9]), .ZN(n_1303));
   AOI22_X1 i_935 (.A1(b[27]), .A2(a[9]), .B1(b[26]), .B2(a[10]), .ZN(n_1304));
   NAND2_X1 i_936 (.A1(b[28]), .A2(a[8]), .ZN(n_1305));
   OAI21_X1 i_937 (.A(n_1303), .B1(n_1304), .B2(n_1305), .ZN(n_3336));
   NAND4_X1 i_938 (.A1(b[24]), .A2(b[23]), .A3(a[13]), .A4(a[12]), .ZN(n_1306));
   AOI22_X1 i_939 (.A1(b[24]), .A2(a[12]), .B1(b[23]), .B2(a[13]), .ZN(n_1319));
   NAND2_X1 i_940 (.A1(b[25]), .A2(a[11]), .ZN(n_1320));
   OAI21_X1 i_941 (.A(n_1306), .B1(n_1319), .B2(n_1320), .ZN(n_3343));
   NAND4_X1 i_942 (.A1(b[21]), .A2(b[20]), .A3(a[16]), .A4(a[15]), .ZN(n_1323));
   AOI22_X1 i_943 (.A1(b[21]), .A2(a[15]), .B1(b[20]), .B2(a[16]), .ZN(n_1324));
   NAND2_X1 i_944 (.A1(b[22]), .A2(a[14]), .ZN(n_1325));
   OAI21_X1 i_945 (.A(n_1323), .B1(n_1324), .B2(n_1325), .ZN(n_3350));
   NAND4_X1 i_946 (.A1(a[19]), .A2(a[18]), .A3(b[18]), .A4(b[17]), .ZN(n_1326));
   AOI22_X1 i_947 (.A1(a[18]), .A2(b[18]), .B1(a[19]), .B2(b[17]), .ZN(n_1327));
   NAND2_X1 i_948 (.A1(b[19]), .A2(a[17]), .ZN(n_1330));
   OAI21_X1 i_949 (.A(n_1326), .B1(n_1327), .B2(n_1330), .ZN(n_3357));
   NAND4_X1 i_950 (.A1(a[22]), .A2(a[21]), .A3(b[15]), .A4(b[14]), .ZN(n_1331));
   AOI22_X1 i_951 (.A1(a[21]), .A2(b[15]), .B1(a[22]), .B2(b[14]), .ZN(n_1332));
   NAND2_X1 i_952 (.A1(a[20]), .A2(b[16]), .ZN(n_1333));
   OAI21_X1 i_953 (.A(n_1331), .B1(n_1332), .B2(n_1333), .ZN(n_3364));
   NAND4_X1 i_954 (.A1(a[25]), .A2(a[24]), .A3(b[12]), .A4(b[11]), .ZN(n_1334));
   AOI22_X1 i_955 (.A1(a[24]), .A2(b[12]), .B1(a[25]), .B2(b[11]), .ZN(n_1337));
   NAND2_X1 i_956 (.A1(a[23]), .A2(b[13]), .ZN(n_1338));
   OAI21_X1 i_957 (.A(n_1334), .B1(n_1337), .B2(n_1338), .ZN(n_3371));
   NAND4_X1 i_958 (.A1(a[28]), .A2(a[27]), .A3(b[9]), .A4(b[8]), .ZN(n_1339));
   AOI22_X1 i_959 (.A1(a[27]), .A2(b[9]), .B1(a[28]), .B2(b[8]), .ZN(n_1340));
   NAND2_X1 i_960 (.A1(a[26]), .A2(b[10]), .ZN(n_1341));
   OAI21_X1 i_961 (.A(n_1339), .B1(n_1340), .B2(n_1341), .ZN(n_3378));
   INV_X1 i_962 (.A(n_1299), .ZN(n_1344));
   NAND2_X1 i_963 (.A1(n_1344), .A2(n_1298), .ZN(n_1345));
   XOR2_X1 i_964 (.A(n_1345), .B(n_1300), .Z(n_3328));
   INV_X1 i_965 (.A(n_1304), .ZN(n_1346));
   NAND2_X1 i_966 (.A1(n_1346), .A2(n_1303), .ZN(n_1347));
   XOR2_X1 i_967 (.A(n_1347), .B(n_1305), .Z(n_3335));
   INV_X1 i_968 (.A(n_1319), .ZN(n_1350));
   NAND2_X1 i_969 (.A1(n_1350), .A2(n_1306), .ZN(n_1351));
   XOR2_X1 i_970 (.A(n_1351), .B(n_1320), .Z(n_3342));
   INV_X1 i_971 (.A(n_1324), .ZN(n_1352));
   NAND2_X1 i_972 (.A1(n_1352), .A2(n_1323), .ZN(n_1353));
   XOR2_X1 i_973 (.A(n_1353), .B(n_1325), .Z(n_3349));
   INV_X1 i_974 (.A(n_1327), .ZN(n_1354));
   NAND2_X1 i_975 (.A1(n_1354), .A2(n_1326), .ZN(n_1369));
   XOR2_X1 i_976 (.A(n_1369), .B(n_1330), .Z(n_3356));
   INV_X1 i_977 (.A(n_1332), .ZN(n_1370));
   NAND2_X1 i_978 (.A1(n_1370), .A2(n_1331), .ZN(n_1373));
   XOR2_X1 i_979 (.A(n_1373), .B(n_1333), .Z(n_3363));
   INV_X1 i_980 (.A(n_1337), .ZN(n_1374));
   NAND2_X1 i_981 (.A1(n_1374), .A2(n_1334), .ZN(n_1375));
   XOR2_X1 i_982 (.A(n_1375), .B(n_1338), .Z(n_3370));
   INV_X1 i_983 (.A(n_1340), .ZN(n_1376));
   NAND2_X1 i_984 (.A1(n_1376), .A2(n_1339), .ZN(n_1377));
   XOR2_X1 i_985 (.A(n_1377), .B(n_1341), .Z(n_3377));
   XNOR2_X1 i_986 (.A(n_1219), .B(n_1220), .ZN(n_1380));
   XOR2_X1 i_987 (.A(n_1380), .B(n_1218), .Z(n_3384));
   NAND4_X1 i_988 (.A1(a[26]), .A2(a[25]), .A3(b[9]), .A4(b[8]), .ZN(n_1381));
   AOI22_X1 i_989 (.A1(a[25]), .A2(b[9]), .B1(a[26]), .B2(b[8]), .ZN(n_1382));
   NAND2_X1 i_990 (.A1(a[24]), .A2(b[10]), .ZN(n_1383));
   OAI21_X1 i_991 (.A(n_1381), .B1(n_1382), .B2(n_1383), .ZN(n_1384));
   NAND4_X1 i_992 (.A1(a[29]), .A2(a[28]), .A3(b[6]), .A4(b[5]), .ZN(n_1387));
   AOI22_X1 i_993 (.A1(a[28]), .A2(b[6]), .B1(a[29]), .B2(b[5]), .ZN(n_1388));
   NAND2_X1 i_994 (.A1(a[27]), .A2(b[7]), .ZN(n_1389));
   OAI21_X1 i_995 (.A(n_1387), .B1(n_1388), .B2(n_1389), .ZN(n_1390));
   NOR2_X1 i_996 (.A1(n_1384), .A2(n_1390), .ZN(n_1391));
   NAND2_X1 i_997 (.A1(a[31]), .A2(b[4]), .ZN(n_1393));
   NAND2_X1 i_998 (.A1(n_1384), .A2(n_1390), .ZN(n_1394));
   AOI21_X1 i_999 (.A(n_1391), .B1(n_1393), .B2(n_1394), .ZN(n_3287));
   NAND4_X1 i_1000 (.A1(b[30]), .A2(b[29]), .A3(a[5]), .A4(a[6]), .ZN(n_1395));
   AOI22_X1 i_1001 (.A1(b[30]), .A2(a[5]), .B1(b[29]), .B2(a[6]), .ZN(n_1396));
   NAND2_X1 i_1002 (.A1(b[31]), .A2(a[4]), .ZN(n_1397));
   OAI21_X1 i_1003 (.A(n_1395), .B1(n_1396), .B2(n_1397), .ZN(n_3224));
   NAND4_X1 i_1004 (.A1(b[27]), .A2(b[26]), .A3(a[8]), .A4(a[9]), .ZN(n_1398));
   AOI22_X1 i_1005 (.A1(b[27]), .A2(a[8]), .B1(b[26]), .B2(a[9]), .ZN(n_1400));
   NAND2_X1 i_1006 (.A1(b[28]), .A2(a[7]), .ZN(n_1401));
   OAI21_X1 i_1007 (.A(n_1398), .B1(n_1400), .B2(n_1401), .ZN(n_3231));
   NAND4_X1 i_1008 (.A1(b[24]), .A2(b[23]), .A3(a[11]), .A4(a[12]), .ZN(n_1402));
   AOI22_X1 i_1009 (.A1(b[24]), .A2(a[11]), .B1(b[23]), .B2(a[12]), .ZN(n_1403));
   NAND2_X1 i_1010 (.A1(b[25]), .A2(a[10]), .ZN(n_1420));
   OAI21_X1 i_1011 (.A(n_1402), .B1(n_1403), .B2(n_1420), .ZN(n_3238));
   NAND4_X1 i_1012 (.A1(b[21]), .A2(b[20]), .A3(a[14]), .A4(a[15]), .ZN(n_1421));
   AOI22_X1 i_1013 (.A1(b[21]), .A2(a[14]), .B1(b[20]), .B2(a[15]), .ZN(n_1424));
   NAND2_X1 i_1014 (.A1(b[22]), .A2(a[13]), .ZN(n_1425));
   OAI21_X1 i_1015 (.A(n_1421), .B1(n_1424), .B2(n_1425), .ZN(n_3245));
   NAND4_X1 i_1016 (.A1(a[17]), .A2(a[18]), .A3(b[18]), .A4(b[17]), .ZN(n_1426));
   AOI22_X1 i_1017 (.A1(a[17]), .A2(b[18]), .B1(a[18]), .B2(b[17]), .ZN(n_1427));
   NAND2_X1 i_1018 (.A1(b[19]), .A2(a[16]), .ZN(n_1428));
   OAI21_X1 i_1019 (.A(n_1426), .B1(n_1427), .B2(n_1428), .ZN(n_3252));
   NAND4_X1 i_1020 (.A1(a[20]), .A2(a[21]), .A3(b[15]), .A4(b[14]), .ZN(n_1431));
   AOI22_X1 i_1021 (.A1(a[20]), .A2(b[15]), .B1(a[21]), .B2(b[14]), .ZN(n_1432));
   NAND2_X1 i_1022 (.A1(a[19]), .A2(b[16]), .ZN(n_1433));
   OAI21_X1 i_1023 (.A(n_1431), .B1(n_1432), .B2(n_1433), .ZN(n_3259));
   NAND4_X1 i_1024 (.A1(a[23]), .A2(a[24]), .A3(b[12]), .A4(b[11]), .ZN(n_1434));
   AOI22_X1 i_1025 (.A1(a[23]), .A2(b[12]), .B1(a[24]), .B2(b[11]), .ZN(n_1435));
   NAND2_X1 i_1026 (.A1(a[22]), .A2(b[13]), .ZN(n_1438));
   OAI21_X1 i_1027 (.A(n_1434), .B1(n_1435), .B2(n_1438), .ZN(n_3266));
   NAND4_X1 i_1028 (.A1(a[26]), .A2(a[27]), .A3(b[9]), .A4(b[8]), .ZN(n_1439));
   AOI22_X1 i_1029 (.A1(a[26]), .A2(b[9]), .B1(a[27]), .B2(b[8]), .ZN(n_1440));
   NAND2_X1 i_1030 (.A1(a[25]), .A2(b[10]), .ZN(n_1441));
   OAI21_X1 i_1031 (.A(n_1439), .B1(n_1440), .B2(n_1441), .ZN(n_3273));
   OR3_X1 i_1032 (.A1(n_1219), .A2(n_497), .A3(n_1232), .ZN(n_1442));
   AOI21_X1 i_1033 (.A(n_1235), .B1(a[29]), .B2(b[6]), .ZN(n_1445));
   NAND2_X1 i_1034 (.A1(a[28]), .A2(b[7]), .ZN(n_1446));
   OAI21_X1 i_1035 (.A(n_1442), .B1(n_1445), .B2(n_1446), .ZN(n_3280));
   INV_X1 i_1036 (.A(n_1391), .ZN(n_1447));
   NAND2_X1 i_1037 (.A1(n_1447), .A2(n_1394), .ZN(n_1448));
   XOR2_X1 i_1038 (.A(n_1448), .B(n_1393), .Z(n_3286));
   INV_X1 i_1039 (.A(n_1396), .ZN(n_1449));
   NAND2_X1 i_1040 (.A1(n_1449), .A2(n_1395), .ZN(n_1451));
   XOR2_X1 i_1041 (.A(n_1451), .B(n_1397), .Z(n_3223));
   INV_X1 i_1042 (.A(n_1400), .ZN(n_1452));
   NAND2_X1 i_1043 (.A1(n_1452), .A2(n_1398), .ZN(n_1453));
   XOR2_X1 i_1044 (.A(n_1453), .B(n_1401), .Z(n_3230));
   INV_X1 i_1045 (.A(n_1403), .ZN(n_1454));
   NAND2_X1 i_1046 (.A1(n_1454), .A2(n_1402), .ZN(n_1455));
   XOR2_X1 i_1047 (.A(n_1455), .B(n_1420), .Z(n_3237));
   INV_X1 i_1048 (.A(n_1424), .ZN(n_1456));
   NAND2_X1 i_1049 (.A1(n_1456), .A2(n_1421), .ZN(n_1459));
   XOR2_X1 i_1050 (.A(n_1459), .B(n_1425), .Z(n_3244));
   INV_X1 i_1051 (.A(n_1427), .ZN(n_1460));
   NAND2_X1 i_1053 (.A1(n_1460), .A2(n_1426), .ZN(n_1461));
   XOR2_X1 i_1054 (.A(n_1461), .B(n_1428), .Z(n_3251));
   INV_X1 i_1055 (.A(n_1432), .ZN(n_1462));
   NAND2_X1 i_1056 (.A1(n_1462), .A2(n_1431), .ZN(n_1479));
   XOR2_X1 i_1057 (.A(n_1479), .B(n_1433), .Z(n_3258));
   INV_X1 i_1058 (.A(n_1435), .ZN(n_1480));
   NAND2_X1 i_1059 (.A1(n_1480), .A2(n_1434), .ZN(n_1483));
   XOR2_X1 i_1060 (.A(n_1483), .B(n_1438), .Z(n_3265));
   INV_X1 i_1061 (.A(n_1440), .ZN(n_1484));
   NAND2_X1 i_1062 (.A1(n_1484), .A2(n_1439), .ZN(n_1485));
   XOR2_X1 i_1063 (.A(n_1485), .B(n_1441), .Z(n_3272));
   INV_X1 i_1064 (.A(n_1445), .ZN(n_1486));
   NAND2_X1 i_1065 (.A1(n_1442), .A2(n_1486), .ZN(n_1487));
   XOR2_X1 i_1066 (.A(n_1487), .B(n_1446), .Z(n_3279));
   NAND4_X1 i_1069 (.A1(b[30]), .A2(b[29]), .A3(a[5]), .A4(a[4]), .ZN(n_1490));
   AOI22_X1 i_1070 (.A1(b[30]), .A2(a[4]), .B1(b[29]), .B2(a[5]), .ZN(n_1491));
   NAND2_X1 i_1071 (.A1(b[31]), .A2(a[3]), .ZN(n_1492));
   OAI21_X1 i_1072 (.A(n_1490), .B1(n_1491), .B2(n_1492), .ZN(n_3117));
   NAND4_X1 i_1073 (.A1(b[27]), .A2(b[26]), .A3(a[8]), .A4(a[7]), .ZN(n_1493));
   AOI22_X1 i_1074 (.A1(b[27]), .A2(a[7]), .B1(b[26]), .B2(a[8]), .ZN(n_1494));
   NAND2_X1 i_1075 (.A1(b[28]), .A2(a[6]), .ZN(n_1497));
   OAI21_X1 i_1076 (.A(n_1493), .B1(n_1494), .B2(n_1497), .ZN(n_3124));
   NAND4_X1 i_1077 (.A1(b[24]), .A2(b[23]), .A3(a[11]), .A4(a[10]), .ZN(n_1498));
   AOI22_X1 i_1078 (.A1(b[24]), .A2(a[10]), .B1(b[23]), .B2(a[11]), .ZN(n_1499));
   NAND2_X1 i_1079 (.A1(b[25]), .A2(a[9]), .ZN(n_1500));
   OAI21_X1 i_1080 (.A(n_1498), .B1(n_1499), .B2(n_1500), .ZN(n_3131));
   NAND4_X1 i_1081 (.A1(b[21]), .A2(b[20]), .A3(a[14]), .A4(a[13]), .ZN(n_1501));
   AOI22_X1 i_1082 (.A1(b[21]), .A2(a[13]), .B1(b[20]), .B2(a[14]), .ZN(n_1504));
   NAND2_X1 i_1083 (.A1(b[22]), .A2(a[12]), .ZN(n_1505));
   OAI21_X1 i_1084 (.A(n_1501), .B1(n_1504), .B2(n_1505), .ZN(n_3138));
   NAND4_X1 i_1085 (.A1(a[17]), .A2(b[18]), .A3(b[17]), .A4(a[16]), .ZN(n_1506));
   AOI22_X1 i_1086 (.A1(b[18]), .A2(a[16]), .B1(a[17]), .B2(b[17]), .ZN(n_1507));
   NAND2_X1 i_1087 (.A1(b[19]), .A2(a[15]), .ZN(n_1508));
   OAI21_X1 i_1088 (.A(n_1506), .B1(n_1507), .B2(n_1508), .ZN(n_3145));
   NAND4_X1 i_1089 (.A1(a[20]), .A2(a[19]), .A3(b[15]), .A4(b[14]), .ZN(n_1511));
   AOI22_X1 i_1090 (.A1(a[19]), .A2(b[15]), .B1(a[20]), .B2(b[14]), .ZN(n_1512));
   NAND2_X1 i_1093 (.A1(a[18]), .A2(b[16]), .ZN(n_1513));
   OAI21_X1 i_1094 (.A(n_1511), .B1(n_1512), .B2(n_1513), .ZN(n_3152));
   NAND4_X1 i_1095 (.A1(a[23]), .A2(a[22]), .A3(b[12]), .A4(b[11]), .ZN(n_1514));
   AOI22_X1 i_1096 (.A1(a[22]), .A2(b[12]), .B1(a[23]), .B2(b[11]), .ZN(n_1517));
   NAND2_X1 i_1097 (.A1(a[21]), .A2(b[13]), .ZN(n_1518));
   OAI21_X1 i_1098 (.A(n_1514), .B1(n_1517), .B2(n_1518), .ZN(n_3159));
   INV_X1 i_1099 (.A(n_1491), .ZN(n_1519));
   NAND2_X1 i_1100 (.A1(n_1519), .A2(n_1490), .ZN(n_1520));
   XOR2_X1 i_1101 (.A(n_1520), .B(n_1492), .Z(n_3116));
   INV_X1 i_1102 (.A(n_1494), .ZN(n_1521));
   NAND2_X1 i_1103 (.A1(n_1521), .A2(n_1493), .ZN(n_1540));
   XOR2_X1 i_1104 (.A(n_1540), .B(n_1497), .Z(n_3123));
   INV_X1 i_1105 (.A(n_1499), .ZN(n_1541));
   NAND2_X1 i_1106 (.A1(n_1541), .A2(n_1498), .ZN(n_1544));
   XOR2_X1 i_1107 (.A(n_1544), .B(n_1500), .Z(n_3130));
   INV_X1 i_1108 (.A(n_1504), .ZN(n_1545));
   NAND2_X1 i_1109 (.A1(n_1545), .A2(n_1501), .ZN(n_1546));
   XOR2_X1 i_1110 (.A(n_1546), .B(n_1505), .Z(n_3137));
   INV_X1 i_1111 (.A(n_1507), .ZN(n_1547));
   NAND2_X1 i_1112 (.A1(n_1547), .A2(n_1506), .ZN(n_1548));
   XOR2_X1 i_1113 (.A(n_1548), .B(n_1508), .Z(n_3144));
   INV_X1 i_1114 (.A(n_1512), .ZN(n_1551));
   NAND2_X1 i_1118 (.A1(n_1551), .A2(n_1511), .ZN(n_1552));
   XOR2_X1 i_1119 (.A(n_1552), .B(n_1513), .Z(n_3151));
   INV_X1 i_1120 (.A(n_1517), .ZN(n_1553));
   NAND2_X1 i_1121 (.A1(n_1553), .A2(n_1514), .ZN(n_1554));
   XOR2_X1 i_1122 (.A(n_1554), .B(n_1518), .Z(n_3158));
   INV_X1 i_1123 (.A(n_1382), .ZN(n_1555));
   NAND2_X1 i_1124 (.A1(n_1555), .A2(n_1381), .ZN(n_1558));
   XOR2_X1 i_1125 (.A(n_1558), .B(n_1383), .Z(n_3165));
   INV_X1 i_1126 (.A(n_1388), .ZN(n_1559));
   NAND2_X1 i_1127 (.A1(n_1559), .A2(n_1387), .ZN(n_1560));
   XOR2_X1 i_1128 (.A(n_1560), .B(n_1389), .Z(n_3172));
   INV_X1 i_1129 (.A(b[4]), .ZN(n_1561));
   NAND2_X1 i_1130 (.A1(a[30]), .A2(b[3]), .ZN(n_1562));
   NAND2_X1 i_1131 (.A1(a[31]), .A2(b[2]), .ZN(n_1565));
   AOI211_X1 i_1132 (.A(n_497), .B(n_1561), .C1(n_1562), .C2(n_1565), .ZN(n_1566));
   INV_X1 i_1133 (.A(b[2]), .ZN(n_1567));
   NOR2_X1 i_1134 (.A1(n_659), .A2(n_1567), .ZN(n_1568));
   OAI211_X1 i_1135 (.A(a[31]), .B(b[3]), .C1(n_1566), .C2(n_1568), .ZN(n_1569));
   AOI21_X1 i_1136 (.A(n_1566), .B1(a[31]), .B2(b[3]), .ZN(n_1571));
   NAND2_X1 i_1137 (.A1(a[30]), .A2(b[4]), .ZN(n_1572));
   OAI21_X1 i_1138 (.A(n_1569), .B1(n_1571), .B2(n_1572), .ZN(n_3179));
   AND2_X1 i_1143 (.A1(n_1571), .A2(n_1572), .ZN(n_1573));
   OAI22_X1 i_1144 (.A1(n_1569), .A2(n_1572), .B1(n_3179), .B2(n_1573), .ZN(
      n_3178));
   NAND2_X1 i_1145 (.A1(b[30]), .A2(a[3]), .ZN(n_1574));
   INV_X1 i_1146 (.A(n_1574), .ZN(n_1575));
   NAND3_X1 i_1147 (.A1(n_1575), .A2(b[29]), .A3(a[4]), .ZN(n_1576));
   AOI21_X1 i_1148 (.A(n_1575), .B1(b[29]), .B2(a[4]), .ZN(n_1578));
   NAND2_X1 i_1149 (.A1(b[31]), .A2(a[2]), .ZN(n_1579));
   OAI21_X1 i_1150 (.A(n_1576), .B1(n_1578), .B2(n_1579), .ZN(n_3009));
   NAND2_X1 i_1151 (.A1(b[27]), .A2(a[6]), .ZN(n_1580));
   INV_X1 i_1152 (.A(n_1580), .ZN(n_1581));
   NAND3_X1 i_1153 (.A1(n_1581), .A2(b[26]), .A3(a[7]), .ZN(n_1602));
   AOI21_X1 i_1154 (.A(n_1581), .B1(b[26]), .B2(a[7]), .ZN(n_1603));
   NAND2_X1 i_1155 (.A1(b[28]), .A2(a[5]), .ZN(n_1606));
   OAI21_X1 i_1156 (.A(n_1602), .B1(n_1603), .B2(n_1606), .ZN(n_3016));
   NAND2_X1 i_1157 (.A1(b[24]), .A2(a[9]), .ZN(n_1607));
   INV_X1 i_1158 (.A(n_1607), .ZN(n_1608));
   NAND3_X1 i_1159 (.A1(n_1608), .A2(b[23]), .A3(a[10]), .ZN(n_1609));
   AOI21_X1 i_1160 (.A(n_1608), .B1(b[23]), .B2(a[10]), .ZN(n_1610));
   NAND2_X1 i_1161 (.A1(b[25]), .A2(a[8]), .ZN(n_1613));
   OAI21_X1 i_1162 (.A(n_1609), .B1(n_1610), .B2(n_1613), .ZN(n_3023));
   NAND2_X1 i_1163 (.A1(b[21]), .A2(a[12]), .ZN(n_1614));
   INV_X1 i_1164 (.A(n_1614), .ZN(n_1615));
   NAND3_X1 i_1165 (.A1(n_1615), .A2(b[20]), .A3(a[13]), .ZN(n_1616));
   AOI21_X1 i_1166 (.A(n_1615), .B1(b[20]), .B2(a[13]), .ZN(n_1617));
   NAND2_X1 i_1167 (.A1(b[22]), .A2(a[11]), .ZN(n_1620));
   OAI21_X1 i_1168 (.A(n_1616), .B1(n_1617), .B2(n_1620), .ZN(n_3030));
   NAND2_X1 i_1169 (.A1(b[18]), .A2(a[15]), .ZN(n_1621));
   INV_X1 i_1170 (.A(n_1621), .ZN(n_1622));
   NAND3_X1 i_1171 (.A1(n_1622), .A2(b[17]), .A3(a[16]), .ZN(n_1623));
   AOI21_X1 i_1176 (.A(n_1622), .B1(b[17]), .B2(a[16]), .ZN(n_1624));
   NAND2_X1 i_1177 (.A1(b[19]), .A2(a[14]), .ZN(n_1627));
   OAI21_X1 i_1178 (.A(n_1623), .B1(n_1624), .B2(n_1627), .ZN(n_3037));
   NAND2_X1 i_1179 (.A1(a[18]), .A2(b[15]), .ZN(n_1628));
   INV_X1 i_1180 (.A(n_1628), .ZN(n_1629));
   NAND3_X1 i_1181 (.A1(n_1629), .A2(a[19]), .A3(b[14]), .ZN(n_1630));
   AOI21_X1 i_1182 (.A(n_1629), .B1(a[19]), .B2(b[14]), .ZN(n_1631));
   NAND2_X1 i_1183 (.A1(a[17]), .A2(b[16]), .ZN(n_1634));
   OAI21_X1 i_1184 (.A(n_1630), .B1(n_1631), .B2(n_1634), .ZN(n_3044));
   NAND2_X1 i_1185 (.A1(a[21]), .A2(b[12]), .ZN(n_1635));
   INV_X1 i_1186 (.A(n_1635), .ZN(n_1636));
   NAND3_X1 i_1187 (.A1(n_1636), .A2(a[22]), .A3(b[11]), .ZN(n_1637));
   AOI21_X1 i_1188 (.A(n_1636), .B1(a[22]), .B2(b[11]), .ZN(n_1638));
   NAND2_X1 i_1189 (.A1(a[20]), .A2(b[13]), .ZN(n_1640));
   OAI21_X1 i_1190 (.A(n_1637), .B1(n_1638), .B2(n_1640), .ZN(n_3051));
   NAND2_X1 i_1191 (.A1(a[24]), .A2(b[9]), .ZN(n_1641));
   INV_X1 i_1192 (.A(n_1641), .ZN(n_1642));
   NAND3_X1 i_1193 (.A1(n_1642), .A2(a[25]), .A3(b[8]), .ZN(n_1643));
   AOI21_X1 i_1194 (.A(n_1642), .B1(a[25]), .B2(b[8]), .ZN(n_1644));
   NAND2_X1 i_1195 (.A1(a[23]), .A2(b[10]), .ZN(n_1645));
   OAI21_X1 i_1196 (.A(n_1643), .B1(n_1644), .B2(n_1645), .ZN(n_3058));
   NAND2_X1 i_1197 (.A1(a[27]), .A2(b[6]), .ZN(n_1648));
   INV_X1 i_1198 (.A(n_1648), .ZN(n_1649));
   NAND3_X1 i_1199 (.A1(n_1649), .A2(a[28]), .A3(b[5]), .ZN(n_1650));
   AOI21_X1 i_1200 (.A(n_1649), .B1(a[28]), .B2(b[5]), .ZN(n_1651));
   NAND2_X1 i_1201 (.A1(a[26]), .A2(b[7]), .ZN(n_1672));
   OAI21_X1 i_1202 (.A(n_1650), .B1(n_1651), .B2(n_1672), .ZN(n_3065));
   INV_X1 i_1203 (.A(n_1578), .ZN(n_1673));
   NAND2_X1 i_1204 (.A1(n_1576), .A2(n_1673), .ZN(n_1676));
   XOR2_X1 i_1210 (.A(n_1676), .B(n_1579), .Z(n_3008));
   INV_X1 i_1211 (.A(n_1603), .ZN(n_1677));
   NAND2_X1 i_1212 (.A1(n_1602), .A2(n_1677), .ZN(n_1678));
   XOR2_X1 i_1213 (.A(n_1678), .B(n_1606), .Z(n_3015));
   INV_X1 i_1214 (.A(n_1610), .ZN(n_1679));
   NAND2_X1 i_1215 (.A1(n_1609), .A2(n_1679), .ZN(n_1680));
   XOR2_X1 i_1216 (.A(n_1680), .B(n_1613), .Z(n_3022));
   INV_X1 i_1217 (.A(n_1617), .ZN(n_1683));
   NAND2_X1 i_1218 (.A1(n_1616), .A2(n_1683), .ZN(n_1684));
   XOR2_X1 i_1219 (.A(n_1684), .B(n_1620), .Z(n_3029));
   INV_X1 i_1220 (.A(n_1624), .ZN(n_1685));
   NAND2_X1 i_1221 (.A1(n_1623), .A2(n_1685), .ZN(n_1686));
   XOR2_X1 i_1222 (.A(n_1686), .B(n_1627), .Z(n_3036));
   INV_X1 i_1223 (.A(n_1631), .ZN(n_1687));
   NAND2_X1 i_1224 (.A1(n_1630), .A2(n_1687), .ZN(n_1690));
   XOR2_X1 i_1225 (.A(n_1690), .B(n_1634), .Z(n_3043));
   INV_X1 i_1226 (.A(n_1638), .ZN(n_1691));
   NAND2_X1 i_1227 (.A1(n_1637), .A2(n_1691), .ZN(n_1692));
   XOR2_X1 i_1228 (.A(n_1692), .B(n_1640), .Z(n_3050));
   INV_X1 i_1229 (.A(n_1644), .ZN(n_1693));
   NAND2_X1 i_1230 (.A1(n_1643), .A2(n_1693), .ZN(n_1694));
   XOR2_X1 i_1231 (.A(n_1694), .B(n_1645), .Z(n_3057));
   INV_X1 i_1232 (.A(n_1651), .ZN(n_1697));
   NAND2_X1 i_1233 (.A1(n_1650), .A2(n_1697), .ZN(n_1698));
   XOR2_X1 i_1234 (.A(n_1698), .B(n_1672), .Z(n_3064));
   XOR2_X1 i_1235 (.A(n_1562), .B(n_1565), .Z(n_1699));
   NAND2_X1 i_1236 (.A1(a[29]), .A2(b[4]), .ZN(n_1700));
   XNOR2_X1 i_1237 (.A(n_1699), .B(n_1700), .ZN(n_3071));
   NAND2_X1 i_1244 (.A1(a[26]), .A2(b[5]), .ZN(n_1701));
   INV_X1 i_1245 (.A(a[25]), .ZN(n_1704));
   INV_X1 i_1246 (.A(b[6]), .ZN(n_1705));
   OR3_X1 i_1247 (.A1(n_1701), .A2(n_1704), .A3(n_1705), .ZN(n_1706));
   INV_X1 i_1248 (.A(n_1706), .ZN(n_1707));
   AND2_X1 i_1249 (.A1(a[24]), .A2(b[7]), .ZN(n_1708));
   OAI21_X1 i_1250 (.A(n_1701), .B1(n_1704), .B2(n_1705), .ZN(n_1711));
   AOI21_X1 i_1251 (.A(n_1707), .B1(n_1708), .B2(n_1711), .ZN(n_1712));
   NAND2_X1 i_1252 (.A1(a[29]), .A2(b[2]), .ZN(n_1713));
   INV_X1 i_1253 (.A(b[3]), .ZN(n_1714));
   OR3_X1 i_1254 (.A1(n_1713), .A2(n_541), .A3(n_1714), .ZN(n_1717));
   INV_X1 i_1255 (.A(n_1717), .ZN(n_1718));
   INV_X1 i_1256 (.A(a[27]), .ZN(n_1719));
   NOR2_X1 i_1257 (.A1(n_1719), .A2(n_1561), .ZN(n_1720));
   OAI21_X1 i_1258 (.A(n_1713), .B1(n_541), .B2(n_1714), .ZN(n_1721));
   AOI21_X1 i_1259 (.A(n_1718), .B1(n_1720), .B2(n_1721), .ZN(n_1744));
   NAND2_X1 i_1260 (.A1(n_1712), .A2(n_1744), .ZN(n_1745));
   INV_X1 i_1261 (.A(n_1745), .ZN(n_1748));
   NAND2_X1 i_1262 (.A1(a[31]), .A2(b[1]), .ZN(n_1749));
   OR2_X1 i_1263 (.A1(n_1712), .A2(n_1744), .ZN(n_1750));
   AOI21_X1 i_1264 (.A(n_1748), .B1(n_1749), .B2(n_1750), .ZN(n_2963));
   NAND2_X1 i_1265 (.A1(b[29]), .A2(a[2]), .ZN(n_1751));
   NOR2_X1 i_1266 (.A1(n_1574), .A2(n_1751), .ZN(n_1752));
   INV_X1 i_1267 (.A(n_1752), .ZN(n_1755));
   AOI22_X1 i_1268 (.A1(b[30]), .A2(a[2]), .B1(b[29]), .B2(a[3]), .ZN(n_1756));
   NAND2_X1 i_1269 (.A1(b[31]), .A2(a[1]), .ZN(n_1757));
   OAI21_X1 i_1270 (.A(n_1755), .B1(n_1756), .B2(n_1757), .ZN(n_2893));
   NAND2_X1 i_1271 (.A1(b[26]), .A2(a[5]), .ZN(n_1758));
   NOR2_X1 i_1272 (.A1(n_1580), .A2(n_1758), .ZN(n_1759));
   INV_X1 i_1273 (.A(n_1759), .ZN(n_1762));
   AOI22_X1 i_1274 (.A1(b[27]), .A2(a[5]), .B1(b[26]), .B2(a[6]), .ZN(n_1763));
   NAND2_X1 i_1275 (.A1(b[28]), .A2(a[4]), .ZN(n_1764));
   OAI21_X1 i_1276 (.A(n_1762), .B1(n_1763), .B2(n_1764), .ZN(n_2900));
   NAND2_X1 i_1277 (.A1(b[23]), .A2(a[8]), .ZN(n_1765));
   NOR2_X1 i_1278 (.A1(n_1607), .A2(n_1765), .ZN(n_1766));
   INV_X1 i_1279 (.A(n_1766), .ZN(n_1769));
   AOI22_X1 i_1286 (.A1(b[24]), .A2(a[8]), .B1(b[23]), .B2(a[9]), .ZN(n_1770));
   NAND2_X1 i_1287 (.A1(b[25]), .A2(a[7]), .ZN(n_1771));
   OAI21_X1 i_1288 (.A(n_1769), .B1(n_1770), .B2(n_1771), .ZN(n_2907));
   NAND2_X1 i_1289 (.A1(b[20]), .A2(a[11]), .ZN(n_1772));
   NOR2_X1 i_1290 (.A1(n_1614), .A2(n_1772), .ZN(n_1773));
   INV_X1 i_1291 (.A(n_1773), .ZN(n_1776));
   AOI22_X1 i_1292 (.A1(b[21]), .A2(a[11]), .B1(b[20]), .B2(a[12]), .ZN(n_1777));
   NAND2_X1 i_1293 (.A1(b[22]), .A2(a[10]), .ZN(n_1778));
   OAI21_X1 i_1294 (.A(n_1776), .B1(n_1777), .B2(n_1778), .ZN(n_2914));
   NAND2_X1 i_1295 (.A1(b[17]), .A2(a[14]), .ZN(n_1779));
   NOR2_X1 i_1296 (.A1(n_1621), .A2(n_1779), .ZN(n_1780));
   INV_X1 i_1297 (.A(n_1780), .ZN(n_1782));
   AOI22_X1 i_1298 (.A1(b[18]), .A2(a[14]), .B1(b[17]), .B2(a[15]), .ZN(n_1783));
   NAND2_X1 i_1299 (.A1(b[19]), .A2(a[13]), .ZN(n_1784));
   OAI21_X1 i_1300 (.A(n_1782), .B1(n_1783), .B2(n_1784), .ZN(n_2921));
   NAND2_X1 i_1301 (.A1(a[17]), .A2(b[14]), .ZN(n_1785));
   NOR2_X1 i_1302 (.A1(n_1628), .A2(n_1785), .ZN(n_1786));
   INV_X1 i_1303 (.A(n_1786), .ZN(n_1787));
   AOI22_X1 i_1304 (.A1(a[17]), .A2(b[15]), .B1(a[18]), .B2(b[14]), .ZN(n_1789));
   NAND2_X1 i_1305 (.A1(a[16]), .A2(b[16]), .ZN(n_1790));
   OAI21_X1 i_1306 (.A(n_1787), .B1(n_1789), .B2(n_1790), .ZN(n_2928));
   NAND2_X1 i_1307 (.A1(a[20]), .A2(b[11]), .ZN(n_1791));
   NOR2_X1 i_1308 (.A1(n_1635), .A2(n_1791), .ZN(n_1792));
   INV_X1 i_1309 (.A(n_1792), .ZN(n_1817));
   AOI22_X1 i_1310 (.A1(a[20]), .A2(b[12]), .B1(a[21]), .B2(b[11]), .ZN(n_1818));
   NAND2_X1 i_1311 (.A1(a[19]), .A2(b[13]), .ZN(n_1821));
   OAI21_X1 i_1312 (.A(n_1817), .B1(n_1818), .B2(n_1821), .ZN(n_2935));
   NAND2_X1 i_1313 (.A1(a[23]), .A2(b[8]), .ZN(n_1822));
   NOR2_X1 i_1314 (.A1(n_1641), .A2(n_1822), .ZN(n_1823));
   INV_X1 i_1315 (.A(n_1823), .ZN(n_1824));
   AOI22_X1 i_1316 (.A1(a[23]), .A2(b[9]), .B1(a[24]), .B2(b[8]), .ZN(n_1825));
   NAND2_X1 i_1317 (.A1(a[22]), .A2(b[10]), .ZN(n_1828));
   OAI21_X1 i_1318 (.A(n_1824), .B1(n_1825), .B2(n_1828), .ZN(n_2942));
   NOR2_X1 i_1319 (.A1(n_1648), .A2(n_1701), .ZN(n_1829));
   INV_X1 i_1320 (.A(n_1829), .ZN(n_1830));
   AOI22_X1 i_1321 (.A1(a[26]), .A2(b[6]), .B1(a[27]), .B2(b[5]), .ZN(n_1831));
   NAND2_X1 i_1329 (.A1(a[25]), .A2(b[7]), .ZN(n_1832));
   OAI21_X1 i_1330 (.A(n_1830), .B1(n_1831), .B2(n_1832), .ZN(n_2949));
   OR2_X1 i_1331 (.A1(n_1562), .A2(n_1713), .ZN(n_1835));
   AOI21_X1 i_1332 (.A(n_1568), .B1(a[29]), .B2(b[3]), .ZN(n_1836));
   NAND2_X1 i_1333 (.A1(a[28]), .A2(b[4]), .ZN(n_1837));
   OAI21_X1 i_1334 (.A(n_1835), .B1(n_1836), .B2(n_1837), .ZN(n_2956));
   NAND2_X1 i_1335 (.A1(n_1750), .A2(n_1745), .ZN(n_1838));
   XOR2_X1 i_1336 (.A(n_1838), .B(n_1749), .Z(n_2962));
   NOR2_X1 i_1337 (.A1(n_1752), .A2(n_1756), .ZN(n_1839));
   XNOR2_X1 i_1338 (.A(n_1839), .B(n_1757), .ZN(n_2892));
   NOR2_X1 i_1339 (.A1(n_1759), .A2(n_1763), .ZN(n_1842));
   XNOR2_X1 i_1340 (.A(n_1842), .B(n_1764), .ZN(n_2899));
   NOR2_X1 i_1341 (.A1(n_1766), .A2(n_1770), .ZN(n_1843));
   XNOR2_X1 i_1342 (.A(n_1843), .B(n_1771), .ZN(n_2906));
   NOR2_X1 i_1343 (.A1(n_1773), .A2(n_1777), .ZN(n_1844));
   XNOR2_X1 i_1344 (.A(n_1844), .B(n_1778), .ZN(n_2913));
   NOR2_X1 i_1345 (.A1(n_1780), .A2(n_1783), .ZN(n_1845));
   XNOR2_X1 i_1346 (.A(n_1845), .B(n_1784), .ZN(n_2920));
   NOR2_X1 i_1347 (.A1(n_1786), .A2(n_1789), .ZN(n_1846));
   XNOR2_X1 i_1348 (.A(n_1846), .B(n_1790), .ZN(n_2927));
   NOR2_X1 i_1349 (.A1(n_1792), .A2(n_1818), .ZN(n_1849));
   XNOR2_X1 i_1350 (.A(n_1849), .B(n_1821), .ZN(n_2934));
   NOR2_X1 i_1351 (.A1(n_1823), .A2(n_1825), .ZN(n_1850));
   XNOR2_X1 i_1352 (.A(n_1850), .B(n_1828), .ZN(n_2941));
   NOR2_X1 i_1353 (.A1(n_1829), .A2(n_1831), .ZN(n_1851));
   XNOR2_X1 i_1354 (.A(n_1851), .B(n_1832), .ZN(n_2948));
   INV_X1 i_1355 (.A(n_1836), .ZN(n_1852));
   NAND2_X1 i_1356 (.A1(n_1835), .A2(n_1852), .ZN(n_1853));
   XOR2_X1 i_1357 (.A(n_1853), .B(n_1837), .Z(n_2955));
   NAND2_X1 i_1358 (.A1(a[28]), .A2(b[1]), .ZN(n_1856));
   NOR2_X1 i_1359 (.A1(n_1713), .A2(n_1856), .ZN(n_1857));
   INV_X1 i_1360 (.A(n_1857), .ZN(n_1858));
   AOI22_X1 i_1361 (.A1(a[29]), .A2(b[1]), .B1(a[28]), .B2(b[2]), .ZN(n_1859));
   NAND2_X1 i_1362 (.A1(a[27]), .A2(b[3]), .ZN(n_1860));
   OAI21_X1 i_1363 (.A(n_1858), .B1(n_1859), .B2(n_1860), .ZN(n_1862));
   AOI21_X1 i_1372 (.A(n_1862), .B1(a[31]), .B2(b[0]), .ZN(n_1863));
   NAND2_X1 i_1373 (.A1(a[30]), .A2(b[1]), .ZN(n_1864));
   NAND3_X1 i_1374 (.A1(n_1862), .A2(a[31]), .A3(b[0]), .ZN(n_1865));
   AOI21_X1 i_1375 (.A(n_1863), .B1(n_1864), .B2(n_1865), .ZN(n_2846));
   INV_X1 i_1376 (.A(n_1751), .ZN(n_1866));
   NAND3_X1 i_1377 (.A1(n_1866), .A2(b[30]), .A3(a[1]), .ZN(n_1867));
   AOI21_X1 i_1378 (.A(n_1866), .B1(b[30]), .B2(a[1]), .ZN(n_1870));
   NAND2_X1 i_1379 (.A1(b[31]), .A2(a[0]), .ZN(n_1871));
   OAI21_X1 i_1380 (.A(n_1867), .B1(n_1870), .B2(n_1871), .ZN(n_2777));
   INV_X1 i_1381 (.A(n_1758), .ZN(n_1872));
   NAND3_X1 i_1382 (.A1(n_1872), .A2(b[27]), .A3(a[4]), .ZN(n_1873));
   AOI21_X1 i_1383 (.A(n_1872), .B1(b[27]), .B2(a[4]), .ZN(n_1898));
   NAND2_X1 i_1384 (.A1(b[28]), .A2(a[3]), .ZN(n_1899));
   OAI21_X1 i_1385 (.A(n_1873), .B1(n_1898), .B2(n_1899), .ZN(n_2784));
   INV_X1 i_1386 (.A(n_1765), .ZN(n_1902));
   NAND3_X1 i_1387 (.A1(n_1902), .A2(b[24]), .A3(a[7]), .ZN(n_1903));
   AOI21_X1 i_1388 (.A(n_1902), .B1(b[24]), .B2(a[7]), .ZN(n_1904));
   NAND2_X1 i_1389 (.A1(b[25]), .A2(a[6]), .ZN(n_1905));
   OAI21_X1 i_1390 (.A(n_1903), .B1(n_1904), .B2(n_1905), .ZN(n_2791));
   INV_X1 i_1391 (.A(n_1772), .ZN(n_1906));
   NAND3_X1 i_1392 (.A1(n_1906), .A2(b[21]), .A3(a[10]), .ZN(n_1909));
   AOI21_X1 i_1393 (.A(n_1906), .B1(b[21]), .B2(a[10]), .ZN(n_1910));
   NAND2_X1 i_1394 (.A1(b[22]), .A2(a[9]), .ZN(n_1911));
   OAI21_X1 i_1395 (.A(n_1909), .B1(n_1910), .B2(n_1911), .ZN(n_2798));
   INV_X1 i_1396 (.A(n_1779), .ZN(n_1912));
   NAND3_X1 i_1397 (.A1(n_1912), .A2(b[18]), .A3(a[13]), .ZN(n_1913));
   AOI21_X1 i_1398 (.A(n_1912), .B1(b[18]), .B2(a[13]), .ZN(n_1916));
   NAND2_X1 i_1399 (.A1(b[19]), .A2(a[12]), .ZN(n_1917));
   OAI21_X1 i_1400 (.A(n_1913), .B1(n_1916), .B2(n_1917), .ZN(n_2805));
   INV_X1 i_1401 (.A(n_1785), .ZN(n_1918));
   NAND3_X1 i_1402 (.A1(n_1918), .A2(a[16]), .A3(b[15]), .ZN(n_1919));
   AOI21_X1 i_1403 (.A(n_1918), .B1(a[16]), .B2(b[15]), .ZN(n_1920));
   NAND2_X1 i_1404 (.A1(b[16]), .A2(a[15]), .ZN(n_1923));
   OAI21_X1 i_1405 (.A(n_1919), .B1(n_1920), .B2(n_1923), .ZN(n_2812));
   INV_X1 i_1406 (.A(n_1791), .ZN(n_1924));
   NAND3_X1 i_1407 (.A1(n_1924), .A2(a[19]), .A3(b[12]), .ZN(n_1925));
   AOI21_X1 i_1408 (.A(n_1924), .B1(a[19]), .B2(b[12]), .ZN(n_1926));
   NAND2_X1 i_1409 (.A1(a[18]), .A2(b[13]), .ZN(n_1927));
   OAI21_X1 i_1410 (.A(n_1925), .B1(n_1926), .B2(n_1927), .ZN(n_2819));
   INV_X1 i_1411 (.A(n_1822), .ZN(n_1930));
   NAND3_X1 i_1412 (.A1(n_1930), .A2(a[22]), .A3(b[9]), .ZN(n_1931));
   AOI21_X1 i_1413 (.A(n_1930), .B1(a[22]), .B2(b[9]), .ZN(n_1932));
   NAND2_X1 i_1414 (.A1(a[21]), .A2(b[10]), .ZN(n_1933));
   OAI21_X1 i_1423 (.A(n_1931), .B1(n_1932), .B2(n_1933), .ZN(n_2826));
   INV_X1 i_1424 (.A(n_1870), .ZN(n_1934));
   NAND2_X1 i_1425 (.A1(n_1867), .A2(n_1934), .ZN(n_1937));
   XOR2_X1 i_1426 (.A(n_1937), .B(n_1871), .Z(n_2776));
   INV_X1 i_1427 (.A(n_1898), .ZN(n_1938));
   NAND2_X1 i_1428 (.A1(n_1873), .A2(n_1938), .ZN(n_1939));
   XOR2_X1 i_1429 (.A(n_1939), .B(n_1899), .Z(n_2783));
   INV_X1 i_1430 (.A(n_1904), .ZN(n_1940));
   NAND2_X1 i_1431 (.A1(n_1903), .A2(n_1940), .ZN(n_1941));
   XOR2_X1 i_1432 (.A(n_1941), .B(n_1905), .Z(n_2790));
   INV_X1 i_1433 (.A(n_1910), .ZN(n_1944));
   NAND2_X1 i_1434 (.A1(n_1909), .A2(n_1944), .ZN(n_1945));
   XOR2_X1 i_1435 (.A(n_1945), .B(n_1911), .Z(n_2797));
   INV_X1 i_1436 (.A(n_1916), .ZN(n_1946));
   NAND2_X1 i_1437 (.A1(n_1913), .A2(n_1946), .ZN(n_1947));
   XOR2_X1 i_1438 (.A(n_1947), .B(n_1917), .Z(n_2804));
   INV_X1 i_1439 (.A(n_1920), .ZN(n_1950));
   NAND2_X1 i_1440 (.A1(n_1919), .A2(n_1950), .ZN(n_1951));
   XOR2_X1 i_1441 (.A(n_1951), .B(n_1923), .Z(n_2811));
   INV_X1 i_1442 (.A(n_1926), .ZN(n_1952));
   NAND2_X1 i_1443 (.A1(n_1925), .A2(n_1952), .ZN(n_1953));
   XOR2_X1 i_1444 (.A(n_1953), .B(n_1927), .Z(n_2818));
   INV_X1 i_1445 (.A(n_1932), .ZN(n_1954));
   NAND2_X1 i_1446 (.A1(n_1931), .A2(n_1954), .ZN(n_1981));
   XOR2_X1 i_1447 (.A(n_1981), .B(n_1933), .Z(n_2825));
   NAND2_X1 i_1448 (.A1(n_1706), .A2(n_1711), .ZN(n_1982));
   XNOR2_X1 i_1449 (.A(n_1982), .B(n_1708), .ZN(n_2832));
   NAND2_X1 i_1450 (.A1(n_1717), .A2(n_1721), .ZN(n_1985));
   XNOR2_X1 i_1451 (.A(n_1985), .B(n_1720), .ZN(n_2839));
   INV_X1 i_1452 (.A(n_1863), .ZN(n_1986));
   NAND2_X1 i_1453 (.A1(n_1986), .A2(n_1865), .ZN(n_1987));
   XOR2_X1 i_1454 (.A(n_1987), .B(n_1864), .Z(n_2845));
   NAND2_X1 i_1455 (.A1(a[25]), .A2(b[4]), .ZN(n_1988));
   INV_X1 i_1456 (.A(a[26]), .ZN(n_1989));
   OR3_X1 i_1457 (.A1(n_1988), .A2(n_1989), .A3(n_1714), .ZN(n_1992));
   INV_X1 i_1458 (.A(n_1992), .ZN(n_1993));
   AND2_X1 i_1459 (.A1(a[24]), .A2(b[5]), .ZN(n_1994));
   OAI21_X1 i_1460 (.A(n_1988), .B1(n_1989), .B2(n_1714), .ZN(n_1995));
   AOI21_X1 i_1461 (.A(n_1993), .B1(n_1994), .B2(n_1995), .ZN(n_1996));
   OR3_X1 i_1462 (.A1(n_1856), .A2(n_497), .A3(n_514), .ZN(n_1999));
   INV_X1 i_1463 (.A(n_1999), .ZN(n_2000));
   NOR2_X1 i_1464 (.A1(n_1719), .A2(n_1567), .ZN(n_2001));
   OAI21_X1 i_1465 (.A(n_1856), .B1(n_497), .B2(n_514), .ZN(n_2002));
   AOI21_X1 i_1475 (.A(n_2000), .B1(n_2001), .B2(n_2002), .ZN(n_2003));
   NAND2_X1 i_1476 (.A1(n_1996), .A2(n_2003), .ZN(n_2006));
   INV_X1 i_1477 (.A(n_2006), .ZN(n_2007));
   NAND2_X1 i_1478 (.A1(a[30]), .A2(b[0]), .ZN(n_2008));
   OR2_X1 i_1479 (.A1(n_1996), .A2(n_2003), .ZN(n_2009));
   AOI21_X1 i_1480 (.A(n_2007), .B1(n_2008), .B2(n_2009), .ZN(n_2733));
   NAND2_X1 i_1481 (.A1(b[28]), .A2(a[1]), .ZN(n_2010));
   NOR2_X1 i_1482 (.A1(n_1751), .A2(n_2010), .ZN(n_2013));
   INV_X1 i_1483 (.A(n_2013), .ZN(n_2014));
   AOI22_X1 i_1484 (.A1(b[28]), .A2(a[2]), .B1(b[29]), .B2(a[1]), .ZN(n_2015));
   NAND2_X1 i_1485 (.A1(b[30]), .A2(a[0]), .ZN(n_2016));
   OAI21_X1 i_1486 (.A(n_2014), .B1(n_2015), .B2(n_2016), .ZN(n_2663));
   NAND2_X1 i_1487 (.A1(b[25]), .A2(a[4]), .ZN(n_2017));
   NOR2_X1 i_1488 (.A1(n_1758), .A2(n_2017), .ZN(n_2020));
   INV_X1 i_1489 (.A(n_2020), .ZN(n_2021));
   AOI22_X1 i_1490 (.A1(b[25]), .A2(a[5]), .B1(b[26]), .B2(a[4]), .ZN(n_2022));
   NAND2_X1 i_1491 (.A1(b[27]), .A2(a[3]), .ZN(n_2023));
   OAI21_X1 i_1492 (.A(n_2021), .B1(n_2022), .B2(n_2023), .ZN(n_2670));
   NAND2_X1 i_1493 (.A1(b[22]), .A2(a[7]), .ZN(n_2024));
   NOR2_X1 i_1494 (.A1(n_1765), .A2(n_2024), .ZN(n_2026));
   INV_X1 i_1495 (.A(n_2026), .ZN(n_2027));
   AOI22_X1 i_1496 (.A1(b[22]), .A2(a[8]), .B1(b[23]), .B2(a[7]), .ZN(n_2028));
   NAND2_X1 i_1497 (.A1(b[24]), .A2(a[6]), .ZN(n_2029));
   OAI21_X1 i_1498 (.A(n_2027), .B1(n_2028), .B2(n_2029), .ZN(n_2677));
   NAND2_X1 i_1499 (.A1(b[19]), .A2(a[10]), .ZN(n_2030));
   NOR2_X1 i_1500 (.A1(n_1772), .A2(n_2030), .ZN(n_2031));
   INV_X1 i_1501 (.A(n_2031), .ZN(n_2033));
   AOI22_X1 i_1502 (.A1(b[19]), .A2(a[11]), .B1(b[20]), .B2(a[10]), .ZN(n_2034));
   NAND2_X1 i_1503 (.A1(b[21]), .A2(a[9]), .ZN(n_2035));
   OAI21_X1 i_1504 (.A(n_2033), .B1(n_2034), .B2(n_2035), .ZN(n_2684));
   NAND2_X1 i_1505 (.A1(b[16]), .A2(a[13]), .ZN(n_2036));
   NOR2_X1 i_1506 (.A1(n_1779), .A2(n_2036), .ZN(n_2065));
   INV_X1 i_1507 (.A(n_2065), .ZN(n_2066));
   AOI22_X1 i_1508 (.A1(b[16]), .A2(a[14]), .B1(b[17]), .B2(a[13]), .ZN(n_2069));
   NAND2_X1 i_1509 (.A1(b[18]), .A2(a[12]), .ZN(n_2070));
   OAI21_X1 i_1510 (.A(n_2066), .B1(n_2069), .B2(n_2070), .ZN(n_2691));
   NAND2_X1 i_1511 (.A1(a[16]), .A2(b[13]), .ZN(n_2071));
   NOR2_X1 i_1512 (.A1(n_1785), .A2(n_2071), .ZN(n_2072));
   INV_X1 i_1513 (.A(n_2072), .ZN(n_2073));
   AOI22_X1 i_1514 (.A1(a[17]), .A2(b[13]), .B1(a[16]), .B2(b[14]), .ZN(n_2076));
   NAND2_X1 i_1515 (.A1(a[15]), .A2(b[15]), .ZN(n_2077));
   OAI21_X1 i_1516 (.A(n_2073), .B1(n_2076), .B2(n_2077), .ZN(n_2698));
   NAND2_X1 i_1527 (.A1(a[19]), .A2(b[10]), .ZN(n_2078));
   NOR2_X1 i_1528 (.A1(n_1791), .A2(n_2078), .ZN(n_2079));
   INV_X1 i_1529 (.A(n_2079), .ZN(n_2080));
   AOI22_X1 i_1530 (.A1(a[20]), .A2(b[10]), .B1(a[19]), .B2(b[11]), .ZN(n_2083));
   NAND2_X1 i_1531 (.A1(a[18]), .A2(b[12]), .ZN(n_2084));
   OAI21_X1 i_1532 (.A(n_2080), .B1(n_2083), .B2(n_2084), .ZN(n_2705));
   NAND2_X1 i_1533 (.A1(a[22]), .A2(b[7]), .ZN(n_2085));
   NOR2_X1 i_1534 (.A1(n_1822), .A2(n_2085), .ZN(n_2086));
   INV_X1 i_1535 (.A(n_2086), .ZN(n_2087));
   AOI22_X1 i_1536 (.A1(a[23]), .A2(b[7]), .B1(a[22]), .B2(b[8]), .ZN(n_2090));
   NAND2_X1 i_1537 (.A1(a[21]), .A2(b[9]), .ZN(n_2091));
   OAI21_X1 i_1538 (.A(n_2087), .B1(n_2090), .B2(n_2091), .ZN(n_2712));
   NOR2_X1 i_1539 (.A1(n_1701), .A2(n_1988), .ZN(n_2092));
   INV_X1 i_1540 (.A(n_2092), .ZN(n_2093));
   AOI22_X1 i_1541 (.A1(a[26]), .A2(b[4]), .B1(a[25]), .B2(b[5]), .ZN(n_2094));
   NAND2_X1 i_1542 (.A1(a[24]), .A2(b[6]), .ZN(n_2097));
   OAI21_X1 i_1543 (.A(n_2093), .B1(n_2094), .B2(n_2097), .ZN(n_2719));
   NAND2_X1 i_1544 (.A1(n_2009), .A2(n_2006), .ZN(n_2098));
   XOR2_X1 i_1545 (.A(n_2098), .B(n_2008), .Z(n_2732));
   NOR2_X1 i_1546 (.A1(n_2013), .A2(n_2015), .ZN(n_2099));
   XNOR2_X1 i_1547 (.A(n_2099), .B(n_2016), .ZN(n_2662));
   NOR2_X1 i_1548 (.A1(n_2020), .A2(n_2022), .ZN(n_2100));
   XNOR2_X1 i_1549 (.A(n_2100), .B(n_2023), .ZN(n_2669));
   NOR2_X1 i_1550 (.A1(n_2026), .A2(n_2028), .ZN(n_2101));
   XNOR2_X1 i_1551 (.A(n_2101), .B(n_2029), .ZN(n_2676));
   NOR2_X1 i_1552 (.A1(n_2031), .A2(n_2034), .ZN(n_2104));
   XNOR2_X1 i_1553 (.A(n_2104), .B(n_2035), .ZN(n_2683));
   NOR2_X1 i_1554 (.A1(n_2065), .A2(n_2069), .ZN(n_2105));
   XNOR2_X1 i_1555 (.A(n_2105), .B(n_2070), .ZN(n_2690));
   NOR2_X1 i_1556 (.A1(n_2072), .A2(n_2076), .ZN(n_2106));
   XNOR2_X1 i_1557 (.A(n_2106), .B(n_2077), .ZN(n_2697));
   NOR2_X1 i_1558 (.A1(n_2079), .A2(n_2083), .ZN(n_2107));
   XNOR2_X1 i_1559 (.A(n_2107), .B(n_2084), .ZN(n_2704));
   NOR2_X1 i_1560 (.A1(n_2086), .A2(n_2090), .ZN(n_2108));
   XNOR2_X1 i_1561 (.A(n_2108), .B(n_2091), .ZN(n_2711));
   NOR2_X1 i_1562 (.A1(n_2092), .A2(n_2094), .ZN(n_2111));
   XNOR2_X1 i_1563 (.A(n_2111), .B(n_2097), .ZN(n_2718));
   NOR2_X1 i_1564 (.A1(n_1857), .A2(n_1859), .ZN(n_2112));
   XNOR2_X1 i_1565 (.A(n_2112), .B(n_1860), .ZN(n_2725));
   INV_X1 i_1566 (.A(n_2010), .ZN(n_2113));
   NAND3_X1 i_1567 (.A1(n_2113), .A2(b[27]), .A3(a[2]), .ZN(n_2114));
   AOI21_X1 i_1568 (.A(n_2113), .B1(b[27]), .B2(a[2]), .ZN(n_2115));
   NAND2_X1 i_1569 (.A1(b[29]), .A2(a[0]), .ZN(n_2117));
   OAI21_X1 i_1570 (.A(n_2114), .B1(n_2115), .B2(n_2117), .ZN(n_2557));
   INV_X1 i_1571 (.A(n_2017), .ZN(n_2118));
   NAND3_X1 i_1572 (.A1(n_2118), .A2(b[24]), .A3(a[5]), .ZN(n_2119));
   AOI21_X1 i_1573 (.A(n_2118), .B1(b[24]), .B2(a[5]), .ZN(n_2120));
   NAND2_X1 i_1574 (.A1(b[26]), .A2(a[3]), .ZN(n_2121));
   OAI21_X1 i_1575 (.A(n_2119), .B1(n_2120), .B2(n_2121), .ZN(n_2564));
   INV_X1 i_1576 (.A(n_2024), .ZN(n_2122));
   NAND3_X1 i_1587 (.A1(n_2122), .A2(b[21]), .A3(a[8]), .ZN(n_2125));
   AOI21_X1 i_1588 (.A(n_2122), .B1(b[21]), .B2(a[8]), .ZN(n_2126));
   NAND2_X1 i_1589 (.A1(b[23]), .A2(a[6]), .ZN(n_2127));
   OAI21_X1 i_1590 (.A(n_2125), .B1(n_2126), .B2(n_2127), .ZN(n_2571));
   INV_X1 i_1591 (.A(n_2030), .ZN(n_2128));
   NAND3_X1 i_1592 (.A1(n_2128), .A2(b[18]), .A3(a[11]), .ZN(n_2157));
   AOI21_X1 i_1593 (.A(n_2128), .B1(b[18]), .B2(a[11]), .ZN(n_2158));
   NAND2_X1 i_1594 (.A1(b[20]), .A2(a[9]), .ZN(n_2161));
   OAI21_X1 i_1595 (.A(n_2157), .B1(n_2158), .B2(n_2161), .ZN(n_2578));
   INV_X1 i_1596 (.A(n_2036), .ZN(n_2162));
   NAND3_X1 i_1597 (.A1(n_2162), .A2(a[14]), .A3(b[15]), .ZN(n_2163));
   AOI21_X1 i_1598 (.A(n_2162), .B1(a[14]), .B2(b[15]), .ZN(n_2164));
   NAND2_X1 i_1599 (.A1(b[17]), .A2(a[12]), .ZN(n_2165));
   OAI21_X1 i_1600 (.A(n_2163), .B1(n_2164), .B2(n_2165), .ZN(n_2585));
   INV_X1 i_1601 (.A(n_2071), .ZN(n_2168));
   NAND3_X1 i_1602 (.A1(n_2168), .A2(a[17]), .A3(b[12]), .ZN(n_2169));
   AOI21_X1 i_1603 (.A(n_2168), .B1(a[17]), .B2(b[12]), .ZN(n_2170));
   NAND2_X1 i_1604 (.A1(a[15]), .A2(b[14]), .ZN(n_2171));
   OAI21_X1 i_1605 (.A(n_2169), .B1(n_2170), .B2(n_2171), .ZN(n_2592));
   INV_X1 i_1606 (.A(n_2078), .ZN(n_2172));
   NAND3_X1 i_1607 (.A1(n_2172), .A2(a[20]), .A3(b[9]), .ZN(n_2175));
   AOI21_X1 i_1608 (.A(n_2172), .B1(a[20]), .B2(b[9]), .ZN(n_2176));
   NAND2_X1 i_1609 (.A1(a[18]), .A2(b[11]), .ZN(n_2177));
   OAI21_X1 i_1610 (.A(n_2175), .B1(n_2176), .B2(n_2177), .ZN(n_2599));
   INV_X1 i_1611 (.A(n_2085), .ZN(n_2178));
   NAND3_X1 i_1612 (.A1(n_2178), .A2(a[23]), .A3(b[6]), .ZN(n_2179));
   AOI21_X1 i_1613 (.A(n_2178), .B1(a[23]), .B2(b[6]), .ZN(n_2182));
   NAND2_X1 i_1614 (.A1(a[21]), .A2(b[8]), .ZN(n_2183));
   OAI21_X1 i_1615 (.A(n_2179), .B1(n_2182), .B2(n_2183), .ZN(n_2606));
   INV_X1 i_1616 (.A(n_2115), .ZN(n_2184));
   NAND2_X1 i_1617 (.A1(n_2114), .A2(n_2184), .ZN(n_2185));
   XOR2_X1 i_1618 (.A(n_2185), .B(n_2117), .Z(n_2556));
   INV_X1 i_1619 (.A(n_2120), .ZN(n_2186));
   NAND2_X1 i_1620 (.A1(n_2119), .A2(n_2186), .ZN(n_2189));
   XOR2_X1 i_1621 (.A(n_2189), .B(n_2121), .Z(n_2563));
   INV_X1 i_1622 (.A(n_2126), .ZN(n_2190));
   NAND2_X1 i_1623 (.A1(n_2125), .A2(n_2190), .ZN(n_2191));
   XOR2_X1 i_1624 (.A(n_2191), .B(n_2127), .Z(n_2570));
   INV_X1 i_1625 (.A(n_2158), .ZN(n_2192));
   NAND2_X1 i_1626 (.A1(n_2157), .A2(n_2192), .ZN(n_2193));
   XOR2_X1 i_1627 (.A(n_2193), .B(n_2161), .Z(n_2577));
   INV_X1 i_1628 (.A(n_2164), .ZN(n_2196));
   NAND2_X1 i_1629 (.A1(n_2163), .A2(n_2196), .ZN(n_2197));
   XOR2_X1 i_1630 (.A(n_2197), .B(n_2165), .Z(n_2584));
   INV_X1 i_1631 (.A(n_2170), .ZN(n_2198));
   NAND2_X1 i_1632 (.A1(n_2169), .A2(n_2198), .ZN(n_2199));
   XOR2_X1 i_1633 (.A(n_2199), .B(n_2171), .Z(n_2591));
   INV_X1 i_1634 (.A(n_2176), .ZN(n_2200));
   NAND2_X1 i_1635 (.A1(n_2175), .A2(n_2200), .ZN(n_2203));
   XOR2_X1 i_1636 (.A(n_2203), .B(n_2177), .Z(n_2598));
   INV_X1 i_1648 (.A(n_2182), .ZN(n_2204));
   NAND2_X1 i_1649 (.A1(n_2179), .A2(n_2204), .ZN(n_2205));
   XOR2_X1 i_1650 (.A(n_2205), .B(n_2183), .Z(n_2605));
   NAND2_X1 i_1651 (.A1(n_1992), .A2(n_1995), .ZN(n_2206));
   XNOR2_X1 i_1652 (.A(n_2206), .B(n_1994), .ZN(n_2612));
   NAND2_X1 i_1653 (.A1(n_1999), .A2(n_2002), .ZN(n_2207));
   XNOR2_X1 i_1654 (.A(n_2207), .B(n_2001), .ZN(n_2619));
   NAND4_X1 i_1655 (.A1(a[26]), .A2(a[25]), .A3(b[2]), .A4(b[1]), .ZN(n_2210));
   AOI22_X1 i_1656 (.A1(a[26]), .A2(b[1]), .B1(a[25]), .B2(b[2]), .ZN(n_2211));
   NAND2_X1 i_1657 (.A1(a[24]), .A2(b[3]), .ZN(n_2212));
   OAI21_X1 i_1658 (.A(n_2210), .B1(n_2211), .B2(n_2212), .ZN(n_2213));
   AOI21_X1 i_1659 (.A(n_2213), .B1(a[28]), .B2(b[0]), .ZN(n_2216));
   NAND2_X1 i_1660 (.A1(a[27]), .A2(b[1]), .ZN(n_2217));
   NAND3_X1 i_1661 (.A1(n_2213), .A2(a[28]), .A3(b[0]), .ZN(n_2218));
   AOI21_X1 i_1662 (.A(n_2216), .B1(n_2217), .B2(n_2218), .ZN(n_2514));
   NAND4_X1 i_1663 (.A1(b[27]), .A2(b[26]), .A3(a[2]), .A4(a[1]), .ZN(n_2219));
   AOI22_X1 i_1664 (.A1(b[26]), .A2(a[2]), .B1(b[27]), .B2(a[1]), .ZN(n_2220));
   NAND2_X1 i_1665 (.A1(b[28]), .A2(a[0]), .ZN(n_2251));
   OAI21_X1 i_1666 (.A(n_2219), .B1(n_2220), .B2(n_2251), .ZN(n_2452));
   NAND4_X1 i_1667 (.A1(b[24]), .A2(b[23]), .A3(a[5]), .A4(a[4]), .ZN(n_2252));
   AOI22_X1 i_1668 (.A1(b[23]), .A2(a[5]), .B1(b[24]), .B2(a[4]), .ZN(n_2255));
   NAND2_X1 i_1669 (.A1(b[25]), .A2(a[3]), .ZN(n_2256));
   OAI21_X1 i_1670 (.A(n_2252), .B1(n_2255), .B2(n_2256), .ZN(n_2459));
   NAND4_X1 i_1671 (.A1(b[21]), .A2(b[20]), .A3(a[8]), .A4(a[7]), .ZN(n_2257));
   AOI22_X1 i_1672 (.A1(b[20]), .A2(a[8]), .B1(b[21]), .B2(a[7]), .ZN(n_2258));
   NAND2_X1 i_1673 (.A1(b[22]), .A2(a[6]), .ZN(n_2259));
   OAI21_X1 i_1674 (.A(n_2257), .B1(n_2258), .B2(n_2259), .ZN(n_2466));
   NAND4_X1 i_1675 (.A1(b[18]), .A2(b[17]), .A3(a[11]), .A4(a[10]), .ZN(n_2262));
   AOI22_X1 i_1676 (.A1(b[17]), .A2(a[11]), .B1(b[18]), .B2(a[10]), .ZN(n_2263));
   NAND2_X1 i_1677 (.A1(b[19]), .A2(a[9]), .ZN(n_2264));
   OAI21_X1 i_1678 (.A(n_2262), .B1(n_2263), .B2(n_2264), .ZN(n_2473));
   NAND4_X1 i_1679 (.A1(a[14]), .A2(b[15]), .A3(b[14]), .A4(a[13]), .ZN(n_2265));
   AOI22_X1 i_1680 (.A1(a[14]), .A2(b[14]), .B1(b[15]), .B2(a[13]), .ZN(n_2266));
   NAND2_X1 i_1681 (.A1(b[16]), .A2(a[12]), .ZN(n_2269));
   OAI21_X1 i_1682 (.A(n_2265), .B1(n_2266), .B2(n_2269), .ZN(n_2480));
   NAND4_X1 i_1683 (.A1(a[17]), .A2(a[16]), .A3(b[12]), .A4(b[11]), .ZN(n_2270));
   AOI22_X1 i_1684 (.A1(a[17]), .A2(b[11]), .B1(a[16]), .B2(b[12]), .ZN(n_2271));
   NAND2_X1 i_1685 (.A1(a[15]), .A2(b[13]), .ZN(n_2272));
   OAI21_X1 i_1686 (.A(n_2270), .B1(n_2271), .B2(n_2272), .ZN(n_2487));
   NAND4_X1 i_1687 (.A1(a[20]), .A2(a[19]), .A3(b[9]), .A4(b[8]), .ZN(n_2273));
   AOI22_X1 i_1688 (.A1(a[20]), .A2(b[8]), .B1(a[19]), .B2(b[9]), .ZN(n_2276));
   NAND2_X1 i_1689 (.A1(a[18]), .A2(b[10]), .ZN(n_2277));
   OAI21_X1 i_1690 (.A(n_2273), .B1(n_2276), .B2(n_2277), .ZN(n_2494));
   NAND4_X1 i_1691 (.A1(a[23]), .A2(a[22]), .A3(b[6]), .A4(b[5]), .ZN(n_2278));
   AOI22_X1 i_1692 (.A1(a[23]), .A2(b[5]), .B1(a[22]), .B2(b[6]), .ZN(n_2279));
   NAND2_X1 i_1693 (.A1(a[21]), .A2(b[7]), .ZN(n_2280));
   OAI21_X1 i_1694 (.A(n_2278), .B1(n_2279), .B2(n_2280), .ZN(n_2501));
   NAND4_X1 i_1695 (.A1(a[26]), .A2(a[25]), .A3(b[3]), .A4(b[2]), .ZN(n_2283));
   AOI22_X1 i_1696 (.A1(a[26]), .A2(b[2]), .B1(a[25]), .B2(b[3]), .ZN(n_2284));
   NAND2_X1 i_1709 (.A1(a[24]), .A2(b[4]), .ZN(n_2285));
   OAI21_X1 i_1710 (.A(n_2283), .B1(n_2284), .B2(n_2285), .ZN(n_2508));
   INV_X1 i_1711 (.A(n_2220), .ZN(n_2286));
   NAND2_X1 i_1712 (.A1(n_2286), .A2(n_2219), .ZN(n_2287));
   XOR2_X1 i_1713 (.A(n_2287), .B(n_2251), .Z(n_2451));
   INV_X1 i_1714 (.A(n_2255), .ZN(n_2290));
   NAND2_X1 i_1715 (.A1(n_2290), .A2(n_2252), .ZN(n_2291));
   XOR2_X1 i_1716 (.A(n_2291), .B(n_2256), .Z(n_2458));
   INV_X1 i_1717 (.A(n_2258), .ZN(n_2292));
   NAND2_X1 i_1718 (.A1(n_2292), .A2(n_2257), .ZN(n_2293));
   XOR2_X1 i_1719 (.A(n_2293), .B(n_2259), .Z(n_2465));
   INV_X1 i_1720 (.A(n_2263), .ZN(n_2294));
   NAND2_X1 i_1721 (.A1(n_2294), .A2(n_2262), .ZN(n_2297));
   XOR2_X1 i_1722 (.A(n_2297), .B(n_2264), .Z(n_2472));
   INV_X1 i_1723 (.A(n_2266), .ZN(n_2298));
   NAND2_X1 i_1724 (.A1(n_2298), .A2(n_2265), .ZN(n_2299));
   XOR2_X1 i_1725 (.A(n_2299), .B(n_2269), .Z(n_2479));
   INV_X1 i_1726 (.A(n_2271), .ZN(n_2300));
   NAND2_X1 i_1727 (.A1(n_2300), .A2(n_2270), .ZN(n_2301));
   XOR2_X1 i_1728 (.A(n_2301), .B(n_2272), .Z(n_2486));
   INV_X1 i_1729 (.A(n_2276), .ZN(n_2303));
   NAND2_X1 i_1730 (.A1(n_2303), .A2(n_2273), .ZN(n_2304));
   XOR2_X1 i_1731 (.A(n_2304), .B(n_2277), .Z(n_2493));
   INV_X1 i_1732 (.A(n_2279), .ZN(n_2305));
   NAND2_X1 i_1733 (.A1(n_2305), .A2(n_2278), .ZN(n_2306));
   XOR2_X1 i_1734 (.A(n_2306), .B(n_2280), .Z(n_2500));
   INV_X1 i_1735 (.A(n_2284), .ZN(n_2307));
   NAND2_X1 i_1736 (.A1(n_2307), .A2(n_2283), .ZN(n_2308));
   XOR2_X1 i_1737 (.A(n_2308), .B(n_2285), .Z(n_2507));
   INV_X1 i_1738 (.A(n_2216), .ZN(n_2310));
   NAND2_X1 i_1739 (.A1(n_2310), .A2(n_2218), .ZN(n_2311));
   XOR2_X1 i_1740 (.A(n_2311), .B(n_2217), .Z(n_2513));
   NAND4_X1 i_1741 (.A1(a[23]), .A2(a[22]), .A3(b[3]), .A4(b[4]), .ZN(n_2312));
   AOI22_X1 i_1742 (.A1(a[23]), .A2(b[3]), .B1(a[22]), .B2(b[4]), .ZN(n_2313));
   NAND2_X1 i_1743 (.A1(a[21]), .A2(b[5]), .ZN(n_2346));
   OAI21_X1 i_1744 (.A(n_2312), .B1(n_2313), .B2(n_2346), .ZN(n_2347));
   NAND4_X1 i_1745 (.A1(a[26]), .A2(a[25]), .A3(b[1]), .A4(b[0]), .ZN(n_2350));
   AOI22_X1 i_1746 (.A1(a[26]), .A2(b[0]), .B1(a[25]), .B2(b[1]), .ZN(n_2351));
   NAND2_X1 i_1747 (.A1(a[24]), .A2(b[2]), .ZN(n_2352));
   OAI21_X1 i_1748 (.A(n_2350), .B1(n_2351), .B2(n_2352), .ZN(n_2353));
   NOR2_X1 i_1749 (.A1(n_2347), .A2(n_2353), .ZN(n_2354));
   NAND2_X1 i_1750 (.A1(a[27]), .A2(b[0]), .ZN(n_2357));
   NAND2_X1 i_1751 (.A1(n_2347), .A2(n_2353), .ZN(n_2358));
   AOI21_X1 i_1752 (.A(n_2354), .B1(n_2357), .B2(n_2358), .ZN(n_2412));
   NAND4_X1 i_1753 (.A1(b[26]), .A2(b[25]), .A3(a[2]), .A4(a[1]), .ZN(n_2359));
   AOI22_X1 i_1754 (.A1(b[25]), .A2(a[2]), .B1(b[26]), .B2(a[1]), .ZN(n_2360));
   NAND2_X1 i_1755 (.A1(b[27]), .A2(a[0]), .ZN(n_2361));
   OAI21_X1 i_1756 (.A(n_2359), .B1(n_2360), .B2(n_2361), .ZN(n_2349));
   NAND4_X1 i_1757 (.A1(b[23]), .A2(b[22]), .A3(a[5]), .A4(a[4]), .ZN(n_2364));
   AOI22_X1 i_1758 (.A1(b[22]), .A2(a[5]), .B1(b[23]), .B2(a[4]), .ZN(n_2365));
   NAND2_X1 i_1759 (.A1(b[24]), .A2(a[3]), .ZN(n_2366));
   OAI21_X1 i_1760 (.A(n_2364), .B1(n_2365), .B2(n_2366), .ZN(n_2356));
   NAND4_X1 i_1761 (.A1(b[20]), .A2(b[19]), .A3(a[8]), .A4(a[7]), .ZN(n_2367));
   AOI22_X1 i_1762 (.A1(b[19]), .A2(a[8]), .B1(b[20]), .B2(a[7]), .ZN(n_2368));
   NAND2_X1 i_1763 (.A1(b[21]), .A2(a[6]), .ZN(n_2371));
   OAI21_X1 i_1764 (.A(n_2367), .B1(n_2368), .B2(n_2371), .ZN(n_2363));
   NAND4_X1 i_1765 (.A1(b[17]), .A2(b[16]), .A3(a[11]), .A4(a[10]), .ZN(n_2372));
   AOI22_X1 i_1778 (.A1(b[16]), .A2(a[11]), .B1(b[17]), .B2(a[10]), .ZN(n_2373));
   NAND2_X1 i_1779 (.A1(b[18]), .A2(a[9]), .ZN(n_2374));
   OAI21_X1 i_1780 (.A(n_2372), .B1(n_2373), .B2(n_2374), .ZN(n_2370));
   NAND4_X1 i_1781 (.A1(a[14]), .A2(b[14]), .A3(a[13]), .A4(b[13]), .ZN(n_2375));
   AOI22_X1 i_1782 (.A1(a[14]), .A2(b[13]), .B1(b[14]), .B2(a[13]), .ZN(n_2378));
   NAND2_X1 i_1783 (.A1(b[15]), .A2(a[12]), .ZN(n_2379));
   OAI21_X1 i_1784 (.A(n_2375), .B1(n_2378), .B2(n_2379), .ZN(n_2377));
   NAND4_X1 i_1785 (.A1(a[17]), .A2(a[16]), .A3(b[11]), .A4(b[10]), .ZN(n_2380));
   AOI22_X1 i_1786 (.A1(a[17]), .A2(b[10]), .B1(a[16]), .B2(b[11]), .ZN(n_2381));
   NAND2_X1 i_1787 (.A1(a[15]), .A2(b[12]), .ZN(n_2382));
   OAI21_X1 i_1788 (.A(n_2380), .B1(n_2381), .B2(n_2382), .ZN(n_2384));
   NAND4_X1 i_1789 (.A1(a[20]), .A2(a[19]), .A3(b[8]), .A4(b[7]), .ZN(n_2385));
   AOI22_X1 i_1790 (.A1(a[20]), .A2(b[7]), .B1(a[19]), .B2(b[8]), .ZN(n_2386));
   NAND2_X1 i_1791 (.A1(a[18]), .A2(b[9]), .ZN(n_2387));
   OAI21_X1 i_1792 (.A(n_2385), .B1(n_2386), .B2(n_2387), .ZN(n_2391));
   NAND4_X1 i_1793 (.A1(a[23]), .A2(a[22]), .A3(b[4]), .A4(b[5]), .ZN(n_2388));
   AOI22_X1 i_1794 (.A1(a[23]), .A2(b[4]), .B1(a[22]), .B2(b[5]), .ZN(n_2389));
   NAND2_X1 i_1795 (.A1(a[21]), .A2(b[6]), .ZN(n_2392));
   OAI21_X1 i_1796 (.A(n_2388), .B1(n_2389), .B2(n_2392), .ZN(n_2398));
   INV_X1 i_1797 (.A(n_2354), .ZN(n_2393));
   NAND2_X1 i_1798 (.A1(n_2393), .A2(n_2358), .ZN(n_2394));
   XOR2_X1 i_1799 (.A(n_2394), .B(n_2357), .Z(n_2411));
   INV_X1 i_1800 (.A(n_2360), .ZN(n_2395));
   NAND2_X1 i_1801 (.A1(n_2395), .A2(n_2359), .ZN(n_2396));
   XOR2_X1 i_1802 (.A(n_2396), .B(n_2361), .Z(n_2348));
   INV_X1 i_1803 (.A(n_2365), .ZN(n_2399));
   NAND2_X1 i_1804 (.A1(n_2399), .A2(n_2364), .ZN(n_2400));
   XOR2_X1 i_1805 (.A(n_2400), .B(n_2366), .Z(n_2355));
   INV_X1 i_1806 (.A(n_2368), .ZN(n_2401));
   NAND2_X1 i_1807 (.A1(n_2401), .A2(n_2367), .ZN(n_2402));
   XOR2_X1 i_1808 (.A(n_2402), .B(n_2371), .Z(n_2362));
   INV_X1 i_1809 (.A(n_2373), .ZN(n_2403));
   NAND2_X1 i_1810 (.A1(n_2403), .A2(n_2372), .ZN(n_2405));
   XOR2_X1 i_1811 (.A(n_2405), .B(n_2374), .Z(n_2369));
   INV_X1 i_1812 (.A(n_2378), .ZN(n_2406));
   NAND2_X1 i_1813 (.A1(n_2406), .A2(n_2375), .ZN(n_2407));
   XOR2_X1 i_1814 (.A(n_2407), .B(n_2379), .Z(n_2376));
   INV_X1 i_1815 (.A(n_2381), .ZN(n_2408));
   NAND2_X1 i_1816 (.A1(n_2408), .A2(n_2380), .ZN(n_2409));
   XOR2_X1 i_1817 (.A(n_2409), .B(n_2382), .Z(n_2383));
   INV_X1 i_1818 (.A(n_2386), .ZN(n_2410));
   NAND2_X1 i_1819 (.A1(n_2410), .A2(n_2385), .ZN(n_2413));
   XOR2_X1 i_1820 (.A(n_2413), .B(n_2387), .Z(n_2390));
   INV_X1 i_1821 (.A(n_2389), .ZN(n_2414));
   NAND2_X1 i_1822 (.A1(n_2414), .A2(n_2388), .ZN(n_2415));
   XOR2_X1 i_1823 (.A(n_2415), .B(n_2392), .Z(n_2397));
   INV_X1 i_1824 (.A(n_2211), .ZN(n_2416));
   NAND2_X1 i_1825 (.A1(n_2416), .A2(n_2210), .ZN(n_2449));
   XOR2_X1 i_1826 (.A(n_2449), .B(n_2212), .Z(n_2404));
   NAND4_X1 i_1827 (.A1(b[25]), .A2(b[24]), .A3(a[2]), .A4(a[1]), .ZN(n_2450));
   AOI22_X1 i_1828 (.A1(b[24]), .A2(a[2]), .B1(b[25]), .B2(a[1]), .ZN(n_2453));
   NAND2_X1 i_1829 (.A1(b[26]), .A2(a[0]), .ZN(n_2454));
   OAI21_X1 i_1830 (.A(n_2450), .B1(n_2453), .B2(n_2454), .ZN(n_2254));
   NAND4_X1 i_1831 (.A1(b[22]), .A2(b[21]), .A3(a[5]), .A4(a[4]), .ZN(n_2455));
   AOI22_X1 i_1832 (.A1(b[21]), .A2(a[5]), .B1(b[22]), .B2(a[4]), .ZN(n_2456));
   NAND2_X1 i_1833 (.A1(b[23]), .A2(a[3]), .ZN(n_2457));
   OAI21_X1 i_1834 (.A(n_2455), .B1(n_2456), .B2(n_2457), .ZN(n_2261));
   NAND4_X1 i_1848 (.A1(b[19]), .A2(b[18]), .A3(a[8]), .A4(a[7]), .ZN(n_2460));
   AOI22_X1 i_1849 (.A1(b[18]), .A2(a[8]), .B1(b[19]), .B2(a[7]), .ZN(n_2461));
   NAND2_X1 i_1850 (.A1(b[20]), .A2(a[6]), .ZN(n_2462));
   OAI21_X1 i_1851 (.A(n_2460), .B1(n_2461), .B2(n_2462), .ZN(n_2268));
   NAND4_X1 i_1852 (.A1(b[16]), .A2(b[15]), .A3(a[11]), .A4(a[10]), .ZN(n_2463));
   AOI22_X1 i_1853 (.A1(b[15]), .A2(a[11]), .B1(b[16]), .B2(a[10]), .ZN(n_2464));
   NAND2_X1 i_1854 (.A1(b[17]), .A2(a[9]), .ZN(n_2467));
   OAI21_X1 i_1855 (.A(n_2463), .B1(n_2464), .B2(n_2467), .ZN(n_2275));
   NAND4_X1 i_1856 (.A1(a[14]), .A2(a[13]), .A3(b[13]), .A4(b[12]), .ZN(n_2468));
   AOI22_X1 i_1857 (.A1(a[14]), .A2(b[12]), .B1(a[13]), .B2(b[13]), .ZN(n_2469));
   NAND2_X1 i_1858 (.A1(b[14]), .A2(a[12]), .ZN(n_2470));
   OAI21_X1 i_1859 (.A(n_2468), .B1(n_2469), .B2(n_2470), .ZN(n_2282));
   NAND4_X1 i_1860 (.A1(a[17]), .A2(a[16]), .A3(b[10]), .A4(b[9]), .ZN(n_2471));
   AOI22_X1 i_1861 (.A1(a[17]), .A2(b[9]), .B1(a[16]), .B2(b[10]), .ZN(n_2474));
   NAND2_X1 i_1862 (.A1(a[15]), .A2(b[11]), .ZN(n_2475));
   OAI21_X1 i_1863 (.A(n_2471), .B1(n_2474), .B2(n_2475), .ZN(n_2289));
   NAND4_X1 i_1864 (.A1(a[20]), .A2(a[19]), .A3(b[7]), .A4(b[6]), .ZN(n_2476));
   AOI22_X1 i_1865 (.A1(a[20]), .A2(b[6]), .B1(a[19]), .B2(b[7]), .ZN(n_2477));
   NAND2_X1 i_1866 (.A1(a[18]), .A2(b[8]), .ZN(n_2478));
   OAI21_X1 i_1867 (.A(n_2476), .B1(n_2477), .B2(n_2478), .ZN(n_2296));
   INV_X1 i_1868 (.A(n_2453), .ZN(n_2481));
   NAND2_X1 i_1869 (.A1(n_2481), .A2(n_2450), .ZN(n_2482));
   XOR2_X1 i_1870 (.A(n_2482), .B(n_2454), .Z(n_2253));
   INV_X1 i_1871 (.A(n_2456), .ZN(n_2483));
   NAND2_X1 i_1872 (.A1(n_2483), .A2(n_2455), .ZN(n_2484));
   XOR2_X1 i_1873 (.A(n_2484), .B(n_2457), .Z(n_2260));
   INV_X1 i_1874 (.A(n_2461), .ZN(n_2485));
   NAND2_X1 i_1875 (.A1(n_2485), .A2(n_2460), .ZN(n_2488));
   XOR2_X1 i_1876 (.A(n_2488), .B(n_2462), .Z(n_2267));
   INV_X1 i_1877 (.A(n_2464), .ZN(n_2489));
   NAND2_X1 i_1878 (.A1(n_2489), .A2(n_2463), .ZN(n_2490));
   XOR2_X1 i_1879 (.A(n_2490), .B(n_2467), .Z(n_2274));
   INV_X1 i_1880 (.A(n_2469), .ZN(n_2491));
   NAND2_X1 i_1881 (.A1(n_2491), .A2(n_2468), .ZN(n_2492));
   XOR2_X1 i_1882 (.A(n_2492), .B(n_2470), .Z(n_2281));
   INV_X1 i_1883 (.A(n_2474), .ZN(n_2495));
   NAND2_X1 i_1884 (.A1(n_2495), .A2(n_2471), .ZN(n_2496));
   XOR2_X1 i_1885 (.A(n_2496), .B(n_2475), .Z(n_2288));
   INV_X1 i_1886 (.A(n_2477), .ZN(n_2497));
   NAND2_X1 i_1887 (.A1(n_2497), .A2(n_2476), .ZN(n_2498));
   XOR2_X1 i_1888 (.A(n_2498), .B(n_2478), .Z(n_2295));
   INV_X1 i_1889 (.A(n_2313), .ZN(n_2499));
   NAND2_X1 i_1890 (.A1(n_2499), .A2(n_2312), .ZN(n_2502));
   XOR2_X1 i_1891 (.A(n_2502), .B(n_2346), .Z(n_2302));
   INV_X1 i_1892 (.A(n_2351), .ZN(n_2503));
   NAND2_X1 i_1893 (.A1(n_2503), .A2(n_2350), .ZN(n_2504));
   XOR2_X1 i_1894 (.A(n_2504), .B(n_2352), .Z(n_2309));
   NAND4_X1 i_1895 (.A1(a[23]), .A2(a[22]), .A3(b[2]), .A4(b[1]), .ZN(n_2505));
   AOI22_X1 i_1896 (.A1(a[23]), .A2(b[1]), .B1(a[22]), .B2(b[2]), .ZN(n_2506));
   NAND2_X1 i_1897 (.A1(a[21]), .A2(b[3]), .ZN(n_2509));
   OAI21_X1 i_1898 (.A(n_2505), .B1(n_2506), .B2(n_2509), .ZN(n_2510));
   AOI21_X1 i_1899 (.A(n_2510), .B1(a[25]), .B2(b[0]), .ZN(n_2511));
   NAND2_X1 i_1900 (.A1(a[24]), .A2(b[1]), .ZN(n_2512));
   NAND3_X1 i_1901 (.A1(n_2510), .A2(a[25]), .A3(b[0]), .ZN(n_2515));
   AOI21_X1 i_1902 (.A(n_2511), .B1(n_2512), .B2(n_2515), .ZN(n_2215));
   NAND4_X1 i_1903 (.A1(b[24]), .A2(b[23]), .A3(a[2]), .A4(a[1]), .ZN(n_2516));
   AOI22_X1 i_1918 (.A1(b[23]), .A2(a[2]), .B1(b[24]), .B2(a[1]), .ZN(n_2517));
   NAND2_X1 i_1919 (.A1(b[25]), .A2(a[0]), .ZN(n_2518));
   OAI21_X1 i_1920 (.A(n_2516), .B1(n_2517), .B2(n_2518), .ZN(n_2160));
   NAND4_X1 i_1921 (.A1(b[21]), .A2(b[20]), .A3(a[5]), .A4(a[4]), .ZN(n_2519));
   AOI22_X1 i_1922 (.A1(b[20]), .A2(a[5]), .B1(b[21]), .B2(a[4]), .ZN(n_2554));
   NAND2_X1 i_1923 (.A1(b[22]), .A2(a[3]), .ZN(n_2555));
   OAI21_X1 i_1924 (.A(n_2519), .B1(n_2554), .B2(n_2555), .ZN(n_2167));
   NAND4_X1 i_1925 (.A1(b[18]), .A2(b[17]), .A3(a[8]), .A4(a[7]), .ZN(n_2558));
   AOI22_X1 i_1926 (.A1(b[17]), .A2(a[8]), .B1(b[18]), .B2(a[7]), .ZN(n_2559));
   NAND2_X1 i_1927 (.A1(b[19]), .A2(a[6]), .ZN(n_2560));
   OAI21_X1 i_1928 (.A(n_2558), .B1(n_2559), .B2(n_2560), .ZN(n_2174));
   NAND4_X1 i_1929 (.A1(b[15]), .A2(b[14]), .A3(a[11]), .A4(a[10]), .ZN(n_2561));
   AOI22_X1 i_1930 (.A1(b[14]), .A2(a[11]), .B1(b[15]), .B2(a[10]), .ZN(n_2562));
   NAND2_X1 i_1931 (.A1(b[16]), .A2(a[9]), .ZN(n_2565));
   OAI21_X1 i_1932 (.A(n_2561), .B1(n_2562), .B2(n_2565), .ZN(n_2181));
   NAND4_X1 i_1933 (.A1(a[14]), .A2(a[13]), .A3(b[12]), .A4(b[11]), .ZN(n_2566));
   AOI22_X1 i_1934 (.A1(a[14]), .A2(b[11]), .B1(a[13]), .B2(b[12]), .ZN(n_2567));
   NAND2_X1 i_1935 (.A1(b[13]), .A2(a[12]), .ZN(n_2568));
   OAI21_X1 i_1936 (.A(n_2566), .B1(n_2567), .B2(n_2568), .ZN(n_2188));
   NAND4_X1 i_1937 (.A1(a[17]), .A2(a[16]), .A3(b[9]), .A4(b[8]), .ZN(n_2569));
   AOI22_X1 i_1938 (.A1(a[17]), .A2(b[8]), .B1(a[16]), .B2(b[9]), .ZN(n_2572));
   NAND2_X1 i_1939 (.A1(a[15]), .A2(b[10]), .ZN(n_2573));
   OAI21_X1 i_1940 (.A(n_2569), .B1(n_2572), .B2(n_2573), .ZN(n_2195));
   NAND4_X1 i_1941 (.A1(a[20]), .A2(a[19]), .A3(b[6]), .A4(b[5]), .ZN(n_2574));
   AOI22_X1 i_1942 (.A1(a[20]), .A2(b[5]), .B1(a[19]), .B2(b[6]), .ZN(n_2575));
   NAND2_X1 i_1943 (.A1(a[18]), .A2(b[7]), .ZN(n_2576));
   OAI21_X1 i_1944 (.A(n_2574), .B1(n_2575), .B2(n_2576), .ZN(n_2202));
   NAND4_X1 i_1945 (.A1(a[23]), .A2(a[22]), .A3(b[3]), .A4(b[2]), .ZN(n_2579));
   AOI22_X1 i_1946 (.A1(a[23]), .A2(b[2]), .B1(a[22]), .B2(b[3]), .ZN(n_2580));
   NAND2_X1 i_1947 (.A1(a[21]), .A2(b[4]), .ZN(n_2581));
   OAI21_X1 i_1948 (.A(n_2579), .B1(n_2580), .B2(n_2581), .ZN(n_2209));
   INV_X1 i_1949 (.A(n_2517), .ZN(n_2582));
   NAND2_X1 i_1950 (.A1(n_2582), .A2(n_2516), .ZN(n_2583));
   XOR2_X1 i_1951 (.A(n_2583), .B(n_2518), .Z(n_2159));
   INV_X1 i_1952 (.A(n_2554), .ZN(n_2586));
   NAND2_X1 i_1953 (.A1(n_2586), .A2(n_2519), .ZN(n_2587));
   XOR2_X1 i_1954 (.A(n_2587), .B(n_2555), .Z(n_2166));
   INV_X1 i_1955 (.A(n_2559), .ZN(n_2588));
   NAND2_X1 i_1956 (.A1(n_2588), .A2(n_2558), .ZN(n_2589));
   XOR2_X1 i_1957 (.A(n_2589), .B(n_2560), .Z(n_2173));
   INV_X1 i_1958 (.A(n_2562), .ZN(n_2590));
   NAND2_X1 i_1959 (.A1(n_2590), .A2(n_2561), .ZN(n_2593));
   XOR2_X1 i_1960 (.A(n_2593), .B(n_2565), .Z(n_2180));
   INV_X1 i_1961 (.A(n_2567), .ZN(n_2594));
   NAND2_X1 i_1962 (.A1(n_2594), .A2(n_2566), .ZN(n_2595));
   XOR2_X1 i_1963 (.A(n_2595), .B(n_2568), .Z(n_2187));
   INV_X1 i_1964 (.A(n_2572), .ZN(n_2596));
   NAND2_X1 i_1965 (.A1(n_2596), .A2(n_2569), .ZN(n_2597));
   XOR2_X1 i_1966 (.A(n_2597), .B(n_2573), .Z(n_2194));
   INV_X1 i_1967 (.A(n_2575), .ZN(n_2600));
   NAND2_X1 i_1968 (.A1(n_2600), .A2(n_2574), .ZN(n_2601));
   XOR2_X1 i_1969 (.A(n_2601), .B(n_2576), .Z(n_2201));
   INV_X1 i_1970 (.A(n_2580), .ZN(n_2602));
   NAND2_X1 i_1971 (.A1(n_2602), .A2(n_2579), .ZN(n_2603));
   XOR2_X1 i_1972 (.A(n_2603), .B(n_2581), .Z(n_2208));
   INV_X1 i_1973 (.A(n_2511), .ZN(n_2604));
   NAND2_X1 i_1974 (.A1(n_2604), .A2(n_2515), .ZN(n_2607));
   XOR2_X1 i_1975 (.A(n_2607), .B(n_2512), .Z(n_2214));
   NAND4_X1 i_1976 (.A1(a[20]), .A2(a[19]), .A3(b[3]), .A4(b[4]), .ZN(n_2608));
   AOI22_X1 i_1977 (.A1(a[20]), .A2(b[3]), .B1(a[19]), .B2(b[4]), .ZN(n_2609));
   NAND2_X1 i_1978 (.A1(a[18]), .A2(b[5]), .ZN(n_2610));
   OAI21_X1 i_1979 (.A(n_2608), .B1(n_2609), .B2(n_2610), .ZN(n_2611));
   NAND4_X1 i_1980 (.A1(a[23]), .A2(a[22]), .A3(b[1]), .A4(b[0]), .ZN(n_2613));
   AOI22_X1 i_1981 (.A1(a[23]), .A2(b[0]), .B1(a[22]), .B2(b[1]), .ZN(n_2614));
   NAND2_X1 i_1996 (.A1(a[21]), .A2(b[2]), .ZN(n_2615));
   OAI21_X1 i_1997 (.A(n_2613), .B1(n_2614), .B2(n_2615), .ZN(n_2616));
   NOR2_X1 i_1998 (.A1(n_2611), .A2(n_2616), .ZN(n_2617));
   NAND2_X1 i_1999 (.A1(a[24]), .A2(b[0]), .ZN(n_2618));
   NAND2_X1 i_2000 (.A1(n_2611), .A2(n_2616), .ZN(n_2620));
   AOI21_X1 i_2001 (.A(n_2617), .B1(n_2618), .B2(n_2620), .ZN(n_2124));
   NAND4_X1 i_2002 (.A1(b[23]), .A2(b[22]), .A3(a[2]), .A4(a[1]), .ZN(n_2621));
   AOI22_X1 i_2003 (.A1(b[22]), .A2(a[2]), .B1(b[23]), .B2(a[1]), .ZN(n_2622));
   NAND2_X1 i_2004 (.A1(b[24]), .A2(a[0]), .ZN(n_2623));
   OAI21_X1 i_2005 (.A(n_2621), .B1(n_2622), .B2(n_2623), .ZN(n_2068));
   NAND4_X1 i_2006 (.A1(b[20]), .A2(b[19]), .A3(a[5]), .A4(a[4]), .ZN(n_2660));
   AOI22_X1 i_2007 (.A1(b[19]), .A2(a[5]), .B1(b[20]), .B2(a[4]), .ZN(n_2661));
   NAND2_X1 i_2008 (.A1(b[21]), .A2(a[3]), .ZN(n_2664));
   OAI21_X1 i_2009 (.A(n_2660), .B1(n_2661), .B2(n_2664), .ZN(n_2075));
   NAND4_X1 i_2010 (.A1(b[17]), .A2(b[16]), .A3(a[8]), .A4(a[7]), .ZN(n_2665));
   AOI22_X1 i_2011 (.A1(b[16]), .A2(a[8]), .B1(b[17]), .B2(a[7]), .ZN(n_2666));
   NAND2_X1 i_2012 (.A1(b[18]), .A2(a[6]), .ZN(n_2667));
   OAI21_X1 i_2013 (.A(n_2665), .B1(n_2666), .B2(n_2667), .ZN(n_2082));
   NAND4_X1 i_2014 (.A1(b[14]), .A2(b[13]), .A3(a[11]), .A4(a[10]), .ZN(n_2668));
   AOI22_X1 i_2015 (.A1(b[13]), .A2(a[11]), .B1(b[14]), .B2(a[10]), .ZN(n_2671));
   NAND2_X1 i_2016 (.A1(b[15]), .A2(a[9]), .ZN(n_2672));
   OAI21_X1 i_2017 (.A(n_2668), .B1(n_2671), .B2(n_2672), .ZN(n_2089));
   NAND4_X1 i_2018 (.A1(a[14]), .A2(a[13]), .A3(b[11]), .A4(b[10]), .ZN(n_2673));
   AOI22_X1 i_2019 (.A1(a[14]), .A2(b[10]), .B1(a[13]), .B2(b[11]), .ZN(n_2674));
   NAND2_X1 i_2020 (.A1(a[12]), .A2(b[12]), .ZN(n_2675));
   OAI21_X1 i_2021 (.A(n_2673), .B1(n_2674), .B2(n_2675), .ZN(n_2096));
   NAND4_X1 i_2022 (.A1(a[17]), .A2(a[16]), .A3(b[8]), .A4(b[7]), .ZN(n_2678));
   AOI22_X1 i_2023 (.A1(a[17]), .A2(b[7]), .B1(a[16]), .B2(b[8]), .ZN(n_2679));
   NAND2_X1 i_2024 (.A1(a[15]), .A2(b[9]), .ZN(n_2680));
   OAI21_X1 i_2025 (.A(n_2678), .B1(n_2679), .B2(n_2680), .ZN(n_2103));
   NAND4_X1 i_2026 (.A1(a[20]), .A2(a[19]), .A3(b[4]), .A4(b[5]), .ZN(n_2681));
   AOI22_X1 i_2027 (.A1(a[20]), .A2(b[4]), .B1(a[19]), .B2(b[5]), .ZN(n_2682));
   NAND2_X1 i_2028 (.A1(a[18]), .A2(b[6]), .ZN(n_2685));
   OAI21_X1 i_2029 (.A(n_2681), .B1(n_2682), .B2(n_2685), .ZN(n_2110));
   INV_X1 i_2030 (.A(n_2617), .ZN(n_2686));
   NAND2_X1 i_2031 (.A1(n_2686), .A2(n_2620), .ZN(n_2687));
   XOR2_X1 i_2032 (.A(n_2687), .B(n_2618), .Z(n_2123));
   INV_X1 i_2033 (.A(n_2622), .ZN(n_2688));
   NAND2_X1 i_2034 (.A1(n_2688), .A2(n_2621), .ZN(n_2689));
   XOR2_X1 i_2035 (.A(n_2689), .B(n_2623), .Z(n_2067));
   INV_X1 i_2036 (.A(n_2661), .ZN(n_2692));
   NAND2_X1 i_2037 (.A1(n_2692), .A2(n_2660), .ZN(n_2693));
   XOR2_X1 i_2038 (.A(n_2693), .B(n_2664), .Z(n_2074));
   INV_X1 i_2039 (.A(n_2666), .ZN(n_2694));
   NAND2_X1 i_2040 (.A1(n_2694), .A2(n_2665), .ZN(n_2695));
   XOR2_X1 i_2041 (.A(n_2695), .B(n_2667), .Z(n_2081));
   INV_X1 i_2042 (.A(n_2671), .ZN(n_2696));
   NAND2_X1 i_2043 (.A1(n_2696), .A2(n_2668), .ZN(n_2699));
   XOR2_X1 i_2044 (.A(n_2699), .B(n_2672), .Z(n_2088));
   INV_X1 i_2045 (.A(n_2674), .ZN(n_2700));
   NAND2_X1 i_2046 (.A1(n_2700), .A2(n_2673), .ZN(n_2701));
   XOR2_X1 i_2047 (.A(n_2701), .B(n_2675), .Z(n_2095));
   INV_X1 i_2048 (.A(n_2679), .ZN(n_2702));
   NAND2_X1 i_2049 (.A1(n_2702), .A2(n_2678), .ZN(n_2703));
   XOR2_X1 i_2050 (.A(n_2703), .B(n_2680), .Z(n_2102));
   INV_X1 i_2051 (.A(n_2682), .ZN(n_2706));
   NAND2_X1 i_2052 (.A1(n_2706), .A2(n_2681), .ZN(n_2707));
   XOR2_X1 i_2053 (.A(n_2707), .B(n_2685), .Z(n_2109));
   INV_X1 i_2054 (.A(n_2506), .ZN(n_2708));
   NAND2_X1 i_2055 (.A1(n_2708), .A2(n_2505), .ZN(n_2709));
   XOR2_X1 i_2056 (.A(n_2709), .B(n_2509), .Z(n_2116));
   NAND4_X1 i_2057 (.A1(b[22]), .A2(b[21]), .A3(a[2]), .A4(a[1]), .ZN(n_2710));
   AOI22_X1 i_2058 (.A1(b[21]), .A2(a[2]), .B1(b[22]), .B2(a[1]), .ZN(n_2713));
   NAND2_X1 i_2059 (.A1(b[23]), .A2(a[0]), .ZN(n_2714));
   OAI21_X1 i_2075 (.A(n_2710), .B1(n_2713), .B2(n_2714), .ZN(n_1984));
   NAND4_X1 i_2076 (.A1(b[19]), .A2(b[18]), .A3(a[5]), .A4(a[4]), .ZN(n_2715));
   AOI22_X1 i_2077 (.A1(b[18]), .A2(a[5]), .B1(b[19]), .B2(a[4]), .ZN(n_2716));
   NAND2_X1 i_2078 (.A1(b[20]), .A2(a[3]), .ZN(n_2717));
   OAI21_X1 i_2079 (.A(n_2715), .B1(n_2716), .B2(n_2717), .ZN(n_1991));
   NAND4_X1 i_2080 (.A1(b[16]), .A2(b[15]), .A3(a[8]), .A4(a[7]), .ZN(n_2720));
   AOI22_X1 i_2081 (.A1(b[15]), .A2(a[8]), .B1(b[16]), .B2(a[7]), .ZN(n_2721));
   NAND2_X1 i_2082 (.A1(b[17]), .A2(a[6]), .ZN(n_2722));
   OAI21_X1 i_2083 (.A(n_2720), .B1(n_2721), .B2(n_2722), .ZN(n_1998));
   NAND4_X1 i_2084 (.A1(b[13]), .A2(a[11]), .A3(b[12]), .A4(a[10]), .ZN(n_2723));
   AOI22_X1 i_2085 (.A1(a[11]), .A2(b[12]), .B1(b[13]), .B2(a[10]), .ZN(n_2724));
   NAND2_X1 i_2086 (.A1(b[14]), .A2(a[9]), .ZN(n_2726));
   OAI21_X1 i_2087 (.A(n_2723), .B1(n_2724), .B2(n_2726), .ZN(n_2005));
   NAND4_X1 i_2088 (.A1(a[14]), .A2(a[13]), .A3(b[10]), .A4(b[9]), .ZN(n_2727));
   AOI22_X1 i_2089 (.A1(a[14]), .A2(b[9]), .B1(a[13]), .B2(b[10]), .ZN(n_2728));
   NAND2_X1 i_2090 (.A1(a[12]), .A2(b[11]), .ZN(n_2729));
   OAI21_X1 i_2091 (.A(n_2727), .B1(n_2728), .B2(n_2729), .ZN(n_2012));
   NAND4_X1 i_2092 (.A1(a[17]), .A2(a[16]), .A3(b[7]), .A4(b[6]), .ZN(n_2730));
   AOI22_X1 i_2093 (.A1(a[17]), .A2(b[6]), .B1(a[16]), .B2(b[7]), .ZN(n_2731));
   NAND2_X1 i_2094 (.A1(a[15]), .A2(b[8]), .ZN(n_2734));
   OAI21_X1 i_2095 (.A(n_2730), .B1(n_2731), .B2(n_2734), .ZN(n_2019));
   INV_X1 i_2096 (.A(n_2713), .ZN(n_2735));
   NAND2_X1 i_2097 (.A1(n_2735), .A2(n_2710), .ZN(n_2736));
   XOR2_X1 i_2098 (.A(n_2736), .B(n_2714), .Z(n_1983));
   INV_X1 i_2099 (.A(n_2716), .ZN(n_2737));
   NAND2_X1 i_2100 (.A1(n_2737), .A2(n_2715), .ZN(n_2774));
   XOR2_X1 i_2101 (.A(n_2774), .B(n_2717), .Z(n_1990));
   INV_X1 i_2102 (.A(n_2721), .ZN(n_2775));
   NAND2_X1 i_2103 (.A1(n_2775), .A2(n_2720), .ZN(n_2778));
   XOR2_X1 i_2104 (.A(n_2778), .B(n_2722), .Z(n_1997));
   INV_X1 i_2105 (.A(n_2724), .ZN(n_2779));
   NAND2_X1 i_2106 (.A1(n_2779), .A2(n_2723), .ZN(n_2780));
   XOR2_X1 i_2107 (.A(n_2780), .B(n_2726), .Z(n_2004));
   INV_X1 i_2108 (.A(n_2728), .ZN(n_2781));
   NAND2_X1 i_2109 (.A1(n_2781), .A2(n_2727), .ZN(n_2782));
   XOR2_X1 i_2110 (.A(n_2782), .B(n_2729), .Z(n_2011));
   INV_X1 i_2111 (.A(n_2731), .ZN(n_2785));
   NAND2_X1 i_2112 (.A1(n_2785), .A2(n_2730), .ZN(n_2786));
   XOR2_X1 i_2113 (.A(n_2786), .B(n_2734), .Z(n_2018));
   INV_X1 i_2114 (.A(n_2609), .ZN(n_2787));
   NAND2_X1 i_2115 (.A1(n_2787), .A2(n_2608), .ZN(n_2788));
   XOR2_X1 i_2116 (.A(n_2788), .B(n_2610), .Z(n_2025));
   INV_X1 i_2117 (.A(n_2614), .ZN(n_2789));
   NAND2_X1 i_2118 (.A1(n_2789), .A2(n_2613), .ZN(n_2792));
   XOR2_X1 i_2119 (.A(n_2792), .B(n_2615), .Z(n_2032));
   NAND4_X1 i_2120 (.A1(a[20]), .A2(a[19]), .A3(b[2]), .A4(b[1]), .ZN(n_2793));
   AOI22_X1 i_2121 (.A1(a[20]), .A2(b[1]), .B1(a[19]), .B2(b[2]), .ZN(n_2794));
   NAND2_X1 i_2122 (.A1(a[18]), .A2(b[3]), .ZN(n_2795));
   OAI21_X1 i_2123 (.A(n_2793), .B1(n_2794), .B2(n_2795), .ZN(n_2796));
   AOI21_X1 i_2124 (.A(n_2796), .B1(a[22]), .B2(b[0]), .ZN(n_2799));
   NAND2_X1 i_2125 (.A1(a[21]), .A2(b[1]), .ZN(n_2800));
   NAND3_X1 i_2126 (.A1(n_2796), .A2(a[22]), .A3(b[0]), .ZN(n_2801));
   AOI21_X1 i_2127 (.A(n_2799), .B1(n_2800), .B2(n_2801), .ZN(n_1949));
   NAND4_X1 i_2128 (.A1(b[21]), .A2(b[20]), .A3(a[2]), .A4(a[1]), .ZN(n_2802));
   AOI22_X1 i_2129 (.A1(b[20]), .A2(a[2]), .B1(b[21]), .B2(a[1]), .ZN(n_2803));
   NAND2_X1 i_2130 (.A1(b[22]), .A2(a[0]), .ZN(n_2806));
   OAI21_X1 i_2131 (.A(n_2802), .B1(n_2803), .B2(n_2806), .ZN(n_1901));
   NAND4_X1 i_2132 (.A1(b[18]), .A2(b[17]), .A3(a[5]), .A4(a[4]), .ZN(n_2807));
   AOI22_X1 i_2133 (.A1(b[17]), .A2(a[5]), .B1(b[18]), .B2(a[4]), .ZN(n_2808));
   NAND2_X1 i_2134 (.A1(b[19]), .A2(a[3]), .ZN(n_2809));
   OAI21_X1 i_2135 (.A(n_2807), .B1(n_2808), .B2(n_2809), .ZN(n_1908));
   NAND4_X1 i_2136 (.A1(b[15]), .A2(b[14]), .A3(a[8]), .A4(a[7]), .ZN(n_2810));
   AOI22_X1 i_2137 (.A1(b[14]), .A2(a[8]), .B1(b[15]), .B2(a[7]), .ZN(n_2813));
   NAND2_X1 i_2154 (.A1(b[16]), .A2(a[6]), .ZN(n_2814));
   OAI21_X1 i_2155 (.A(n_2810), .B1(n_2813), .B2(n_2814), .ZN(n_1915));
   NAND4_X1 i_2156 (.A1(a[11]), .A2(b[12]), .A3(b[11]), .A4(a[10]), .ZN(n_2815));
   AOI22_X1 i_2157 (.A1(a[11]), .A2(b[11]), .B1(b[12]), .B2(a[10]), .ZN(n_2816));
   NAND2_X1 i_2158 (.A1(b[13]), .A2(a[9]), .ZN(n_2817));
   OAI21_X1 i_2159 (.A(n_2815), .B1(n_2816), .B2(n_2817), .ZN(n_1922));
   NAND4_X1 i_2160 (.A1(a[14]), .A2(a[13]), .A3(b[9]), .A4(b[8]), .ZN(n_2820));
   AOI22_X1 i_2161 (.A1(a[14]), .A2(b[8]), .B1(a[13]), .B2(b[9]), .ZN(n_2821));
   NAND2_X1 i_2162 (.A1(a[12]), .A2(b[10]), .ZN(n_2822));
   OAI21_X1 i_2163 (.A(n_2820), .B1(n_2821), .B2(n_2822), .ZN(n_1929));
   NAND4_X1 i_2164 (.A1(a[17]), .A2(a[16]), .A3(b[6]), .A4(b[5]), .ZN(n_2823));
   AOI22_X1 i_2165 (.A1(a[17]), .A2(b[5]), .B1(a[16]), .B2(b[6]), .ZN(n_2824));
   NAND2_X1 i_2166 (.A1(a[15]), .A2(b[7]), .ZN(n_2827));
   OAI21_X1 i_2167 (.A(n_2823), .B1(n_2824), .B2(n_2827), .ZN(n_1936));
   NAND4_X1 i_2168 (.A1(a[20]), .A2(a[19]), .A3(b[3]), .A4(b[2]), .ZN(n_2828));
   AOI22_X1 i_2169 (.A1(a[20]), .A2(b[2]), .B1(a[19]), .B2(b[3]), .ZN(n_2829));
   NAND2_X1 i_2170 (.A1(a[18]), .A2(b[4]), .ZN(n_2830));
   OAI21_X1 i_2171 (.A(n_2828), .B1(n_2829), .B2(n_2830), .ZN(n_1943));
   INV_X1 i_2172 (.A(n_2803), .ZN(n_2831));
   NAND2_X1 i_2173 (.A1(n_2831), .A2(n_2802), .ZN(n_2833));
   XOR2_X1 i_2174 (.A(n_2833), .B(n_2806), .Z(n_1900));
   INV_X1 i_2175 (.A(n_2808), .ZN(n_2834));
   NAND2_X1 i_2176 (.A1(n_2834), .A2(n_2807), .ZN(n_2835));
   XOR2_X1 i_2177 (.A(n_2835), .B(n_2809), .Z(n_1907));
   INV_X1 i_2178 (.A(n_2813), .ZN(n_2836));
   NAND2_X1 i_2179 (.A1(n_2836), .A2(n_2810), .ZN(n_2837));
   XOR2_X1 i_2180 (.A(n_2837), .B(n_2814), .Z(n_1914));
   INV_X1 i_2181 (.A(n_2816), .ZN(n_2838));
   NAND2_X1 i_2182 (.A1(n_2838), .A2(n_2815), .ZN(n_2840));
   XOR2_X1 i_2183 (.A(n_2840), .B(n_2817), .Z(n_1921));
   INV_X1 i_2184 (.A(n_2821), .ZN(n_2841));
   NAND2_X1 i_2185 (.A1(n_2841), .A2(n_2820), .ZN(n_2842));
   XOR2_X1 i_2186 (.A(n_2842), .B(n_2822), .Z(n_1928));
   INV_X1 i_2187 (.A(n_2824), .ZN(n_2843));
   NAND2_X1 i_2188 (.A1(n_2843), .A2(n_2823), .ZN(n_2844));
   XOR2_X1 i_2189 (.A(n_2844), .B(n_2827), .Z(n_1935));
   INV_X1 i_2190 (.A(n_2829), .ZN(n_2847));
   NAND2_X1 i_2191 (.A1(n_2847), .A2(n_2828), .ZN(n_2848));
   XOR2_X1 i_2192 (.A(n_2848), .B(n_2830), .Z(n_1942));
   INV_X1 i_2193 (.A(n_2799), .ZN(n_2849));
   NAND2_X1 i_2194 (.A1(n_2849), .A2(n_2801), .ZN(n_2850));
   XOR2_X1 i_2195 (.A(n_2850), .B(n_2800), .Z(n_1948));
   NAND4_X1 i_2196 (.A1(a[17]), .A2(a[16]), .A3(b[3]), .A4(b[4]), .ZN(n_2851));
   AOI22_X1 i_2197 (.A1(a[17]), .A2(b[3]), .B1(a[16]), .B2(b[4]), .ZN(n_2890));
   NAND2_X1 i_2198 (.A1(a[15]), .A2(b[5]), .ZN(n_2891));
   OAI21_X1 i_2199 (.A(n_2851), .B1(n_2890), .B2(n_2891), .ZN(n_2894));
   NAND4_X1 i_2200 (.A1(a[20]), .A2(a[19]), .A3(b[1]), .A4(b[0]), .ZN(n_2895));
   AOI22_X1 i_2201 (.A1(a[20]), .A2(b[0]), .B1(a[19]), .B2(b[1]), .ZN(n_2896));
   NAND2_X1 i_2202 (.A1(a[18]), .A2(b[2]), .ZN(n_2897));
   OAI21_X1 i_2203 (.A(n_2895), .B1(n_2896), .B2(n_2897), .ZN(n_2898));
   NOR2_X1 i_2204 (.A1(n_2894), .A2(n_2898), .ZN(n_2901));
   NAND2_X1 i_2205 (.A1(a[21]), .A2(b[0]), .ZN(n_2902));
   NAND2_X1 i_2206 (.A1(n_2894), .A2(n_2898), .ZN(n_2903));
   AOI21_X1 i_2207 (.A(n_2901), .B1(n_2902), .B2(n_2903), .ZN(n_1869));
   NAND4_X1 i_2208 (.A1(b[20]), .A2(b[19]), .A3(a[2]), .A4(a[1]), .ZN(n_2904));
   AOI22_X1 i_2209 (.A1(b[19]), .A2(a[2]), .B1(b[20]), .B2(a[1]), .ZN(n_2905));
   NAND2_X1 i_2210 (.A1(b[21]), .A2(a[0]), .ZN(n_2908));
   OAI21_X1 i_2211 (.A(n_2904), .B1(n_2905), .B2(n_2908), .ZN(n_1820));
   NAND4_X1 i_2212 (.A1(b[17]), .A2(b[16]), .A3(a[5]), .A4(a[4]), .ZN(n_2909));
   AOI22_X1 i_2213 (.A1(b[16]), .A2(a[5]), .B1(b[17]), .B2(a[4]), .ZN(n_2910));
   NAND2_X1 i_2214 (.A1(b[18]), .A2(a[3]), .ZN(n_2911));
   OAI21_X1 i_2215 (.A(n_2909), .B1(n_2910), .B2(n_2911), .ZN(n_1827));
   NAND4_X1 i_2216 (.A1(b[14]), .A2(b[13]), .A3(a[8]), .A4(a[7]), .ZN(n_2912));
   AOI22_X1 i_2217 (.A1(b[13]), .A2(a[8]), .B1(b[14]), .B2(a[7]), .ZN(n_2915));
   NAND2_X1 i_2218 (.A1(b[15]), .A2(a[6]), .ZN(n_2916));
   OAI21_X1 i_2219 (.A(n_2912), .B1(n_2915), .B2(n_2916), .ZN(n_1834));
   NAND4_X1 i_2220 (.A1(a[11]), .A2(b[11]), .A3(a[10]), .A4(b[10]), .ZN(n_2917));
   AOI22_X1 i_2221 (.A1(a[11]), .A2(b[10]), .B1(b[11]), .B2(a[10]), .ZN(n_2918));
   NAND2_X1 i_2222 (.A1(b[12]), .A2(a[9]), .ZN(n_2919));
   OAI21_X1 i_2223 (.A(n_2917), .B1(n_2918), .B2(n_2919), .ZN(n_1841));
   NAND4_X1 i_2224 (.A1(a[14]), .A2(a[13]), .A3(b[8]), .A4(b[7]), .ZN(n_2922));
   AOI22_X1 i_2241 (.A1(a[14]), .A2(b[7]), .B1(a[13]), .B2(b[8]), .ZN(n_2923));
   NAND2_X1 i_2242 (.A1(a[12]), .A2(b[9]), .ZN(n_2924));
   OAI21_X1 i_2243 (.A(n_2922), .B1(n_2923), .B2(n_2924), .ZN(n_1848));
   NAND4_X1 i_2244 (.A1(a[17]), .A2(a[16]), .A3(b[4]), .A4(b[5]), .ZN(n_2925));
   AOI22_X1 i_2245 (.A1(a[17]), .A2(b[4]), .B1(a[16]), .B2(b[5]), .ZN(n_2926));
   NAND2_X1 i_2246 (.A1(a[15]), .A2(b[6]), .ZN(n_2929));
   OAI21_X1 i_2247 (.A(n_2925), .B1(n_2926), .B2(n_2929), .ZN(n_1855));
   INV_X1 i_2248 (.A(n_2901), .ZN(n_2930));
   NAND2_X1 i_2249 (.A1(n_2930), .A2(n_2903), .ZN(n_2931));
   XOR2_X1 i_2250 (.A(n_2931), .B(n_2902), .Z(n_1868));
   INV_X1 i_2251 (.A(n_2905), .ZN(n_2932));
   NAND2_X1 i_2252 (.A1(n_2932), .A2(n_2904), .ZN(n_2933));
   XOR2_X1 i_2253 (.A(n_2933), .B(n_2908), .Z(n_1819));
   INV_X1 i_2254 (.A(n_2910), .ZN(n_2936));
   NAND2_X1 i_2255 (.A1(n_2936), .A2(n_2909), .ZN(n_2937));
   XOR2_X1 i_2256 (.A(n_2937), .B(n_2911), .Z(n_1826));
   INV_X1 i_2257 (.A(n_2915), .ZN(n_2938));
   NAND2_X1 i_2258 (.A1(n_2938), .A2(n_2912), .ZN(n_2939));
   XOR2_X1 i_2259 (.A(n_2939), .B(n_2916), .Z(n_1833));
   INV_X1 i_2260 (.A(n_2918), .ZN(n_2940));
   NAND2_X1 i_2261 (.A1(n_2940), .A2(n_2917), .ZN(n_2943));
   XOR2_X1 i_2262 (.A(n_2943), .B(n_2919), .Z(n_1840));
   INV_X1 i_2263 (.A(n_2923), .ZN(n_2944));
   NAND2_X1 i_2264 (.A1(n_2944), .A2(n_2922), .ZN(n_2945));
   XOR2_X1 i_2265 (.A(n_2945), .B(n_2924), .Z(n_1847));
   INV_X1 i_2266 (.A(n_2926), .ZN(n_2946));
   NAND2_X1 i_2267 (.A1(n_2946), .A2(n_2925), .ZN(n_2947));
   XOR2_X1 i_2268 (.A(n_2947), .B(n_2929), .Z(n_1854));
   INV_X1 i_2269 (.A(n_2794), .ZN(n_2950));
   NAND2_X1 i_2270 (.A1(n_2950), .A2(n_2793), .ZN(n_2951));
   XOR2_X1 i_2271 (.A(n_2951), .B(n_2795), .Z(n_1861));
   NAND4_X1 i_2272 (.A1(b[19]), .A2(b[18]), .A3(a[2]), .A4(a[1]), .ZN(n_2952));
   AOI22_X1 i_2273 (.A1(b[18]), .A2(a[2]), .B1(b[19]), .B2(a[1]), .ZN(n_2953));
   NAND2_X1 i_2274 (.A1(b[20]), .A2(a[0]), .ZN(n_2954));
   OAI21_X1 i_2275 (.A(n_2952), .B1(n_2953), .B2(n_2954), .ZN(n_1747));
   NAND4_X1 i_2276 (.A1(b[16]), .A2(b[15]), .A3(a[5]), .A4(a[4]), .ZN(n_2957));
   AOI22_X1 i_2277 (.A1(b[15]), .A2(a[5]), .B1(b[16]), .B2(a[4]), .ZN(n_2958));
   NAND2_X1 i_2278 (.A1(b[17]), .A2(a[3]), .ZN(n_2959));
   OAI21_X1 i_2279 (.A(n_2957), .B1(n_2958), .B2(n_2959), .ZN(n_1754));
   NAND4_X1 i_2280 (.A1(b[13]), .A2(b[12]), .A3(a[8]), .A4(a[7]), .ZN(n_2960));
   AOI22_X1 i_2281 (.A1(b[12]), .A2(a[8]), .B1(b[13]), .B2(a[7]), .ZN(n_2961));
   NAND2_X1 i_2282 (.A1(b[14]), .A2(a[6]), .ZN(n_2964));
   OAI21_X1 i_2283 (.A(n_2960), .B1(n_2961), .B2(n_2964), .ZN(n_1761));
   NAND4_X1 i_2284 (.A1(a[11]), .A2(a[10]), .A3(b[10]), .A4(b[9]), .ZN(n_2965));
   AOI22_X1 i_2285 (.A1(a[11]), .A2(b[9]), .B1(a[10]), .B2(b[10]), .ZN(n_2966));
   NAND2_X1 i_2286 (.A1(b[11]), .A2(a[9]), .ZN(n_2967));
   OAI21_X1 i_2287 (.A(n_2965), .B1(n_2966), .B2(n_2967), .ZN(n_1768));
   NAND4_X1 i_2288 (.A1(a[14]), .A2(a[13]), .A3(b[7]), .A4(b[6]), .ZN(n_3006));
   AOI22_X1 i_2289 (.A1(a[14]), .A2(b[6]), .B1(a[13]), .B2(b[7]), .ZN(n_3007));
   NAND2_X1 i_2290 (.A1(a[12]), .A2(b[8]), .ZN(n_3010));
   OAI21_X1 i_2291 (.A(n_3006), .B1(n_3007), .B2(n_3010), .ZN(n_1775));
   INV_X1 i_2292 (.A(n_2953), .ZN(n_3011));
   NAND2_X1 i_2293 (.A1(n_3011), .A2(n_2952), .ZN(n_3012));
   XOR2_X1 i_2294 (.A(n_3012), .B(n_2954), .Z(n_1746));
   INV_X1 i_2295 (.A(n_2958), .ZN(n_3013));
   NAND2_X1 i_2296 (.A1(n_3013), .A2(n_2957), .ZN(n_3014));
   XOR2_X1 i_2297 (.A(n_3014), .B(n_2959), .Z(n_1753));
   INV_X1 i_2298 (.A(n_2961), .ZN(n_3017));
   NAND2_X1 i_2299 (.A1(n_3017), .A2(n_2960), .ZN(n_3018));
   XOR2_X1 i_2300 (.A(n_3018), .B(n_2964), .Z(n_1760));
   INV_X1 i_2301 (.A(n_2966), .ZN(n_3019));
   NAND2_X1 i_2302 (.A1(n_3019), .A2(n_2965), .ZN(n_3020));
   XOR2_X1 i_2303 (.A(n_3020), .B(n_2967), .Z(n_1767));
   INV_X1 i_2304 (.A(n_3007), .ZN(n_3021));
   NAND2_X1 i_2305 (.A1(n_3021), .A2(n_3006), .ZN(n_3024));
   XOR2_X1 i_2306 (.A(n_3024), .B(n_3010), .Z(n_1774));
   INV_X1 i_2307 (.A(n_2890), .ZN(n_3025));
   NAND2_X1 i_2308 (.A1(n_3025), .A2(n_2851), .ZN(n_3026));
   XOR2_X1 i_2309 (.A(n_3026), .B(n_2891), .Z(n_1781));
   INV_X1 i_2310 (.A(n_2896), .ZN(n_3027));
   NAND2_X1 i_2311 (.A1(n_3027), .A2(n_2895), .ZN(n_3028));
   XOR2_X1 i_2329 (.A(n_3028), .B(n_2897), .Z(n_1788));
   NAND4_X1 i_2330 (.A1(a[17]), .A2(a[16]), .A3(b[2]), .A4(b[1]), .ZN(n_3031));
   AOI22_X1 i_2331 (.A1(a[17]), .A2(b[1]), .B1(a[16]), .B2(b[2]), .ZN(n_3032));
   NAND2_X1 i_2332 (.A1(a[15]), .A2(b[3]), .ZN(n_3033));
   OAI21_X1 i_2333 (.A(n_3031), .B1(n_3032), .B2(n_3033), .ZN(n_3034));
   AOI21_X1 i_2334 (.A(n_3034), .B1(a[19]), .B2(b[0]), .ZN(n_3035));
   NAND2_X1 i_2335 (.A1(a[18]), .A2(b[1]), .ZN(n_3038));
   NAND3_X1 i_2336 (.A1(n_3034), .A2(a[19]), .A3(b[0]), .ZN(n_3039));
   AOI21_X1 i_2337 (.A(n_3035), .B1(n_3038), .B2(n_3039), .ZN(n_1716));
   NAND4_X1 i_2338 (.A1(b[18]), .A2(b[17]), .A3(a[2]), .A4(a[1]), .ZN(n_3040));
   AOI22_X1 i_2339 (.A1(b[17]), .A2(a[2]), .B1(b[18]), .B2(a[1]), .ZN(n_3041));
   NAND2_X1 i_2340 (.A1(b[19]), .A2(a[0]), .ZN(n_3042));
   OAI21_X1 i_2341 (.A(n_3040), .B1(n_3041), .B2(n_3042), .ZN(n_1675));
   NAND4_X1 i_2342 (.A1(b[15]), .A2(b[14]), .A3(a[5]), .A4(a[4]), .ZN(n_3045));
   AOI22_X1 i_2343 (.A1(b[14]), .A2(a[5]), .B1(b[15]), .B2(a[4]), .ZN(n_3046));
   NAND2_X1 i_2344 (.A1(b[16]), .A2(a[3]), .ZN(n_3047));
   OAI21_X1 i_2345 (.A(n_3045), .B1(n_3046), .B2(n_3047), .ZN(n_1682));
   NAND4_X1 i_2346 (.A1(b[12]), .A2(b[11]), .A3(a[8]), .A4(a[7]), .ZN(n_3048));
   AOI22_X1 i_2347 (.A1(b[11]), .A2(a[8]), .B1(b[12]), .B2(a[7]), .ZN(n_3049));
   NAND2_X1 i_2348 (.A1(b[13]), .A2(a[6]), .ZN(n_3052));
   OAI21_X1 i_2349 (.A(n_3048), .B1(n_3049), .B2(n_3052), .ZN(n_1689));
   NAND4_X1 i_2350 (.A1(a[11]), .A2(a[10]), .A3(b[9]), .A4(b[8]), .ZN(n_3053));
   AOI22_X1 i_2351 (.A1(a[11]), .A2(b[8]), .B1(a[10]), .B2(b[9]), .ZN(n_3054));
   NAND2_X1 i_2352 (.A1(b[10]), .A2(a[9]), .ZN(n_3055));
   OAI21_X1 i_2353 (.A(n_3053), .B1(n_3054), .B2(n_3055), .ZN(n_1696));
   NAND4_X1 i_2354 (.A1(a[14]), .A2(a[13]), .A3(b[6]), .A4(b[5]), .ZN(n_3056));
   AOI22_X1 i_2355 (.A1(a[14]), .A2(b[5]), .B1(a[13]), .B2(b[6]), .ZN(n_3059));
   NAND2_X1 i_2356 (.A1(a[12]), .A2(b[7]), .ZN(n_3060));
   OAI21_X1 i_2357 (.A(n_3056), .B1(n_3059), .B2(n_3060), .ZN(n_1703));
   NAND4_X1 i_2358 (.A1(a[17]), .A2(a[16]), .A3(b[3]), .A4(b[2]), .ZN(n_3061));
   AOI22_X1 i_2359 (.A1(a[17]), .A2(b[2]), .B1(a[16]), .B2(b[3]), .ZN(n_3062));
   NAND2_X1 i_2360 (.A1(a[15]), .A2(b[4]), .ZN(n_3063));
   OAI21_X1 i_2361 (.A(n_3061), .B1(n_3062), .B2(n_3063), .ZN(n_1710));
   INV_X1 i_2362 (.A(n_3041), .ZN(n_3066));
   NAND2_X1 i_2363 (.A1(n_3066), .A2(n_3040), .ZN(n_3067));
   XOR2_X1 i_2364 (.A(n_3067), .B(n_3042), .Z(n_1674));
   INV_X1 i_2365 (.A(n_3046), .ZN(n_3068));
   NAND2_X1 i_2366 (.A1(n_3068), .A2(n_3045), .ZN(n_3069));
   XOR2_X1 i_2367 (.A(n_3069), .B(n_3047), .Z(n_1681));
   INV_X1 i_2368 (.A(n_3049), .ZN(n_3070));
   NAND2_X1 i_2369 (.A1(n_3070), .A2(n_3048), .ZN(n_3072));
   XOR2_X1 i_2370 (.A(n_3072), .B(n_3052), .Z(n_1688));
   INV_X1 i_2371 (.A(n_3054), .ZN(n_3073));
   NAND2_X1 i_2372 (.A1(n_3073), .A2(n_3053), .ZN(n_3074));
   XOR2_X1 i_2373 (.A(n_3074), .B(n_3055), .Z(n_1695));
   INV_X1 i_2374 (.A(n_3059), .ZN(n_3075));
   NAND2_X1 i_2375 (.A1(n_3075), .A2(n_3056), .ZN(n_3114));
   XOR2_X1 i_2376 (.A(n_3114), .B(n_3060), .Z(n_1702));
   INV_X1 i_2377 (.A(n_3062), .ZN(n_3115));
   NAND2_X1 i_2378 (.A1(n_3115), .A2(n_3061), .ZN(n_3118));
   XOR2_X1 i_2379 (.A(n_3118), .B(n_3063), .Z(n_1709));
   INV_X1 i_2380 (.A(n_3035), .ZN(n_3119));
   NAND2_X1 i_2381 (.A1(n_3119), .A2(n_3039), .ZN(n_3120));
   XOR2_X1 i_2382 (.A(n_3120), .B(n_3038), .Z(n_1715));
   NAND4_X1 i_2383 (.A1(a[14]), .A2(a[13]), .A3(b[3]), .A4(b[4]), .ZN(n_3121));
   AOI22_X1 i_2384 (.A1(a[14]), .A2(b[3]), .B1(a[13]), .B2(b[4]), .ZN(n_3122));
   NAND2_X1 i_2385 (.A1(a[12]), .A2(b[5]), .ZN(n_3125));
   OAI21_X1 i_2386 (.A(n_3121), .B1(n_3122), .B2(n_3125), .ZN(n_3126));
   NAND4_X1 i_2387 (.A1(a[17]), .A2(a[16]), .A3(b[1]), .A4(b[0]), .ZN(n_3127));
   AOI22_X1 i_2388 (.A1(a[17]), .A2(b[0]), .B1(a[16]), .B2(b[1]), .ZN(n_3128));
   NAND2_X1 i_2389 (.A1(a[15]), .A2(b[2]), .ZN(n_3129));
   OAI21_X1 i_2390 (.A(n_3127), .B1(n_3128), .B2(n_3129), .ZN(n_3132));
   NOR2_X1 i_2391 (.A1(n_3126), .A2(n_3132), .ZN(n_3133));
   NAND2_X1 i_2392 (.A1(a[18]), .A2(b[0]), .ZN(n_3134));
   NAND2_X1 i_2393 (.A1(n_3126), .A2(n_3132), .ZN(n_3135));
   AOI21_X1 i_2394 (.A(n_3133), .B1(n_3134), .B2(n_3135), .ZN(n_1647));
   NAND4_X1 i_2395 (.A1(b[17]), .A2(b[16]), .A3(a[2]), .A4(a[1]), .ZN(n_3136));
   AOI22_X1 i_2396 (.A1(b[16]), .A2(a[2]), .B1(b[17]), .B2(a[1]), .ZN(n_3139));
   NAND2_X1 i_2397 (.A1(b[18]), .A2(a[0]), .ZN(n_3140));
   OAI21_X1 i_2398 (.A(n_3136), .B1(n_3139), .B2(n_3140), .ZN(n_1605));
   NAND4_X1 i_2417 (.A1(b[14]), .A2(b[13]), .A3(a[5]), .A4(a[4]), .ZN(n_3141));
   AOI22_X1 i_2418 (.A1(b[13]), .A2(a[5]), .B1(b[14]), .B2(a[4]), .ZN(n_3142));
   NAND2_X1 i_2419 (.A1(b[15]), .A2(a[3]), .ZN(n_3143));
   OAI21_X1 i_2420 (.A(n_3141), .B1(n_3142), .B2(n_3143), .ZN(n_1612));
   NAND4_X1 i_2421 (.A1(b[11]), .A2(b[10]), .A3(a[8]), .A4(a[7]), .ZN(n_3146));
   AOI22_X1 i_2422 (.A1(b[10]), .A2(a[8]), .B1(b[11]), .B2(a[7]), .ZN(n_3147));
   NAND2_X1 i_2423 (.A1(b[12]), .A2(a[6]), .ZN(n_3148));
   OAI21_X1 i_2424 (.A(n_3146), .B1(n_3147), .B2(n_3148), .ZN(n_1619));
   NAND4_X1 i_2425 (.A1(a[11]), .A2(a[10]), .A3(b[8]), .A4(b[7]), .ZN(n_3149));
   AOI22_X1 i_2426 (.A1(a[11]), .A2(b[7]), .B1(a[10]), .B2(b[8]), .ZN(n_3150));
   NAND2_X1 i_2427 (.A1(a[9]), .A2(b[9]), .ZN(n_3153));
   OAI21_X1 i_2428 (.A(n_3149), .B1(n_3150), .B2(n_3153), .ZN(n_1626));
   NAND4_X1 i_2429 (.A1(a[14]), .A2(a[13]), .A3(b[4]), .A4(b[5]), .ZN(n_3154));
   AOI22_X1 i_2430 (.A1(a[14]), .A2(b[4]), .B1(a[13]), .B2(b[5]), .ZN(n_3155));
   NAND2_X1 i_2431 (.A1(a[12]), .A2(b[6]), .ZN(n_3156));
   OAI21_X1 i_2432 (.A(n_3154), .B1(n_3155), .B2(n_3156), .ZN(n_1633));
   INV_X1 i_2433 (.A(n_3133), .ZN(n_3157));
   NAND2_X1 i_2434 (.A1(n_3157), .A2(n_3135), .ZN(n_3160));
   XOR2_X1 i_2435 (.A(n_3160), .B(n_3134), .Z(n_1646));
   INV_X1 i_2436 (.A(n_3139), .ZN(n_3161));
   NAND2_X1 i_2437 (.A1(n_3161), .A2(n_3136), .ZN(n_3162));
   XOR2_X1 i_2438 (.A(n_3162), .B(n_3140), .Z(n_1604));
   INV_X1 i_2439 (.A(n_3142), .ZN(n_3163));
   NAND2_X1 i_2440 (.A1(n_3163), .A2(n_3141), .ZN(n_3164));
   XOR2_X1 i_2441 (.A(n_3164), .B(n_3143), .Z(n_1611));
   INV_X1 i_2442 (.A(n_3147), .ZN(n_3166));
   NAND2_X1 i_2443 (.A1(n_3166), .A2(n_3146), .ZN(n_3167));
   XOR2_X1 i_2444 (.A(n_3167), .B(n_3148), .Z(n_1618));
   INV_X1 i_2445 (.A(n_3150), .ZN(n_3168));
   NAND2_X1 i_2446 (.A1(n_3168), .A2(n_3149), .ZN(n_3169));
   XOR2_X1 i_2447 (.A(n_3169), .B(n_3153), .Z(n_1625));
   INV_X1 i_2448 (.A(n_3155), .ZN(n_3170));
   NAND2_X1 i_2449 (.A1(n_3170), .A2(n_3154), .ZN(n_3171));
   XOR2_X1 i_2450 (.A(n_3171), .B(n_3156), .Z(n_1632));
   INV_X1 i_2451 (.A(n_3032), .ZN(n_3173));
   NAND2_X1 i_2452 (.A1(n_3173), .A2(n_3031), .ZN(n_3174));
   XOR2_X1 i_2453 (.A(n_3174), .B(n_3033), .Z(n_1639));
   NAND4_X1 i_2454 (.A1(b[16]), .A2(b[15]), .A3(a[2]), .A4(a[1]), .ZN(n_3175));
   AOI22_X1 i_2455 (.A1(b[15]), .A2(a[2]), .B1(b[16]), .B2(a[1]), .ZN(n_3176));
   NAND2_X1 i_2456 (.A1(b[17]), .A2(a[0]), .ZN(n_3177));
   OAI21_X1 i_2457 (.A(n_3175), .B1(n_3176), .B2(n_3177), .ZN(n_1543));
   NAND4_X1 i_2458 (.A1(b[13]), .A2(b[12]), .A3(a[5]), .A4(a[4]), .ZN(n_3180));
   AOI22_X1 i_2459 (.A1(b[12]), .A2(a[5]), .B1(b[13]), .B2(a[4]), .ZN(n_3181));
   NAND2_X1 i_2460 (.A1(b[14]), .A2(a[3]), .ZN(n_3182));
   OAI21_X1 i_2461 (.A(n_3180), .B1(n_3181), .B2(n_3182), .ZN(n_1550));
   NAND4_X1 i_2462 (.A1(b[10]), .A2(a[8]), .A3(b[9]), .A4(a[7]), .ZN(n_3183));
   AOI22_X1 i_2463 (.A1(a[8]), .A2(b[9]), .B1(b[10]), .B2(a[7]), .ZN(n_3184));
   NAND2_X1 i_2464 (.A1(b[11]), .A2(a[6]), .ZN(n_3221));
   OAI21_X1 i_2465 (.A(n_3183), .B1(n_3184), .B2(n_3221), .ZN(n_1557));
   NAND4_X1 i_2466 (.A1(a[11]), .A2(a[10]), .A3(b[7]), .A4(b[6]), .ZN(n_3222));
   AOI22_X1 i_2467 (.A1(a[11]), .A2(b[6]), .B1(a[10]), .B2(b[7]), .ZN(n_3225));
   NAND2_X1 i_2468 (.A1(a[9]), .A2(b[8]), .ZN(n_3226));
   OAI21_X1 i_2469 (.A(n_3222), .B1(n_3225), .B2(n_3226), .ZN(n_1564));
   INV_X1 i_2470 (.A(n_3176), .ZN(n_3227));
   NAND2_X1 i_2471 (.A1(n_3227), .A2(n_3175), .ZN(n_3228));
   XOR2_X1 i_2472 (.A(n_3228), .B(n_3177), .Z(n_1542));
   INV_X1 i_2473 (.A(n_3181), .ZN(n_3229));
   NAND2_X1 i_2474 (.A1(n_3229), .A2(n_3180), .ZN(n_3232));
   XOR2_X1 i_2475 (.A(n_3232), .B(n_3182), .Z(n_1549));
   INV_X1 i_2476 (.A(n_3184), .ZN(n_3233));
   NAND2_X1 i_2477 (.A1(n_3233), .A2(n_3183), .ZN(n_3234));
   XOR2_X1 i_2478 (.A(n_3234), .B(n_3221), .Z(n_1556));
   INV_X1 i_2479 (.A(n_3225), .ZN(n_3235));
   NAND2_X1 i_2480 (.A1(n_3235), .A2(n_3222), .ZN(n_3236));
   XOR2_X1 i_2481 (.A(n_3236), .B(n_3226), .Z(n_1563));
   INV_X1 i_2482 (.A(n_3122), .ZN(n_3239));
   NAND2_X1 i_2483 (.A1(n_3239), .A2(n_3121), .ZN(n_3240));
   XOR2_X1 i_2484 (.A(n_3240), .B(n_3125), .Z(n_1570));
   INV_X1 i_2485 (.A(n_3128), .ZN(n_3241));
   NAND2_X1 i_2486 (.A1(n_3241), .A2(n_3127), .ZN(n_3242));
   XOR2_X1 i_2487 (.A(n_3242), .B(n_3129), .Z(n_1577));
   NAND4_X1 i_2488 (.A1(a[14]), .A2(a[13]), .A3(b[2]), .A4(b[1]), .ZN(n_3243));
   AOI22_X1 i_2489 (.A1(a[14]), .A2(b[1]), .B1(a[13]), .B2(b[2]), .ZN(n_3246));
   NAND2_X1 i_2490 (.A1(a[12]), .A2(b[3]), .ZN(n_3247));
   OAI21_X1 i_2491 (.A(n_3243), .B1(n_3246), .B2(n_3247), .ZN(n_3248));
   AOI21_X1 i_2492 (.A(n_3248), .B1(a[16]), .B2(b[0]), .ZN(n_3249));
   NAND2_X1 i_2493 (.A1(a[15]), .A2(b[1]), .ZN(n_3250));
   NAND3_X1 i_2494 (.A1(n_3248), .A2(a[16]), .A3(b[0]), .ZN(n_3253));
   AOI21_X1 i_2513 (.A(n_3249), .B1(n_3250), .B2(n_3253), .ZN(n_1516));
   NAND4_X1 i_2514 (.A1(b[15]), .A2(b[14]), .A3(a[2]), .A4(a[1]), .ZN(n_3254));
   AOI22_X1 i_2515 (.A1(b[14]), .A2(a[2]), .B1(b[15]), .B2(a[1]), .ZN(n_3255));
   NAND2_X1 i_2516 (.A1(b[16]), .A2(a[0]), .ZN(n_3256));
   OAI21_X1 i_2517 (.A(n_3254), .B1(n_3255), .B2(n_3256), .ZN(n_1482));
   NAND4_X1 i_2518 (.A1(b[12]), .A2(b[11]), .A3(a[5]), .A4(a[4]), .ZN(n_3257));
   AOI22_X1 i_2519 (.A1(b[11]), .A2(a[5]), .B1(b[12]), .B2(a[4]), .ZN(n_3260));
   NAND2_X1 i_2520 (.A1(b[13]), .A2(a[3]), .ZN(n_3261));
   OAI21_X1 i_2521 (.A(n_3257), .B1(n_3260), .B2(n_3261), .ZN(n_1489));
   NAND4_X1 i_2522 (.A1(a[8]), .A2(b[9]), .A3(b[8]), .A4(a[7]), .ZN(n_3262));
   AOI22_X1 i_2523 (.A1(a[8]), .A2(b[8]), .B1(b[9]), .B2(a[7]), .ZN(n_3263));
   NAND2_X1 i_2524 (.A1(b[10]), .A2(a[6]), .ZN(n_3264));
   OAI21_X1 i_2525 (.A(n_3262), .B1(n_3263), .B2(n_3264), .ZN(n_1496));
   NAND4_X1 i_2526 (.A1(a[11]), .A2(a[10]), .A3(b[6]), .A4(b[5]), .ZN(n_3267));
   AOI22_X1 i_2527 (.A1(a[11]), .A2(b[5]), .B1(a[10]), .B2(b[6]), .ZN(n_3268));
   NAND2_X1 i_2528 (.A1(a[9]), .A2(b[7]), .ZN(n_3269));
   OAI21_X1 i_2529 (.A(n_3267), .B1(n_3268), .B2(n_3269), .ZN(n_1503));
   NAND4_X1 i_2530 (.A1(a[14]), .A2(a[13]), .A3(b[3]), .A4(b[2]), .ZN(n_3270));
   AOI22_X1 i_2531 (.A1(a[14]), .A2(b[2]), .B1(a[13]), .B2(b[3]), .ZN(n_3271));
   NAND2_X1 i_2532 (.A1(a[12]), .A2(b[4]), .ZN(n_3274));
   OAI21_X1 i_2533 (.A(n_3270), .B1(n_3271), .B2(n_3274), .ZN(n_1510));
   INV_X1 i_2534 (.A(n_3255), .ZN(n_3275));
   NAND2_X1 i_2535 (.A1(n_3275), .A2(n_3254), .ZN(n_3276));
   XOR2_X1 i_2536 (.A(n_3276), .B(n_3256), .Z(n_1481));
   INV_X1 i_2537 (.A(n_3260), .ZN(n_3277));
   NAND2_X1 i_2538 (.A1(n_3277), .A2(n_3257), .ZN(n_3278));
   XOR2_X1 i_2539 (.A(n_3278), .B(n_3261), .Z(n_1488));
   INV_X1 i_2540 (.A(n_3263), .ZN(n_3281));
   NAND2_X1 i_2541 (.A1(n_3281), .A2(n_3262), .ZN(n_3282));
   XOR2_X1 i_2542 (.A(n_3282), .B(n_3264), .Z(n_1495));
   INV_X1 i_2543 (.A(n_3268), .ZN(n_3283));
   NAND2_X1 i_2544 (.A1(n_3283), .A2(n_3267), .ZN(n_3284));
   XOR2_X1 i_2545 (.A(n_3284), .B(n_3269), .Z(n_1502));
   INV_X1 i_2546 (.A(n_3271), .ZN(n_3285));
   NAND2_X1 i_2547 (.A1(n_3285), .A2(n_3270), .ZN(n_3288));
   XOR2_X1 i_2548 (.A(n_3288), .B(n_3274), .Z(n_1509));
   INV_X1 i_2549 (.A(n_3249), .ZN(n_3289));
   NAND2_X1 i_2550 (.A1(n_3289), .A2(n_3253), .ZN(n_3290));
   XOR2_X1 i_2551 (.A(n_3290), .B(n_3250), .Z(n_1515));
   NAND4_X1 i_2552 (.A1(a[11]), .A2(a[10]), .A3(b[3]), .A4(b[4]), .ZN(n_3291));
   AOI22_X1 i_2553 (.A1(a[11]), .A2(b[3]), .B1(a[10]), .B2(b[4]), .ZN(n_3326));
   NAND2_X1 i_2554 (.A1(a[9]), .A2(b[5]), .ZN(n_3327));
   OAI21_X1 i_2555 (.A(n_3291), .B1(n_3326), .B2(n_3327), .ZN(n_3330));
   NAND4_X1 i_2556 (.A1(a[14]), .A2(a[13]), .A3(b[1]), .A4(b[0]), .ZN(n_3331));
   AOI22_X1 i_2557 (.A1(a[14]), .A2(b[0]), .B1(a[13]), .B2(b[1]), .ZN(n_3332));
   NAND2_X1 i_2558 (.A1(a[12]), .A2(b[2]), .ZN(n_3333));
   OAI21_X1 i_2559 (.A(n_3331), .B1(n_3332), .B2(n_3333), .ZN(n_3334));
   NOR2_X1 i_2560 (.A1(n_3330), .A2(n_3334), .ZN(n_3337));
   NAND2_X1 i_2561 (.A1(a[15]), .A2(b[0]), .ZN(n_3338));
   NAND2_X1 i_2562 (.A1(n_3330), .A2(n_3334), .ZN(n_3339));
   AOI21_X1 i_2563 (.A(n_3337), .B1(n_3338), .B2(n_3339), .ZN(n_1458));
   NAND4_X1 i_2564 (.A1(b[14]), .A2(b[13]), .A3(a[2]), .A4(a[1]), .ZN(n_3340));
   AOI22_X1 i_2565 (.A1(b[13]), .A2(a[2]), .B1(b[14]), .B2(a[1]), .ZN(n_3341));
   NAND2_X1 i_2566 (.A1(b[15]), .A2(a[0]), .ZN(n_3344));
   OAI21_X1 i_2567 (.A(n_3340), .B1(n_3341), .B2(n_3344), .ZN(n_1423));
   NAND4_X1 i_2568 (.A1(b[11]), .A2(b[10]), .A3(a[5]), .A4(a[4]), .ZN(n_3345));
   AOI22_X1 i_2569 (.A1(b[10]), .A2(a[5]), .B1(b[11]), .B2(a[4]), .ZN(n_3346));
   NAND2_X1 i_2570 (.A1(b[12]), .A2(a[3]), .ZN(n_3347));
   OAI21_X1 i_2571 (.A(n_3345), .B1(n_3346), .B2(n_3347), .ZN(n_1430));
   NAND4_X1 i_2572 (.A1(a[8]), .A2(b[8]), .A3(a[7]), .A4(b[7]), .ZN(n_3348));
   AOI22_X1 i_2573 (.A1(a[8]), .A2(b[7]), .B1(b[8]), .B2(a[7]), .ZN(n_3351));
   NAND2_X1 i_2574 (.A1(b[9]), .A2(a[6]), .ZN(n_3352));
   OAI21_X1 i_2575 (.A(n_3348), .B1(n_3351), .B2(n_3352), .ZN(n_1437));
   NAND4_X1 i_2576 (.A1(a[11]), .A2(a[10]), .A3(b[4]), .A4(b[5]), .ZN(n_3353));
   AOI22_X1 i_2577 (.A1(a[11]), .A2(b[4]), .B1(a[10]), .B2(b[5]), .ZN(n_3354));
   NAND2_X1 i_2578 (.A1(a[9]), .A2(b[6]), .ZN(n_3355));
   OAI21_X1 i_2579 (.A(n_3353), .B1(n_3354), .B2(n_3355), .ZN(n_1444));
   INV_X1 i_2580 (.A(n_3337), .ZN(n_3358));
   NAND2_X1 i_2581 (.A1(n_3358), .A2(n_3339), .ZN(n_3359));
   XOR2_X1 i_2582 (.A(n_3359), .B(n_3338), .Z(n_1457));
   INV_X1 i_2583 (.A(n_3341), .ZN(n_3360));
   NAND2_X1 i_2584 (.A1(n_3360), .A2(n_3340), .ZN(n_3361));
   XOR2_X1 i_2585 (.A(n_3361), .B(n_3344), .Z(n_1422));
   INV_X1 i_2586 (.A(n_3346), .ZN(n_3362));
   NAND2_X1 i_2587 (.A1(n_3362), .A2(n_3345), .ZN(n_3365));
   XOR2_X1 i_2588 (.A(n_3365), .B(n_3347), .Z(n_1429));
   INV_X1 i_2589 (.A(n_3351), .ZN(n_3366));
   NAND2_X1 i_2590 (.A1(n_3366), .A2(n_3348), .ZN(n_3367));
   XOR2_X1 i_2610 (.A(n_3367), .B(n_3352), .Z(n_1436));
   INV_X1 i_2611 (.A(n_3354), .ZN(n_3368));
   NAND2_X1 i_2612 (.A1(n_3368), .A2(n_3353), .ZN(n_3369));
   XOR2_X1 i_2613 (.A(n_3369), .B(n_3355), .Z(n_1443));
   INV_X1 i_2614 (.A(n_3246), .ZN(n_3372));
   NAND2_X1 i_2615 (.A1(n_3372), .A2(n_3243), .ZN(n_3373));
   XOR2_X1 i_2616 (.A(n_3373), .B(n_3247), .Z(n_1450));
   NAND4_X1 i_2617 (.A1(b[13]), .A2(b[12]), .A3(a[2]), .A4(a[1]), .ZN(n_3374));
   AOI22_X1 i_2618 (.A1(b[12]), .A2(a[2]), .B1(b[13]), .B2(a[1]), .ZN(n_3375));
   NAND2_X1 i_2619 (.A1(b[14]), .A2(a[0]), .ZN(n_3376));
   OAI21_X1 i_2620 (.A(n_3374), .B1(n_3375), .B2(n_3376), .ZN(n_1372));
   NAND4_X1 i_2621 (.A1(b[10]), .A2(b[9]), .A3(a[5]), .A4(a[4]), .ZN(n_3379));
   AOI22_X1 i_2622 (.A1(b[9]), .A2(a[5]), .B1(b[10]), .B2(a[4]), .ZN(n_3380));
   NAND2_X1 i_2623 (.A1(b[11]), .A2(a[3]), .ZN(n_3381));
   OAI21_X1 i_2624 (.A(n_3379), .B1(n_3380), .B2(n_3381), .ZN(n_1379));
   NAND4_X1 i_2625 (.A1(a[8]), .A2(a[7]), .A3(b[7]), .A4(b[6]), .ZN(n_3382));
   AOI22_X1 i_2626 (.A1(a[8]), .A2(b[6]), .B1(a[7]), .B2(b[7]), .ZN(n_3383));
   NAND2_X1 i_2627 (.A1(b[8]), .A2(a[6]), .ZN(n_3385));
   OAI21_X1 i_2628 (.A(n_3382), .B1(n_3383), .B2(n_3385), .ZN(n_1386));
   INV_X1 i_2629 (.A(n_3375), .ZN(n_3386));
   NAND2_X1 i_2630 (.A1(n_3386), .A2(n_3374), .ZN(n_3387));
   XOR2_X1 i_2631 (.A(n_3387), .B(n_3376), .Z(n_1371));
   INV_X1 i_2632 (.A(n_3380), .ZN(n_3388));
   NAND2_X1 i_2633 (.A1(n_3388), .A2(n_3379), .ZN(n_3423));
   XOR2_X1 i_2634 (.A(n_3423), .B(n_3381), .Z(n_1378));
   INV_X1 i_2635 (.A(n_3383), .ZN(n_3424));
   NAND2_X1 i_2636 (.A1(n_3424), .A2(n_3382), .ZN(n_3427));
   XOR2_X1 i_2637 (.A(n_3427), .B(n_3385), .Z(n_1385));
   INV_X1 i_2638 (.A(n_3326), .ZN(n_3428));
   NAND2_X1 i_2639 (.A1(n_3428), .A2(n_3291), .ZN(n_3429));
   XOR2_X1 i_2640 (.A(n_3429), .B(n_3327), .Z(n_1392));
   INV_X1 i_2641 (.A(n_3332), .ZN(n_3430));
   NAND2_X1 i_2642 (.A1(n_3430), .A2(n_3331), .ZN(n_3431));
   XOR2_X1 i_2643 (.A(n_3431), .B(n_3333), .Z(n_1399));
   NAND4_X1 i_2644 (.A1(a[11]), .A2(a[10]), .A3(b[2]), .A4(b[1]), .ZN(n_3434));
   AOI22_X1 i_2645 (.A1(a[11]), .A2(b[1]), .B1(a[10]), .B2(b[2]), .ZN(n_3435));
   NAND2_X1 i_2646 (.A1(a[9]), .A2(b[3]), .ZN(n_3436));
   OAI21_X1 i_2647 (.A(n_3434), .B1(n_3435), .B2(n_3436), .ZN(n_3437));
   AOI21_X1 i_2648 (.A(n_3437), .B1(a[13]), .B2(b[0]), .ZN(n_3438));
   NAND2_X1 i_2649 (.A1(a[12]), .A2(b[1]), .ZN(n_3441));
   NAND3_X1 i_2650 (.A1(n_3437), .A2(a[13]), .A3(b[0]), .ZN(n_3442));
   AOI21_X1 i_2651 (.A(n_3438), .B1(n_3441), .B2(n_3442), .ZN(n_1349));
   NAND4_X1 i_2652 (.A1(b[12]), .A2(b[11]), .A3(a[2]), .A4(a[1]), .ZN(n_3443));
   AOI22_X1 i_2653 (.A1(b[11]), .A2(a[2]), .B1(b[12]), .B2(a[1]), .ZN(n_3444));
   NAND2_X1 i_2654 (.A1(b[13]), .A2(a[0]), .ZN(n_3445));
   OAI21_X1 i_2655 (.A(n_3443), .B1(n_3444), .B2(n_3445), .ZN(n_1322));
   NAND4_X1 i_2656 (.A1(b[9]), .A2(b[8]), .A3(a[5]), .A4(a[4]), .ZN(n_3448));
   AOI22_X1 i_2657 (.A1(b[8]), .A2(a[5]), .B1(b[9]), .B2(a[4]), .ZN(n_3449));
   NAND2_X1 i_2658 (.A1(b[10]), .A2(a[3]), .ZN(n_3450));
   OAI21_X1 i_2659 (.A(n_3448), .B1(n_3449), .B2(n_3450), .ZN(n_1329));
   NAND4_X1 i_2660 (.A1(a[8]), .A2(a[7]), .A3(b[6]), .A4(b[5]), .ZN(n_3451));
   AOI22_X1 i_2661 (.A1(a[8]), .A2(b[5]), .B1(a[7]), .B2(b[6]), .ZN(n_3452));
   NAND2_X1 i_2662 (.A1(b[7]), .A2(a[6]), .ZN(n_3455));
   OAI21_X1 i_2663 (.A(n_3451), .B1(n_3452), .B2(n_3455), .ZN(n_1336));
   NAND4_X1 i_2664 (.A1(a[11]), .A2(a[10]), .A3(b[3]), .A4(b[2]), .ZN(n_3456));
   AOI22_X1 i_2665 (.A1(a[11]), .A2(b[2]), .B1(a[10]), .B2(b[3]), .ZN(n_3457));
   NAND2_X1 i_2666 (.A1(a[9]), .A2(b[4]), .ZN(n_3458));
   OAI21_X1 i_2667 (.A(n_3456), .B1(n_3457), .B2(n_3458), .ZN(n_1343));
   INV_X1 i_2668 (.A(n_3444), .ZN(n_3459));
   NAND2_X1 i_2669 (.A1(n_3459), .A2(n_3443), .ZN(n_3462));
   XOR2_X1 i_2670 (.A(n_3462), .B(n_3445), .Z(n_1321));
   INV_X1 i_2671 (.A(n_3449), .ZN(n_3463));
   NAND2_X1 i_2672 (.A1(n_3463), .A2(n_3448), .ZN(n_3464));
   XOR2_X1 i_2673 (.A(n_3464), .B(n_3450), .Z(n_1328));
   INV_X1 i_2674 (.A(n_3452), .ZN(n_3465));
   NAND2_X1 i_2675 (.A1(n_3465), .A2(n_3451), .ZN(n_3466));
   XOR2_X1 i_2676 (.A(n_3466), .B(n_3455), .Z(n_1335));
   INV_X1 i_2677 (.A(n_3457), .ZN(n_3468));
   NAND2_X1 i_2678 (.A1(n_3468), .A2(n_3456), .ZN(n_3469));
   XOR2_X1 i_2679 (.A(n_3469), .B(n_3458), .Z(n_1342));
   INV_X1 i_2680 (.A(n_3438), .ZN(n_3470));
   NAND2_X1 i_2681 (.A1(n_3470), .A2(n_3442), .ZN(n_3471));
   XOR2_X1 i_2682 (.A(n_3471), .B(n_3441), .Z(n_1348));
   NAND4_X1 i_2683 (.A1(a[8]), .A2(a[7]), .A3(b[3]), .A4(b[4]), .ZN(n_3472));
   AOI22_X1 i_2684 (.A1(a[8]), .A2(b[3]), .B1(a[7]), .B2(b[4]), .ZN(n_3473));
   NAND2_X1 i_2685 (.A1(a[6]), .A2(b[5]), .ZN(n_3475));
   OAI21_X1 i_2686 (.A(n_3472), .B1(n_3473), .B2(n_3475), .ZN(n_3476));
   NAND4_X1 i_2687 (.A1(a[11]), .A2(a[10]), .A3(b[1]), .A4(b[0]), .ZN(n_3477));
   AOI22_X1 i_2707 (.A1(a[11]), .A2(b[0]), .B1(a[10]), .B2(b[1]), .ZN(n_3478));
   NAND2_X1 i_2708 (.A1(a[9]), .A2(b[2]), .ZN(n_3479));
   OAI21_X1 i_2709 (.A(n_3477), .B1(n_3478), .B2(n_3479), .ZN(n_3482));
   NOR2_X1 i_2710 (.A1(n_3476), .A2(n_3482), .ZN(n_3483));
   NAND2_X1 i_2711 (.A1(a[12]), .A2(b[0]), .ZN(n_3484));
   NAND2_X1 i_2712 (.A1(n_3476), .A2(n_3482), .ZN(n_3485));
   AOI21_X1 i_2713 (.A(n_3483), .B1(n_3484), .B2(n_3485), .ZN(n_1302));
   NAND4_X1 i_2714 (.A1(b[11]), .A2(b[10]), .A3(a[2]), .A4(a[1]), .ZN(n_3486));
   AOI22_X1 i_2715 (.A1(b[10]), .A2(a[2]), .B1(b[11]), .B2(a[1]), .ZN(n_3519));
   NAND2_X1 i_2716 (.A1(b[12]), .A2(a[0]), .ZN(n_3520));
   OAI21_X1 i_2717 (.A(n_3486), .B1(n_3519), .B2(n_3520), .ZN(n_1274));
   NAND4_X1 i_2718 (.A1(b[8]), .A2(b[7]), .A3(a[5]), .A4(a[4]), .ZN(n_3523));
   AOI22_X1 i_2719 (.A1(b[7]), .A2(a[5]), .B1(b[8]), .B2(a[4]), .ZN(n_3524));
   NAND2_X1 i_2720 (.A1(b[9]), .A2(a[3]), .ZN(n_3525));
   OAI21_X1 i_2721 (.A(n_3523), .B1(n_3524), .B2(n_3525), .ZN(n_1281));
   NAND4_X1 i_2722 (.A1(a[8]), .A2(a[7]), .A3(b[4]), .A4(b[5]), .ZN(n_3526));
   AOI22_X1 i_2723 (.A1(a[8]), .A2(b[4]), .B1(a[7]), .B2(b[5]), .ZN(n_3527));
   NAND2_X1 i_2724 (.A1(a[6]), .A2(b[6]), .ZN(n_3530));
   OAI21_X1 i_2725 (.A(n_3526), .B1(n_3527), .B2(n_3530), .ZN(n_1288));
   INV_X1 i_2726 (.A(n_3483), .ZN(n_3531));
   NAND2_X1 i_2727 (.A1(n_3531), .A2(n_3485), .ZN(n_3532));
   XOR2_X1 i_2728 (.A(n_3532), .B(n_3484), .Z(n_1301));
   INV_X1 i_2729 (.A(n_3519), .ZN(n_3533));
   NAND2_X1 i_2730 (.A1(n_3533), .A2(n_3486), .ZN(n_3534));
   XOR2_X1 i_2731 (.A(n_3534), .B(n_3520), .Z(n_1273));
   INV_X1 i_2732 (.A(n_3524), .ZN(n_3537));
   NAND2_X1 i_2733 (.A1(n_3537), .A2(n_3523), .ZN(n_3538));
   XOR2_X1 i_2734 (.A(n_3538), .B(n_3525), .Z(n_1280));
   INV_X1 i_2735 (.A(n_3527), .ZN(n_3539));
   NAND2_X1 i_2736 (.A1(n_3539), .A2(n_3526), .ZN(n_3540));
   XOR2_X1 i_2737 (.A(n_3540), .B(n_3530), .Z(n_1287));
   INV_X1 i_2738 (.A(n_3435), .ZN(n_3541));
   NAND2_X1 i_2739 (.A1(n_3541), .A2(n_3434), .ZN(n_3544));
   XOR2_X1 i_2740 (.A(n_3544), .B(n_3436), .Z(n_1294));
   NAND4_X1 i_2741 (.A1(b[10]), .A2(b[9]), .A3(a[2]), .A4(a[1]), .ZN(n_3545));
   AOI22_X1 i_2742 (.A1(b[9]), .A2(a[2]), .B1(b[10]), .B2(a[1]), .ZN(n_3546));
   NAND2_X1 i_2743 (.A1(b[11]), .A2(a[0]), .ZN(n_3547));
   OAI21_X1 i_2744 (.A(n_3545), .B1(n_3546), .B2(n_3547), .ZN(n_1234));
   NAND4_X1 i_2745 (.A1(b[7]), .A2(a[5]), .A3(b[6]), .A4(a[4]), .ZN(n_3548));
   AOI22_X1 i_2746 (.A1(a[5]), .A2(b[6]), .B1(b[7]), .B2(a[4]), .ZN(n_3551));
   NAND2_X1 i_2747 (.A1(b[8]), .A2(a[3]), .ZN(n_3552));
   OAI21_X1 i_2748 (.A(n_3548), .B1(n_3551), .B2(n_3552), .ZN(n_1241));
   INV_X1 i_2749 (.A(n_3546), .ZN(n_3553));
   NAND2_X1 i_2750 (.A1(n_3553), .A2(n_3545), .ZN(n_3554));
   XOR2_X1 i_2751 (.A(n_3554), .B(n_3547), .Z(n_1233));
   INV_X1 i_2752 (.A(n_3551), .ZN(n_3555));
   NAND2_X1 i_2753 (.A1(n_3555), .A2(n_3548), .ZN(n_3558));
   XOR2_X1 i_2754 (.A(n_3558), .B(n_3552), .Z(n_1240));
   INV_X1 i_2755 (.A(n_3473), .ZN(n_3559));
   NAND2_X1 i_2756 (.A1(n_3559), .A2(n_3472), .ZN(n_3560));
   XOR2_X1 i_2757 (.A(n_3560), .B(n_3475), .Z(n_1247));
   INV_X1 i_2758 (.A(n_3478), .ZN(n_3561));
   NAND2_X1 i_2759 (.A1(n_3561), .A2(n_3477), .ZN(n_3562));
   XOR2_X1 i_2760 (.A(n_3562), .B(n_3479), .Z(n_1254));
   NAND4_X1 i_2761 (.A1(a[8]), .A2(a[7]), .A3(b[2]), .A4(b[1]), .ZN(n_3565));
   AOI22_X1 i_2762 (.A1(a[8]), .A2(b[1]), .B1(a[7]), .B2(b[2]), .ZN(n_3566));
   NAND2_X1 i_2763 (.A1(b[3]), .A2(a[6]), .ZN(n_3567));
   OAI21_X1 i_2764 (.A(n_3565), .B1(n_3566), .B2(n_3567), .ZN(n_3568));
   AOI21_X1 i_2765 (.A(n_3568), .B1(a[10]), .B2(b[0]), .ZN(n_3569));
   NAND2_X1 i_2766 (.A1(a[9]), .A2(b[1]), .ZN(n_3572));
   NAND3_X1 i_2767 (.A1(n_3568), .A2(a[10]), .A3(b[0]), .ZN(n_3573));
   AOI21_X1 i_2768 (.A(n_3569), .B1(n_3572), .B2(n_3573), .ZN(n_1215));
   NAND4_X1 i_2769 (.A1(b[9]), .A2(b[8]), .A3(a[2]), .A4(a[1]), .ZN(n_3574));
   AOI22_X1 i_2770 (.A1(b[8]), .A2(a[2]), .B1(b[9]), .B2(a[1]), .ZN(n_3575));
   NAND2_X1 i_2771 (.A1(b[10]), .A2(a[0]), .ZN(n_3576));
   OAI21_X1 i_2772 (.A(n_3574), .B1(n_3575), .B2(n_3576), .ZN(n_1195));
   NAND4_X1 i_2773 (.A1(a[5]), .A2(b[6]), .A3(b[5]), .A4(a[4]), .ZN(n_3579));
   AOI22_X1 i_2774 (.A1(a[5]), .A2(b[5]), .B1(b[6]), .B2(a[4]), .ZN(n_3580));
   NAND2_X1 i_2775 (.A1(b[7]), .A2(a[3]), .ZN(n_3581));
   OAI21_X1 i_2776 (.A(n_3579), .B1(n_3580), .B2(n_3581), .ZN(n_1202));
   NAND4_X1 i_2796 (.A1(a[8]), .A2(a[7]), .A3(b[3]), .A4(b[2]), .ZN(n_3582));
   AOI22_X1 i_2797 (.A1(a[8]), .A2(b[2]), .B1(a[7]), .B2(b[3]), .ZN(n_3613));
   NAND2_X1 i_2798 (.A1(a[6]), .A2(b[4]), .ZN(n_3614));
   OAI21_X1 i_2799 (.A(n_3582), .B1(n_3613), .B2(n_3614), .ZN(n_1209));
   INV_X1 i_2800 (.A(n_3575), .ZN(n_3617));
   NAND2_X1 i_2801 (.A1(n_3617), .A2(n_3574), .ZN(n_3618));
   XOR2_X1 i_2802 (.A(n_3618), .B(n_3576), .Z(n_1194));
   INV_X1 i_2803 (.A(n_3580), .ZN(n_3619));
   NAND2_X1 i_2804 (.A1(n_3619), .A2(n_3579), .ZN(n_3620));
   XOR2_X1 i_2805 (.A(n_3620), .B(n_3581), .Z(n_1201));
   INV_X1 i_2806 (.A(n_3613), .ZN(n_3621));
   NAND2_X1 i_2807 (.A1(n_3621), .A2(n_3582), .ZN(n_3624));
   XOR2_X1 i_2808 (.A(n_3624), .B(n_3614), .Z(n_1208));
   INV_X1 i_2809 (.A(n_3569), .ZN(n_3625));
   NAND2_X1 i_2810 (.A1(n_3625), .A2(n_3573), .ZN(n_3626));
   XOR2_X1 i_2811 (.A(n_3626), .B(n_3572), .Z(n_1214));
   NAND4_X1 i_2812 (.A1(b[3]), .A2(a[5]), .A3(b[4]), .A4(a[4]), .ZN(n_3627));
   AOI22_X1 i_2813 (.A1(b[3]), .A2(a[5]), .B1(b[4]), .B2(a[4]), .ZN(n_3628));
   NAND2_X1 i_2814 (.A1(b[5]), .A2(a[3]), .ZN(n_3631));
   OAI21_X1 i_2815 (.A(n_3627), .B1(n_3628), .B2(n_3631), .ZN(n_3632));
   NAND4_X1 i_2816 (.A1(a[8]), .A2(a[7]), .A3(b[1]), .A4(b[0]), .ZN(n_3633));
   AOI22_X1 i_2817 (.A1(a[8]), .A2(b[0]), .B1(a[7]), .B2(b[1]), .ZN(n_3634));
   NAND2_X1 i_2818 (.A1(b[2]), .A2(a[6]), .ZN(n_3635));
   OAI21_X1 i_2819 (.A(n_3633), .B1(n_3634), .B2(n_3635), .ZN(n_3638));
   NOR2_X1 i_2820 (.A1(n_3632), .A2(n_3638), .ZN(n_3639));
   NAND2_X1 i_2821 (.A1(a[9]), .A2(b[0]), .ZN(n_3640));
   NAND2_X1 i_2822 (.A1(n_3632), .A2(n_3638), .ZN(n_3641));
   AOI21_X1 i_2823 (.A(n_3639), .B1(n_3640), .B2(n_3641), .ZN(n_1179));
   NAND4_X1 i_2824 (.A1(b[8]), .A2(b[7]), .A3(a[2]), .A4(a[1]), .ZN(n_3642));
   AOI22_X1 i_2825 (.A1(b[7]), .A2(a[2]), .B1(b[8]), .B2(a[1]), .ZN(n_3645));
   NAND2_X1 i_2826 (.A1(b[9]), .A2(a[0]), .ZN(n_3646));
   OAI21_X1 i_2827 (.A(n_3642), .B1(n_3645), .B2(n_3646), .ZN(n_1158));
   NAND4_X1 i_2828 (.A1(a[5]), .A2(b[4]), .A3(b[5]), .A4(a[4]), .ZN(n_3647));
   AOI22_X1 i_2829 (.A1(a[5]), .A2(b[4]), .B1(b[5]), .B2(a[4]), .ZN(n_3648));
   NAND2_X1 i_2830 (.A1(b[6]), .A2(a[3]), .ZN(n_3649));
   OAI21_X1 i_2831 (.A(n_3647), .B1(n_3648), .B2(n_3649), .ZN(n_1165));
   INV_X1 i_2832 (.A(n_3639), .ZN(n_3652));
   NAND2_X1 i_2833 (.A1(n_3652), .A2(n_3641), .ZN(n_3653));
   XOR2_X1 i_2834 (.A(n_3653), .B(n_3640), .Z(n_1178));
   INV_X1 i_2835 (.A(n_3645), .ZN(n_3654));
   NAND2_X1 i_2836 (.A1(n_3654), .A2(n_3642), .ZN(n_3655));
   XOR2_X1 i_2837 (.A(n_3655), .B(n_3646), .Z(n_1157));
   INV_X1 i_2838 (.A(n_3648), .ZN(n_3656));
   NAND2_X1 i_2839 (.A1(n_3656), .A2(n_3647), .ZN(n_3659));
   XOR2_X1 i_2840 (.A(n_3659), .B(n_3649), .Z(n_1164));
   INV_X1 i_2841 (.A(n_3566), .ZN(n_3660));
   NAND2_X1 i_2842 (.A1(n_3660), .A2(n_3565), .ZN(n_3661));
   XOR2_X1 i_2843 (.A(n_3661), .B(n_3567), .Z(n_1171));
   NAND4_X1 i_2844 (.A1(b[7]), .A2(b[6]), .A3(a[2]), .A4(a[1]), .ZN(n_3662));
   AOI22_X1 i_2845 (.A1(b[6]), .A2(a[2]), .B1(b[7]), .B2(a[1]), .ZN(n_3663));
   NAND2_X1 i_2846 (.A1(b[8]), .A2(a[0]), .ZN(n_3665));
   OAI21_X1 i_2847 (.A(n_3662), .B1(n_3663), .B2(n_3665), .ZN(n_1129));
   INV_X1 i_2848 (.A(n_3663), .ZN(n_3666));
   NAND2_X1 i_2849 (.A1(n_3666), .A2(n_3662), .ZN(n_3667));
   XOR2_X1 i_2850 (.A(n_3667), .B(n_3665), .Z(n_1128));
   INV_X1 i_2851 (.A(n_3628), .ZN(n_3668));
   NAND2_X1 i_2852 (.A1(n_3668), .A2(n_3627), .ZN(n_3699));
   XOR2_X1 i_2853 (.A(n_3699), .B(n_3631), .Z(n_1135));
   INV_X1 i_2854 (.A(n_3634), .ZN(n_3700));
   NAND2_X1 i_2855 (.A1(n_3700), .A2(n_3633), .ZN(n_3703));
   XOR2_X1 i_2856 (.A(n_3703), .B(n_3635), .Z(n_1142));
   NAND2_X1 i_2857 (.A1(a[4]), .A2(b[1]), .ZN(n_3704));
   NAND2_X1 i_2858 (.A1(b[2]), .A2(a[5]), .ZN(n_3705));
   NOR2_X1 i_2859 (.A1(n_3704), .A2(n_3705), .ZN(n_3706));
   INV_X1 i_2860 (.A(n_3706), .ZN(n_3707));
   AOI22_X1 i_2861 (.A1(a[5]), .A2(b[1]), .B1(b[2]), .B2(a[4]), .ZN(n_3710));
   NAND2_X1 i_2862 (.A1(b[3]), .A2(a[3]), .ZN(n_3711));
   OAI21_X1 i_2863 (.A(n_3707), .B1(n_3710), .B2(n_3711), .ZN(n_3712));
   AOI21_X1 i_2864 (.A(n_3712), .B1(a[7]), .B2(b[0]), .ZN(n_3713));
   NAND2_X1 i_2865 (.A1(a[6]), .A2(b[1]), .ZN(n_3714));
   NAND3_X1 i_2866 (.A1(n_3712), .A2(a[7]), .A3(b[0]), .ZN(n_3717));
   AOI21_X1 i_2885 (.A(n_3713), .B1(n_3714), .B2(n_3717), .ZN(n_1114));
   NAND4_X1 i_2886 (.A1(b[6]), .A2(a[2]), .A3(b[5]), .A4(a[1]), .ZN(n_3718));
   AOI22_X1 i_2887 (.A1(a[2]), .A2(b[5]), .B1(b[6]), .B2(a[1]), .ZN(n_3719));
   NAND2_X1 i_2888 (.A1(b[7]), .A2(a[0]), .ZN(n_3720));
   OAI21_X1 i_2889 (.A(n_3718), .B1(n_3719), .B2(n_3720), .ZN(n_1101));
   INV_X1 i_2890 (.A(n_3705), .ZN(n_3721));
   NAND3_X1 i_2891 (.A1(n_3721), .A2(b[3]), .A3(a[4]), .ZN(n_3724));
   AOI21_X1 i_2892 (.A(n_3721), .B1(b[3]), .B2(a[4]), .ZN(n_3725));
   NAND2_X1 i_2893 (.A1(b[4]), .A2(a[3]), .ZN(n_3726));
   OAI21_X1 i_2894 (.A(n_3724), .B1(n_3725), .B2(n_3726), .ZN(n_1108));
   INV_X1 i_2895 (.A(n_3719), .ZN(n_3727));
   NAND2_X1 i_2896 (.A1(n_3727), .A2(n_3718), .ZN(n_3728));
   XOR2_X1 i_2897 (.A(n_3728), .B(n_3720), .Z(n_1100));
   INV_X1 i_2898 (.A(n_3725), .ZN(n_3731));
   NAND2_X1 i_2899 (.A1(n_3724), .A2(n_3731), .ZN(n_3732));
   XOR2_X1 i_2900 (.A(n_3732), .B(n_3726), .Z(n_1107));
   INV_X1 i_2901 (.A(n_3713), .ZN(n_3733));
   NAND2_X1 i_2902 (.A1(n_3733), .A2(n_3717), .ZN(n_3734));
   XOR2_X1 i_2903 (.A(n_3734), .B(n_3714), .Z(n_1113));
   INV_X1 i_2904 (.A(a[1]), .ZN(n_3735));
   OR3_X1 i_2905 (.A1(n_508), .A2(n_1561), .A3(n_3735), .ZN(n_3737));
   INV_X1 i_2906 (.A(n_3737), .ZN(n_3738));
   NOR2_X1 i_2907 (.A1(n_1232), .A2(n_513), .ZN(n_3739));
   OAI21_X1 i_2908 (.A(n_508), .B1(n_1561), .B2(n_3735), .ZN(n_3740));
   AOI21_X1 i_2909 (.A(n_3738), .B1(n_3739), .B2(n_3740), .ZN(n_3741));
   INV_X1 i_2910 (.A(a[5]), .ZN(n_3742));
   OR3_X1 i_2911 (.A1(n_3704), .A2(n_3742), .A3(n_514), .ZN(n_3744));
   INV_X1 i_2912 (.A(n_3744), .ZN(n_3745));
   AND2_X1 i_2913 (.A1(b[2]), .A2(a[3]), .ZN(n_3746));
   OAI21_X1 i_2914 (.A(n_3704), .B1(n_3742), .B2(n_514), .ZN(n_3747));
   AOI21_X1 i_2915 (.A(n_3745), .B1(n_3746), .B2(n_3747), .ZN(n_3748));
   NAND2_X1 i_2916 (.A1(n_3741), .A2(n_3748), .ZN(n_3751));
   INV_X1 i_2917 (.A(n_3751), .ZN(n_3752));
   NAND2_X1 i_2918 (.A1(a[6]), .A2(b[0]), .ZN(n_3753));
   OR2_X1 i_2919 (.A1(n_3741), .A2(n_3748), .ZN(n_3754));
   AOI21_X1 i_2920 (.A(n_3752), .B1(n_3753), .B2(n_3754), .ZN(n_1089));
   NAND4_X1 i_2921 (.A1(b[4]), .A2(a[2]), .A3(b[5]), .A4(a[1]), .ZN(n_3755));
   AOI22_X1 i_2922 (.A1(b[4]), .A2(a[2]), .B1(b[5]), .B2(a[1]), .ZN(n_3784));
   NAND2_X1 i_2923 (.A1(b[6]), .A2(a[0]), .ZN(n_3785));
   OAI21_X1 i_2924 (.A(n_3755), .B1(n_3784), .B2(n_3785), .ZN(n_1075));
   NAND2_X1 i_2925 (.A1(n_3754), .A2(n_3751), .ZN(n_3788));
   XOR2_X1 i_2926 (.A(n_3788), .B(n_3753), .Z(n_1088));
   INV_X1 i_2927 (.A(n_3784), .ZN(n_3789));
   NAND2_X1 i_2928 (.A1(n_3789), .A2(n_3755), .ZN(n_3790));
   XOR2_X1 i_2929 (.A(n_3790), .B(n_3785), .Z(n_1074));
   NOR2_X1 i_2930 (.A1(n_3706), .A2(n_3710), .ZN(n_3791));
   XNOR2_X1 i_2931 (.A(n_3791), .B(n_3711), .ZN(n_1081));
   NAND2_X1 i_2932 (.A1(n_3737), .A2(n_3740), .ZN(n_3792));
   XNOR2_X1 i_2933 (.A(n_3792), .B(n_3739), .ZN(n_1056));
   NAND2_X1 i_2934 (.A1(n_3744), .A2(n_3747), .ZN(n_3795));
   XNOR2_X1 i_2935 (.A(n_3795), .B(n_3746), .ZN(n_1063));
   INV_X1 i_2936 (.A(n_509), .ZN(n_3796));
   AOI21_X1 i_2937 (.A(n_510), .B1(n_3796), .B2(n_512), .ZN(n_1040));
   AOI21_X1 i_2938 (.A(n_528), .B1(n_516), .B2(n_3704), .ZN(n_1046));
   AOI22_X1 i_2939 (.A1(a[3]), .A2(b[1]), .B1(a[4]), .B2(b[0]), .ZN(n_3797));
   NAND3_X1 i_2940 (.A1(a[4]), .A2(a[3]), .A3(b[0]), .ZN(n_3798));
   OAI22_X1 i_2941 (.A1(n_1046), .A2(n_3797), .B1(n_516), .B2(n_3798), .ZN(
      n_1045));
   OAI21_X1 i_2942 (.A(n_523), .B1(n_524), .B2(n_527), .ZN(n_1030));
   INV_X1 i_2943 (.A(n_521), .ZN(n_3799));
   AOI22_X1 i_2944 (.A1(b[1]), .A2(a[0]), .B1(b[0]), .B2(a[1]), .ZN(n_3802));
   NOR2_X1 i_2945 (.A1(n_3799), .A2(n_3802), .ZN(p_0[1]));
   INV_X1 i_2946 (.A(n_520), .ZN(n_3803));
   NAND2_X1 i_2947 (.A1(n_3803), .A2(n_522), .ZN(n_3804));
   XOR2_X1 i_2948 (.A(n_3804), .B(n_521), .Z(p_0[2]));
   INV_X1 i_2949 (.A(n_504), .ZN(n_3805));
   OAI21_X1 i_2950 (.A(n_3805), .B1(n_502), .B2(n_505), .ZN(n_3806));
   INV_X1 i_2951 (.A(n_503), .ZN(n_3809));
   NAND2_X1 i_2952 (.A1(n_3809), .A2(n_338), .ZN(n_3810));
   NOR2_X1 i_2953 (.A1(n_3809), .A2(n_338), .ZN(n_3811));
   INV_X1 i_2954 (.A(n_3811), .ZN(n_3812));
   NAND2_X1 i_2955 (.A1(n_3810), .A2(n_3812), .ZN(n_3813));
   XNOR2_X1 i_2973 (.A(n_3806), .B(n_3813), .ZN(p_0[62]));
   INV_X1 i_2974 (.A(n_3806), .ZN(n_3816));
   OAI21_X1 i_2975 (.A(n_3810), .B1(n_3816), .B2(n_3811), .ZN(p_0[63]));
endmodule

module multOperator(clk, rst, a, b, c);
   input clk;
   input rst;
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   DFFR_X1 \c_reg[63]  (.D(n_64), .RN(n_0), .CK(clk), .Q(c[63]), .QN());
   INV_X1 i_0_0 (.A(rst), .ZN(n_0));
   DFFR_X1 \c_reg[62]  (.D(n_63), .RN(n_0), .CK(clk), .Q(c[62]), .QN());
   DFFR_X1 \c_reg[61]  (.D(n_62), .RN(n_0), .CK(clk), .Q(c[61]), .QN());
   DFFR_X1 \c_reg[60]  (.D(n_61), .RN(n_0), .CK(clk), .Q(c[60]), .QN());
   DFFR_X1 \c_reg[59]  (.D(n_60), .RN(n_0), .CK(clk), .Q(c[59]), .QN());
   DFFR_X1 \c_reg[58]  (.D(n_59), .RN(n_0), .CK(clk), .Q(c[58]), .QN());
   DFFR_X1 \c_reg[57]  (.D(n_58), .RN(n_0), .CK(clk), .Q(c[57]), .QN());
   DFFR_X1 \c_reg[56]  (.D(n_57), .RN(n_0), .CK(clk), .Q(c[56]), .QN());
   DFFR_X1 \c_reg[55]  (.D(n_56), .RN(n_0), .CK(clk), .Q(c[55]), .QN());
   DFFR_X1 \c_reg[54]  (.D(n_55), .RN(n_0), .CK(clk), .Q(c[54]), .QN());
   DFFR_X1 \c_reg[53]  (.D(n_54), .RN(n_0), .CK(clk), .Q(c[53]), .QN());
   DFFR_X1 \c_reg[52]  (.D(n_53), .RN(n_0), .CK(clk), .Q(c[52]), .QN());
   DFFR_X1 \c_reg[51]  (.D(n_52), .RN(n_0), .CK(clk), .Q(c[51]), .QN());
   DFFR_X1 \c_reg[50]  (.D(n_51), .RN(n_0), .CK(clk), .Q(c[50]), .QN());
   DFFR_X1 \c_reg[49]  (.D(n_50), .RN(n_0), .CK(clk), .Q(c[49]), .QN());
   DFFR_X1 \c_reg[48]  (.D(n_49), .RN(n_0), .CK(clk), .Q(c[48]), .QN());
   DFFR_X1 \c_reg[47]  (.D(n_48), .RN(n_0), .CK(clk), .Q(c[47]), .QN());
   DFFR_X1 \c_reg[46]  (.D(n_47), .RN(n_0), .CK(clk), .Q(c[46]), .QN());
   DFFR_X1 \c_reg[45]  (.D(n_46), .RN(n_0), .CK(clk), .Q(c[45]), .QN());
   DFFR_X1 \c_reg[44]  (.D(n_45), .RN(n_0), .CK(clk), .Q(c[44]), .QN());
   DFFR_X1 \c_reg[43]  (.D(n_44), .RN(n_0), .CK(clk), .Q(c[43]), .QN());
   DFFR_X1 \c_reg[42]  (.D(n_43), .RN(n_0), .CK(clk), .Q(c[42]), .QN());
   DFFR_X1 \c_reg[41]  (.D(n_42), .RN(n_0), .CK(clk), .Q(c[41]), .QN());
   DFFR_X1 \c_reg[40]  (.D(n_41), .RN(n_0), .CK(clk), .Q(c[40]), .QN());
   DFFR_X1 \c_reg[39]  (.D(n_40), .RN(n_0), .CK(clk), .Q(c[39]), .QN());
   DFFR_X1 \c_reg[38]  (.D(n_39), .RN(n_0), .CK(clk), .Q(c[38]), .QN());
   DFFR_X1 \c_reg[37]  (.D(n_38), .RN(n_0), .CK(clk), .Q(c[37]), .QN());
   DFFR_X1 \c_reg[36]  (.D(n_37), .RN(n_0), .CK(clk), .Q(c[36]), .QN());
   DFFR_X1 \c_reg[35]  (.D(n_36), .RN(n_0), .CK(clk), .Q(c[35]), .QN());
   DFFR_X1 \c_reg[34]  (.D(n_35), .RN(n_0), .CK(clk), .Q(c[34]), .QN());
   DFFR_X1 \c_reg[33]  (.D(n_34), .RN(n_0), .CK(clk), .Q(c[33]), .QN());
   DFFR_X1 \c_reg[32]  (.D(n_33), .RN(n_0), .CK(clk), .Q(c[32]), .QN());
   DFFR_X1 \c_reg[31]  (.D(n_32), .RN(n_0), .CK(clk), .Q(c[31]), .QN());
   DFFR_X1 \c_reg[30]  (.D(n_31), .RN(n_0), .CK(clk), .Q(c[30]), .QN());
   DFFR_X1 \c_reg[29]  (.D(n_30), .RN(n_0), .CK(clk), .Q(c[29]), .QN());
   DFFR_X1 \c_reg[28]  (.D(n_29), .RN(n_0), .CK(clk), .Q(c[28]), .QN());
   DFFR_X1 \c_reg[27]  (.D(n_28), .RN(n_0), .CK(clk), .Q(c[27]), .QN());
   DFFR_X1 \c_reg[26]  (.D(n_27), .RN(n_0), .CK(clk), .Q(c[26]), .QN());
   DFFR_X1 \c_reg[25]  (.D(n_26), .RN(n_0), .CK(clk), .Q(c[25]), .QN());
   DFFR_X1 \c_reg[24]  (.D(n_25), .RN(n_0), .CK(clk), .Q(c[24]), .QN());
   DFFR_X1 \c_reg[23]  (.D(n_24), .RN(n_0), .CK(clk), .Q(c[23]), .QN());
   DFFR_X1 \c_reg[22]  (.D(n_23), .RN(n_0), .CK(clk), .Q(c[22]), .QN());
   DFFR_X1 \c_reg[21]  (.D(n_22), .RN(n_0), .CK(clk), .Q(c[21]), .QN());
   DFFR_X1 \c_reg[20]  (.D(n_21), .RN(n_0), .CK(clk), .Q(c[20]), .QN());
   DFFR_X1 \c_reg[19]  (.D(n_20), .RN(n_0), .CK(clk), .Q(c[19]), .QN());
   DFFR_X1 \c_reg[18]  (.D(n_19), .RN(n_0), .CK(clk), .Q(c[18]), .QN());
   DFFR_X1 \c_reg[17]  (.D(n_18), .RN(n_0), .CK(clk), .Q(c[17]), .QN());
   DFFR_X1 \c_reg[16]  (.D(n_17), .RN(n_0), .CK(clk), .Q(c[16]), .QN());
   DFFR_X1 \c_reg[15]  (.D(n_16), .RN(n_0), .CK(clk), .Q(c[15]), .QN());
   DFFR_X1 \c_reg[14]  (.D(n_15), .RN(n_0), .CK(clk), .Q(c[14]), .QN());
   DFFR_X1 \c_reg[13]  (.D(n_14), .RN(n_0), .CK(clk), .Q(c[13]), .QN());
   DFFR_X1 \c_reg[12]  (.D(n_13), .RN(n_0), .CK(clk), .Q(c[12]), .QN());
   DFFR_X1 \c_reg[11]  (.D(n_12), .RN(n_0), .CK(clk), .Q(c[11]), .QN());
   DFFR_X1 \c_reg[10]  (.D(n_11), .RN(n_0), .CK(clk), .Q(c[10]), .QN());
   DFFR_X1 \c_reg[9]  (.D(n_10), .RN(n_0), .CK(clk), .Q(c[9]), .QN());
   DFFR_X1 \c_reg[8]  (.D(n_9), .RN(n_0), .CK(clk), .Q(c[8]), .QN());
   DFFR_X1 \c_reg[7]  (.D(n_8), .RN(n_0), .CK(clk), .Q(c[7]), .QN());
   DFFR_X1 \c_reg[6]  (.D(n_7), .RN(n_0), .CK(clk), .Q(c[6]), .QN());
   DFFR_X1 \c_reg[5]  (.D(n_6), .RN(n_0), .CK(clk), .Q(c[5]), .QN());
   DFFR_X1 \c_reg[4]  (.D(n_5), .RN(n_0), .CK(clk), .Q(c[4]), .QN());
   DFFR_X1 \c_reg[3]  (.D(n_4), .RN(n_0), .CK(clk), .Q(c[3]), .QN());
   DFFR_X1 \c_reg[2]  (.D(n_3), .RN(n_0), .CK(clk), .Q(c[2]), .QN());
   DFFR_X1 \c_reg[1]  (.D(n_2), .RN(n_0), .CK(clk), .Q(c[1]), .QN());
   DFFR_X1 \c_reg[0]  (.D(n_1), .RN(n_0), .CK(clk), .Q(c[0]), .QN());
   datapath i_1 (.b(b), .a(a), .p_0({n_64, n_63, n_62, n_61, n_60, n_59, n_58, 
      n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, 
      n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, 
      n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, 
      n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, 
      n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1}));
endmodule

module buffer__parameterized0(clk, rst, D, Q);
   input clk;
   input rst;
   input [63:0]D;
   output [63:0]Q;

   wire n_0_0;

   DFF_X1 \Q_reg[63]  (.D(n_63), .CK(clk), .Q(Q[63]), .QN());
   DFF_X1 \Q_reg[62]  (.D(n_62), .CK(clk), .Q(Q[62]), .QN());
   DFF_X1 \Q_reg[61]  (.D(n_61), .CK(clk), .Q(Q[61]), .QN());
   DFF_X1 \Q_reg[60]  (.D(n_60), .CK(clk), .Q(Q[60]), .QN());
   DFF_X1 \Q_reg[59]  (.D(n_59), .CK(clk), .Q(Q[59]), .QN());
   DFF_X1 \Q_reg[58]  (.D(n_58), .CK(clk), .Q(Q[58]), .QN());
   DFF_X1 \Q_reg[57]  (.D(n_57), .CK(clk), .Q(Q[57]), .QN());
   DFF_X1 \Q_reg[56]  (.D(n_56), .CK(clk), .Q(Q[56]), .QN());
   DFF_X1 \Q_reg[55]  (.D(n_55), .CK(clk), .Q(Q[55]), .QN());
   DFF_X1 \Q_reg[54]  (.D(n_54), .CK(clk), .Q(Q[54]), .QN());
   DFF_X1 \Q_reg[53]  (.D(n_53), .CK(clk), .Q(Q[53]), .QN());
   DFF_X1 \Q_reg[52]  (.D(n_52), .CK(clk), .Q(Q[52]), .QN());
   DFF_X1 \Q_reg[51]  (.D(n_51), .CK(clk), .Q(Q[51]), .QN());
   DFF_X1 \Q_reg[50]  (.D(n_50), .CK(clk), .Q(Q[50]), .QN());
   DFF_X1 \Q_reg[49]  (.D(n_49), .CK(clk), .Q(Q[49]), .QN());
   DFF_X1 \Q_reg[48]  (.D(n_48), .CK(clk), .Q(Q[48]), .QN());
   DFF_X1 \Q_reg[47]  (.D(n_47), .CK(clk), .Q(Q[47]), .QN());
   DFF_X1 \Q_reg[46]  (.D(n_46), .CK(clk), .Q(Q[46]), .QN());
   DFF_X1 \Q_reg[45]  (.D(n_45), .CK(clk), .Q(Q[45]), .QN());
   DFF_X1 \Q_reg[44]  (.D(n_44), .CK(clk), .Q(Q[44]), .QN());
   DFF_X1 \Q_reg[43]  (.D(n_43), .CK(clk), .Q(Q[43]), .QN());
   DFF_X1 \Q_reg[42]  (.D(n_42), .CK(clk), .Q(Q[42]), .QN());
   DFF_X1 \Q_reg[41]  (.D(n_41), .CK(clk), .Q(Q[41]), .QN());
   DFF_X1 \Q_reg[40]  (.D(n_40), .CK(clk), .Q(Q[40]), .QN());
   DFF_X1 \Q_reg[39]  (.D(n_39), .CK(clk), .Q(Q[39]), .QN());
   DFF_X1 \Q_reg[38]  (.D(n_38), .CK(clk), .Q(Q[38]), .QN());
   DFF_X1 \Q_reg[37]  (.D(n_37), .CK(clk), .Q(Q[37]), .QN());
   DFF_X1 \Q_reg[36]  (.D(n_36), .CK(clk), .Q(Q[36]), .QN());
   DFF_X1 \Q_reg[35]  (.D(n_35), .CK(clk), .Q(Q[35]), .QN());
   DFF_X1 \Q_reg[34]  (.D(n_34), .CK(clk), .Q(Q[34]), .QN());
   DFF_X1 \Q_reg[33]  (.D(n_33), .CK(clk), .Q(Q[33]), .QN());
   DFF_X1 \Q_reg[32]  (.D(n_32), .CK(clk), .Q(Q[32]), .QN());
   DFF_X1 \Q_reg[31]  (.D(n_31), .CK(clk), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_30), .CK(clk), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_29), .CK(clk), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_28), .CK(clk), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_27), .CK(clk), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_26), .CK(clk), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_25), .CK(clk), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_24), .CK(clk), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_23), .CK(clk), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_22), .CK(clk), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_21), .CK(clk), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_20), .CK(clk), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_19), .CK(clk), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_18), .CK(clk), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_17), .CK(clk), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_16), .CK(clk), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(clk), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(clk), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(clk), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(clk), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(clk), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(clk), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(clk), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(clk), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(clk), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(clk), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(clk), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(clk), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(clk), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(clk), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(clk), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(clk), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_1 (.A1(n_0_0), .A2(D[0]), .ZN(n_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[1]), .ZN(n_1));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[2]), .ZN(n_2));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[3]), .ZN(n_3));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[4]), .ZN(n_4));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[5]), .ZN(n_5));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[6]), .ZN(n_6));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[7]), .ZN(n_7));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[8]), .ZN(n_8));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[9]), .ZN(n_9));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[10]), .ZN(n_10));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[11]), .ZN(n_11));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[12]), .ZN(n_12));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[13]), .ZN(n_13));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[14]), .ZN(n_14));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[15]), .ZN(n_15));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[16]), .ZN(n_16));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[17]), .ZN(n_17));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[18]), .ZN(n_18));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[19]), .ZN(n_19));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[20]), .ZN(n_20));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[21]), .ZN(n_21));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[22]), .ZN(n_22));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[23]), .ZN(n_23));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[24]), .ZN(n_24));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[25]), .ZN(n_25));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[26]), .ZN(n_26));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[27]), .ZN(n_27));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[28]), .ZN(n_28));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[29]), .ZN(n_29));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[30]), .ZN(n_30));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[31]), .ZN(n_31));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(D[32]), .ZN(n_32));
   AND2_X1 i_0_34 (.A1(n_0_0), .A2(D[33]), .ZN(n_33));
   AND2_X1 i_0_35 (.A1(n_0_0), .A2(D[34]), .ZN(n_34));
   AND2_X1 i_0_36 (.A1(n_0_0), .A2(D[35]), .ZN(n_35));
   AND2_X1 i_0_37 (.A1(n_0_0), .A2(D[36]), .ZN(n_36));
   AND2_X1 i_0_38 (.A1(n_0_0), .A2(D[37]), .ZN(n_37));
   AND2_X1 i_0_39 (.A1(n_0_0), .A2(D[38]), .ZN(n_38));
   AND2_X1 i_0_40 (.A1(n_0_0), .A2(D[39]), .ZN(n_39));
   AND2_X1 i_0_41 (.A1(n_0_0), .A2(D[40]), .ZN(n_40));
   AND2_X1 i_0_42 (.A1(n_0_0), .A2(D[41]), .ZN(n_41));
   AND2_X1 i_0_43 (.A1(n_0_0), .A2(D[42]), .ZN(n_42));
   AND2_X1 i_0_44 (.A1(n_0_0), .A2(D[43]), .ZN(n_43));
   AND2_X1 i_0_45 (.A1(n_0_0), .A2(D[44]), .ZN(n_44));
   AND2_X1 i_0_46 (.A1(n_0_0), .A2(D[45]), .ZN(n_45));
   AND2_X1 i_0_47 (.A1(n_0_0), .A2(D[46]), .ZN(n_46));
   AND2_X1 i_0_48 (.A1(n_0_0), .A2(D[47]), .ZN(n_47));
   AND2_X1 i_0_49 (.A1(n_0_0), .A2(D[48]), .ZN(n_48));
   AND2_X1 i_0_50 (.A1(n_0_0), .A2(D[49]), .ZN(n_49));
   AND2_X1 i_0_51 (.A1(n_0_0), .A2(D[50]), .ZN(n_50));
   AND2_X1 i_0_52 (.A1(n_0_0), .A2(D[51]), .ZN(n_51));
   AND2_X1 i_0_53 (.A1(n_0_0), .A2(D[52]), .ZN(n_52));
   AND2_X1 i_0_54 (.A1(n_0_0), .A2(D[53]), .ZN(n_53));
   AND2_X1 i_0_55 (.A1(n_0_0), .A2(D[54]), .ZN(n_54));
   AND2_X1 i_0_56 (.A1(n_0_0), .A2(D[55]), .ZN(n_55));
   AND2_X1 i_0_57 (.A1(n_0_0), .A2(D[56]), .ZN(n_56));
   AND2_X1 i_0_58 (.A1(n_0_0), .A2(D[57]), .ZN(n_57));
   AND2_X1 i_0_59 (.A1(n_0_0), .A2(D[58]), .ZN(n_58));
   AND2_X1 i_0_60 (.A1(n_0_0), .A2(D[59]), .ZN(n_59));
   AND2_X1 i_0_61 (.A1(n_0_0), .A2(D[60]), .ZN(n_60));
   AND2_X1 i_0_62 (.A1(n_0_0), .A2(D[61]), .ZN(n_61));
   AND2_X1 i_0_63 (.A1(n_0_0), .A2(D[62]), .ZN(n_62));
   AND2_X1 i_0_64 (.A1(n_0_0), .A2(D[63]), .ZN(n_63));
endmodule

module simpleMultiplier(clk, rst, a, b, c);
   input clk;
   input rst;
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   wire [31:0]a_out;
   wire [31:0]b_out;
   wire [63:0]c_out;

   buffer__0_65 inRegA (.clk(clk), .rst(rst), .D(a), .Q(a_out));
   buffer inRegB (.clk(clk), .rst(rst), .D(b), .Q(b_out));
   multOperator M64 (.clk(clk), .rst(rst), .a(a_out), .b(b_out), .c(c_out));
   buffer__parameterized0 outReg (.clk(clk), .rst(rst), .D(c_out), .Q(c));
endmodule
