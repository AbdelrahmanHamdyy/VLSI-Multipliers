/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Dec 27 13:48:12 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3445685297 */

module datapath(a, p_0);
   input [31:0]a;
   output [31:0]p_0;

   AOI21_X1 i_0 (.A(n_62), .B1(a[1]), .B2(a[0]), .ZN(p_0[1]));
   AOI21_X1 i_1 (.A(n_60), .B1(a[2]), .B2(n_61), .ZN(p_0[2]));
   AOI21_X1 i_2 (.A(n_58), .B1(a[3]), .B2(n_59), .ZN(p_0[3]));
   AOI21_X1 i_3 (.A(n_5), .B1(a[4]), .B2(n_57), .ZN(p_0[4]));
   AOI21_X1 i_4 (.A(n_3), .B1(a[5]), .B2(n_4), .ZN(p_0[5]));
   AOI21_X1 i_5 (.A(n_1), .B1(a[6]), .B2(n_2), .ZN(p_0[6]));
   AOI21_X1 i_6 (.A(n_55), .B1(a[7]), .B2(n_0), .ZN(p_0[7]));
   INV_X1 i_7 (.A(n_1), .ZN(n_0));
   NOR2_X1 i_8 (.A1(n_57), .A2(n_56), .ZN(n_1));
   INV_X1 i_9 (.A(n_3), .ZN(n_2));
   NOR2_X1 i_10 (.A1(a[5]), .A2(n_4), .ZN(n_3));
   INV_X1 i_11 (.A(n_5), .ZN(n_4));
   NOR2_X1 i_12 (.A1(a[4]), .A2(n_57), .ZN(n_5));
   AOI21_X1 i_13 (.A(n_11), .B1(a[8]), .B2(n_54), .ZN(p_0[8]));
   AOI21_X1 i_14 (.A(n_9), .B1(a[9]), .B2(n_10), .ZN(p_0[9]));
   AOI21_X1 i_15 (.A(n_7), .B1(a[10]), .B2(n_8), .ZN(p_0[10]));
   AOI21_X1 i_16 (.A(n_52), .B1(a[11]), .B2(n_6), .ZN(p_0[11]));
   INV_X1 i_17 (.A(n_7), .ZN(n_6));
   NOR2_X1 i_18 (.A1(n_54), .A2(n_53), .ZN(n_7));
   INV_X1 i_19 (.A(n_9), .ZN(n_8));
   NOR2_X1 i_20 (.A1(a[9]), .A2(n_10), .ZN(n_9));
   INV_X1 i_21 (.A(n_11), .ZN(n_10));
   NOR2_X1 i_22 (.A1(a[8]), .A2(n_54), .ZN(n_11));
   AOI21_X1 i_23 (.A(n_17), .B1(a[12]), .B2(n_51), .ZN(p_0[12]));
   AOI21_X1 i_24 (.A(n_15), .B1(a[13]), .B2(n_16), .ZN(p_0[13]));
   AOI21_X1 i_25 (.A(n_13), .B1(a[14]), .B2(n_14), .ZN(p_0[14]));
   AOI21_X1 i_26 (.A(n_49), .B1(a[15]), .B2(n_12), .ZN(p_0[15]));
   INV_X1 i_27 (.A(n_13), .ZN(n_12));
   NOR2_X1 i_28 (.A1(n_51), .A2(n_50), .ZN(n_13));
   INV_X1 i_29 (.A(n_15), .ZN(n_14));
   NOR2_X1 i_30 (.A1(a[13]), .A2(n_16), .ZN(n_15));
   INV_X1 i_31 (.A(n_17), .ZN(n_16));
   NOR2_X1 i_32 (.A1(a[12]), .A2(n_51), .ZN(n_17));
   AOI21_X1 i_33 (.A(n_23), .B1(a[16]), .B2(n_48), .ZN(p_0[16]));
   AOI21_X1 i_34 (.A(n_21), .B1(a[17]), .B2(n_22), .ZN(p_0[17]));
   AOI21_X1 i_35 (.A(n_19), .B1(a[18]), .B2(n_20), .ZN(p_0[18]));
   AOI21_X1 i_36 (.A(n_45), .B1(a[19]), .B2(n_18), .ZN(p_0[19]));
   INV_X1 i_37 (.A(n_19), .ZN(n_18));
   NOR2_X1 i_38 (.A1(n_48), .A2(n_46), .ZN(n_19));
   INV_X1 i_39 (.A(n_21), .ZN(n_20));
   NOR2_X1 i_40 (.A1(a[17]), .A2(n_22), .ZN(n_21));
   INV_X1 i_41 (.A(n_23), .ZN(n_22));
   NOR2_X1 i_42 (.A1(a[16]), .A2(n_48), .ZN(n_23));
   AOI21_X1 i_43 (.A(n_25), .B1(a[20]), .B2(n_44), .ZN(p_0[20]));
   AOI21_X1 i_44 (.A(n_27), .B1(a[21]), .B2(n_24), .ZN(p_0[21]));
   INV_X1 i_45 (.A(n_25), .ZN(n_24));
   NOR2_X1 i_46 (.A1(a[20]), .A2(n_44), .ZN(n_25));
   AOI21_X1 i_47 (.A(n_43), .B1(a[22]), .B2(n_26), .ZN(p_0[22]));
   INV_X1 i_48 (.A(n_27), .ZN(n_26));
   NOR3_X1 i_49 (.A1(a[21]), .A2(a[20]), .A3(n_44), .ZN(n_27));
   AOI21_X1 i_50 (.A(n_41), .B1(a[23]), .B2(n_42), .ZN(p_0[23]));
   AOI21_X1 i_51 (.A(n_29), .B1(a[24]), .B2(n_40), .ZN(p_0[24]));
   AOI21_X1 i_61 (.A(n_36), .B1(a[29]), .B2(n_33), .ZN(p_0[29]));
   INV_X1 i_62 (.A(n_34), .ZN(n_33));
   AOI21_X1 i_64 (.A(n_37), .B1(a[30]), .B2(n_35), .ZN(p_0[30]));
   INV_X1 i_65 (.A(n_36), .ZN(n_35));
   NOR3_X1 i_66 (.A1(a[29]), .A2(a[28]), .A3(n_38), .ZN(n_36));
   XNOR2_X1 i_67 (.A(a[31]), .B(n_37), .ZN(p_0[31]));
   NOR4_X1 i_68 (.A1(a[29]), .A2(a[28]), .A3(a[30]), .A4(n_38), .ZN(n_37));
   INV_X1 i_52 (.A(n_28), .ZN(n_29));
   NAND3_X1 i_53 (.A1(n_81), .A2(n_80), .A3(n_79), .ZN(n_46));
   NAND3_X1 i_54 (.A1(n_87), .A2(n_86), .A3(n_85), .ZN(n_50));
   NAND3_X1 i_55 (.A1(n_93), .A2(n_92), .A3(n_91), .ZN(n_53));
   NAND3_X1 i_56 (.A1(n_99), .A2(n_98), .A3(n_97), .ZN(n_56));
   INV_X1 i_57 (.A(n_59), .ZN(n_60));
   NAND2_X1 i_58 (.A1(n_62), .A2(n_103), .ZN(n_59));
   INV_X1 i_59 (.A(n_61), .ZN(n_62));
   NAND2_X1 i_60 (.A1(n_102), .A2(n_101), .ZN(n_61));
   AOI21_X1 i_63 (.A(n_31), .B1(n_28), .B2(a[25]), .ZN(p_0[25]));
   NAND2_X1 i_69 (.A1(n_41), .A2(n_30), .ZN(n_28));
   INV_X1 i_70 (.A(a[24]), .ZN(n_30));
   INV_X1 i_71 (.A(n_32), .ZN(n_31));
   AOI22_X1 i_72 (.A1(n_32), .A2(a[26]), .B1(n_41), .B2(n_69), .ZN(p_0[26]));
   NAND4_X1 i_73 (.A1(n_45), .A2(n_105), .A3(n_72), .A4(n_39), .ZN(n_32));
   INV_X1 i_74 (.A(n_47), .ZN(n_39));
   OR2_X1 i_75 (.A1(a[25]), .A2(a[24]), .ZN(n_47));
   INV_X1 i_76 (.A(n_44), .ZN(n_45));
   NAND4_X1 i_77 (.A1(n_55), .A2(n_89), .A3(n_83), .A4(n_77), .ZN(n_44));
   INV_X1 i_78 (.A(n_54), .ZN(n_55));
   NAND2_X1 i_79 (.A1(n_58), .A2(n_95), .ZN(n_54));
   AOI21_X1 i_80 (.A(n_64), .B1(n_63), .B2(a[27]), .ZN(p_0[27]));
   NAND2_X1 i_81 (.A1(n_41), .A2(n_69), .ZN(n_63));
   INV_X1 i_82 (.A(n_38), .ZN(n_64));
   NAND3_X1 i_83 (.A1(n_43), .A2(n_105), .A3(n_67), .ZN(n_38));
   NOR2_X1 i_84 (.A1(n_65), .A2(n_34), .ZN(p_0[28]));
   AOI21_X1 i_85 (.A(n_106), .B1(n_41), .B2(n_67), .ZN(n_65));
   INV_X1 i_86 (.A(n_40), .ZN(n_41));
   NAND4_X1 i_87 (.A1(n_49), .A2(n_105), .A3(n_77), .A4(n_72), .ZN(n_40));
   INV_X1 i_88 (.A(n_48), .ZN(n_49));
   NAND4_X1 i_89 (.A1(n_58), .A2(n_95), .A3(n_89), .A4(n_83), .ZN(n_48));
   INV_X1 i_90 (.A(n_66), .ZN(n_34));
   NAND4_X1 i_91 (.A1(n_43), .A2(n_106), .A3(n_105), .A4(n_67), .ZN(n_66));
   INV_X1 i_92 (.A(n_68), .ZN(n_67));
   NAND2_X1 i_93 (.A1(n_69), .A2(n_71), .ZN(n_68));
   INV_X1 i_94 (.A(n_70), .ZN(n_69));
   OR3_X1 i_95 (.A1(a[26]), .A2(a[25]), .A3(a[24]), .ZN(n_70));
   INV_X1 i_96 (.A(a[27]), .ZN(n_71));
   INV_X1 i_97 (.A(n_42), .ZN(n_43));
   NAND4_X1 i_98 (.A1(n_52), .A2(n_83), .A3(n_77), .A4(n_72), .ZN(n_42));
   INV_X1 i_99 (.A(n_73), .ZN(n_72));
   NAND3_X1 i_100 (.A1(n_76), .A2(n_75), .A3(n_74), .ZN(n_73));
   INV_X1 i_101 (.A(a[20]), .ZN(n_74));
   INV_X1 i_102 (.A(a[21]), .ZN(n_75));
   INV_X1 i_103 (.A(a[22]), .ZN(n_76));
   INV_X1 i_104 (.A(n_78), .ZN(n_77));
   NAND4_X1 i_105 (.A1(n_82), .A2(n_81), .A3(n_80), .A4(n_79), .ZN(n_78));
   INV_X1 i_106 (.A(a[16]), .ZN(n_79));
   INV_X1 i_107 (.A(a[17]), .ZN(n_80));
   INV_X1 i_108 (.A(a[18]), .ZN(n_81));
   INV_X1 i_109 (.A(a[19]), .ZN(n_82));
   INV_X1 i_110 (.A(n_84), .ZN(n_83));
   NAND4_X1 i_111 (.A1(n_88), .A2(n_87), .A3(n_86), .A4(n_85), .ZN(n_84));
   INV_X1 i_112 (.A(a[12]), .ZN(n_85));
   INV_X1 i_113 (.A(a[13]), .ZN(n_86));
   INV_X1 i_114 (.A(a[14]), .ZN(n_87));
   INV_X1 i_115 (.A(a[15]), .ZN(n_88));
   INV_X1 i_116 (.A(n_51), .ZN(n_52));
   NAND3_X1 i_117 (.A1(n_58), .A2(n_95), .A3(n_89), .ZN(n_51));
   INV_X1 i_118 (.A(n_90), .ZN(n_89));
   NAND4_X1 i_119 (.A1(n_94), .A2(n_93), .A3(n_92), .A4(n_91), .ZN(n_90));
   INV_X1 i_120 (.A(a[8]), .ZN(n_91));
   INV_X1 i_121 (.A(a[9]), .ZN(n_92));
   INV_X1 i_122 (.A(a[10]), .ZN(n_93));
   INV_X1 i_123 (.A(a[11]), .ZN(n_94));
   INV_X1 i_124 (.A(n_96), .ZN(n_95));
   NAND4_X1 i_125 (.A1(n_100), .A2(n_99), .A3(n_98), .A4(n_97), .ZN(n_96));
   INV_X1 i_126 (.A(a[4]), .ZN(n_97));
   INV_X1 i_127 (.A(a[5]), .ZN(n_98));
   INV_X1 i_128 (.A(a[6]), .ZN(n_99));
   INV_X1 i_129 (.A(a[7]), .ZN(n_100));
   INV_X1 i_130 (.A(n_57), .ZN(n_58));
   NAND4_X1 i_131 (.A1(n_104), .A2(n_103), .A3(n_102), .A4(n_101), .ZN(n_57));
   INV_X1 i_132 (.A(a[0]), .ZN(n_101));
   INV_X1 i_133 (.A(a[1]), .ZN(n_102));
   INV_X1 i_134 (.A(a[2]), .ZN(n_103));
   INV_X1 i_135 (.A(a[3]), .ZN(n_104));
   INV_X1 i_136 (.A(a[23]), .ZN(n_105));
   INV_X1 i_137 (.A(a[28]), .ZN(n_106));
endmodule

module datapath__0_2(b, p_0);
   input [31:0]b;
   output [31:0]p_0;

   AOI21_X1 i_35 (.A(n_19), .B1(b[18]), .B2(n_20), .ZN(p_0[18]));
   AOI21_X1 i_36 (.A(n_45), .B1(b[19]), .B2(n_18), .ZN(p_0[19]));
   INV_X1 i_37 (.A(n_19), .ZN(n_18));
   NOR2_X1 i_38 (.A1(n_48), .A2(n_46), .ZN(n_19));
   INV_X1 i_39 (.A(n_21), .ZN(n_20));
   AOI21_X1 i_43 (.A(n_25), .B1(b[20]), .B2(n_44), .ZN(p_0[20]));
   AOI21_X1 i_44 (.A(n_27), .B1(b[21]), .B2(n_24), .ZN(p_0[21]));
   INV_X1 i_45 (.A(n_25), .ZN(n_24));
   NOR2_X1 i_46 (.A1(b[20]), .A2(n_44), .ZN(n_25));
   AOI21_X1 i_47 (.A(n_43), .B1(b[22]), .B2(n_26), .ZN(p_0[22]));
   INV_X1 i_48 (.A(n_27), .ZN(n_26));
   NOR3_X1 i_49 (.A1(b[21]), .A2(b[20]), .A3(n_44), .ZN(n_27));
   AOI21_X1 i_50 (.A(n_41), .B1(b[23]), .B2(n_42), .ZN(p_0[23]));
   AOI21_X1 i_51 (.A(n_29), .B1(b[24]), .B2(n_40), .ZN(p_0[24]));
   INV_X1 i_52 (.A(n_28), .ZN(p_0[25]));
   OAI21_X1 i_53 (.A(n_30), .B1(n_63), .B2(n_29), .ZN(n_28));
   NOR2_X1 i_54 (.A1(b[24]), .A2(n_40), .ZN(n_29));
   AOI21_X1 i_55 (.A(n_32), .B1(b[26]), .B2(n_30), .ZN(p_0[26]));
   OR3_X1 i_56 (.A1(b[25]), .A2(b[24]), .A3(n_40), .ZN(n_30));
   AOI21_X1 i_57 (.A(n_39), .B1(b[27]), .B2(n_31), .ZN(p_0[27]));
   INV_X1 i_58 (.A(n_32), .ZN(n_31));
   NOR2_X1 i_59 (.A1(n_47), .A2(n_40), .ZN(n_32));
   AOI21_X1 i_60 (.A(n_34), .B1(b[28]), .B2(n_38), .ZN(p_0[28]));
   AOI21_X1 i_61 (.A(n_36), .B1(b[29]), .B2(n_33), .ZN(p_0[29]));
   INV_X1 i_62 (.A(n_34), .ZN(n_33));
   NOR2_X1 i_63 (.A1(b[28]), .A2(n_38), .ZN(n_34));
   AOI21_X1 i_64 (.A(n_37), .B1(b[30]), .B2(n_35), .ZN(p_0[30]));
   INV_X1 i_65 (.A(n_36), .ZN(n_35));
   NOR3_X1 i_66 (.A1(b[29]), .A2(b[28]), .A3(n_38), .ZN(n_36));
   XNOR2_X1 i_67 (.A(b[31]), .B(n_37), .ZN(p_0[31]));
   NOR4_X1 i_68 (.A1(b[29]), .A2(b[28]), .A3(b[30]), .A4(n_38), .ZN(n_37));
   INV_X1 i_69 (.A(n_39), .ZN(n_38));
   NOR3_X1 i_70 (.A1(b[27]), .A2(n_47), .A3(n_40), .ZN(n_39));
   INV_X1 i_71 (.A(n_41), .ZN(n_40));
   NOR2_X1 i_72 (.A1(b[23]), .A2(n_42), .ZN(n_41));
   INV_X1 i_73 (.A(n_43), .ZN(n_42));
   NOR4_X1 i_74 (.A1(b[22]), .A2(b[21]), .A3(b[20]), .A4(n_44), .ZN(n_43));
   INV_X1 i_75 (.A(n_45), .ZN(n_44));
   NOR3_X1 i_76 (.A1(b[19]), .A2(n_46), .A3(n_48), .ZN(n_45));
   OR3_X1 i_77 (.A1(b[18]), .A2(b[16]), .A3(b[17]), .ZN(n_46));
   OR3_X1 i_78 (.A1(b[26]), .A2(b[25]), .A3(b[24]), .ZN(n_47));
   INV_X1 i_94 (.A(b[25]), .ZN(n_63));
   INV_X1 i_0 (.A(n_4), .ZN(n_15));
   INV_X1 i_1 (.A(n_52), .ZN(n_9));
   INV_X1 i_2 (.A(n_0), .ZN(n_3));
   NAND2_X1 i_3 (.A1(n_5), .A2(n_1), .ZN(n_0));
   XNOR2_X1 i_4 (.A(n_17), .B(n_1), .ZN(p_0[5]));
   INV_X1 i_5 (.A(b[5]), .ZN(n_1));
   OR2_X1 i_6 (.A1(n_50), .A2(b[15]), .ZN(n_2));
   OR2_X1 i_7 (.A1(n_61), .A2(b[13]), .ZN(n_4));
   INV_X1 i_8 (.A(n_72), .ZN(n_21));
   INV_X1 i_9 (.A(n_17), .ZN(n_5));
   INV_X1 i_10 (.A(n_6), .ZN(p_0[1]));
   NAND2_X1 i_11 (.A1(n_11), .A2(n_7), .ZN(n_6));
   NAND2_X1 i_12 (.A1(b[1]), .A2(b[0]), .ZN(n_7));
   INV_X1 i_13 (.A(n_8), .ZN(p_0[2]));
   NAND2_X1 i_14 (.A1(n_10), .A2(n_92), .ZN(n_8));
   NAND2_X1 i_15 (.A1(n_11), .A2(b[2]), .ZN(n_10));
   NAND2_X1 i_16 (.A1(n_94), .A2(n_93), .ZN(n_11));
   INV_X1 i_17 (.A(n_12), .ZN(p_0[3]));
   NAND2_X1 i_18 (.A1(n_90), .A2(n_13), .ZN(n_12));
   NAND2_X1 i_19 (.A1(n_92), .A2(b[3]), .ZN(n_13));
   INV_X1 i_20 (.A(n_14), .ZN(p_0[4]));
   NAND2_X1 i_21 (.A1(n_17), .A2(n_16), .ZN(n_14));
   NAND2_X1 i_22 (.A1(n_90), .A2(b[4]), .ZN(n_16));
   NAND2_X1 i_23 (.A1(n_89), .A2(n_86), .ZN(n_17));
   AOI22_X1 i_24 (.A1(n_22), .A2(b[6]), .B1(n_89), .B2(n_49), .ZN(p_0[6]));
   INV_X1 i_25 (.A(n_3), .ZN(n_22));
   AOI21_X1 i_26 (.A(n_81), .B1(b[7]), .B2(n_23), .ZN(p_0[7]));
   NAND2_X1 i_27 (.A1(n_89), .A2(n_49), .ZN(n_23));
   INV_X1 i_28 (.A(n_85), .ZN(n_49));
   XNOR2_X1 i_29 (.A(n_82), .B(n_77), .ZN(p_0[8]));
   INV_X1 i_30 (.A(n_51), .ZN(p_0[9]));
   NAND2_X1 i_31 (.A1(n_53), .A2(n_52), .ZN(n_51));
   NAND3_X1 i_32 (.A1(n_81), .A2(n_78), .A3(n_77), .ZN(n_52));
   OAI21_X1 i_33 (.A(b[9]), .B1(n_82), .B2(b[8]), .ZN(n_53));
   AOI21_X1 i_34 (.A(n_56), .B1(n_54), .B2(b[10]), .ZN(p_0[10]));
   INV_X1 i_40 (.A(n_9), .ZN(n_54));
   INV_X1 i_41 (.A(n_55), .ZN(p_0[11]));
   OAI21_X1 i_42 (.A(n_74), .B1(n_56), .B2(n_80), .ZN(n_55));
   INV_X1 i_79 (.A(n_57), .ZN(n_56));
   NAND4_X1 i_80 (.A1(n_81), .A2(n_79), .A3(n_78), .A4(n_77), .ZN(n_57));
   INV_X1 i_81 (.A(n_58), .ZN(p_0[12]));
   NAND2_X1 i_82 (.A1(n_61), .A2(n_59), .ZN(n_58));
   NAND2_X1 i_83 (.A1(n_74), .A2(b[12]), .ZN(n_59));
   INV_X1 i_84 (.A(n_60), .ZN(p_0[13]));
   XNOR2_X1 i_85 (.A(n_61), .B(b[13]), .ZN(n_60));
   NAND2_X1 i_86 (.A1(n_73), .A2(n_62), .ZN(n_61));
   INV_X1 i_87 (.A(b[12]), .ZN(n_62));
   AOI21_X1 i_88 (.A(n_64), .B1(n_65), .B2(b[14]), .ZN(p_0[14]));
   INV_X1 i_89 (.A(n_66), .ZN(n_64));
   INV_X1 i_90 (.A(n_15), .ZN(n_65));
   AOI22_X1 i_91 (.A1(n_97), .A2(n_73), .B1(b[15]), .B2(n_66), .ZN(p_0[15]));
   OR2_X1 i_92 (.A1(n_74), .A2(n_50), .ZN(n_66));
   OR3_X1 i_93 (.A1(b[14]), .A2(b[13]), .A3(b[12]), .ZN(n_50));
   INV_X1 i_95 (.A(n_67), .ZN(p_0[16]));
   NAND2_X1 i_96 (.A1(n_68), .A2(n_71), .ZN(n_67));
   NAND2_X1 i_97 (.A1(n_48), .A2(b[16]), .ZN(n_68));
   NAND2_X1 i_98 (.A1(n_97), .A2(n_73), .ZN(n_48));
   INV_X1 i_99 (.A(n_69), .ZN(p_0[17]));
   NAND2_X1 i_100 (.A1(n_70), .A2(n_72), .ZN(n_69));
   NAND2_X1 i_101 (.A1(n_71), .A2(b[17]), .ZN(n_70));
   NAND3_X1 i_102 (.A1(n_97), .A2(n_98), .A3(n_73), .ZN(n_71));
   NAND4_X1 i_103 (.A1(n_97), .A2(n_99), .A3(n_98), .A4(n_73), .ZN(n_72));
   INV_X1 i_104 (.A(n_74), .ZN(n_73));
   NAND2_X1 i_105 (.A1(n_81), .A2(n_75), .ZN(n_74));
   INV_X1 i_106 (.A(n_76), .ZN(n_75));
   NAND4_X1 i_107 (.A1(n_80), .A2(n_79), .A3(n_78), .A4(n_77), .ZN(n_76));
   INV_X1 i_108 (.A(b[8]), .ZN(n_77));
   INV_X1 i_109 (.A(b[9]), .ZN(n_78));
   INV_X1 i_110 (.A(b[10]), .ZN(n_79));
   INV_X1 i_111 (.A(b[11]), .ZN(n_80));
   INV_X1 i_112 (.A(n_82), .ZN(n_81));
   NAND2_X1 i_113 (.A1(n_83), .A2(n_89), .ZN(n_82));
   INV_X1 i_114 (.A(n_84), .ZN(n_83));
   OR2_X1 i_115 (.A1(n_85), .A2(b[7]), .ZN(n_84));
   NAND3_X1 i_116 (.A1(n_88), .A2(n_87), .A3(n_86), .ZN(n_85));
   INV_X1 i_117 (.A(b[4]), .ZN(n_86));
   INV_X1 i_118 (.A(b[5]), .ZN(n_87));
   INV_X1 i_119 (.A(b[6]), .ZN(n_88));
   INV_X1 i_120 (.A(n_90), .ZN(n_89));
   NAND2_X1 i_121 (.A1(n_91), .A2(n_96), .ZN(n_90));
   INV_X1 i_122 (.A(n_92), .ZN(n_91));
   NAND3_X1 i_123 (.A1(n_95), .A2(n_94), .A3(n_93), .ZN(n_92));
   INV_X1 i_124 (.A(b[0]), .ZN(n_93));
   INV_X1 i_125 (.A(b[1]), .ZN(n_94));
   INV_X1 i_126 (.A(b[2]), .ZN(n_95));
   INV_X1 i_127 (.A(b[3]), .ZN(n_96));
   INV_X1 i_128 (.A(n_2), .ZN(n_97));
   INV_X1 i_129 (.A(b[16]), .ZN(n_98));
   INV_X1 i_130 (.A(b[17]), .ZN(n_99));
endmodule

module datapath__0_6(p_0, Accumulator, Accumulator1);
   input [31:0]p_0;
   input [31:0]Accumulator;
   output [31:0]Accumulator1;

   INV_X1 i_0 (.A(n_0), .ZN(Accumulator1[0]));
   OAI21_X1 i_1 (.A(n_159), .B1(p_0[0]), .B2(Accumulator[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_159), .B(n_1), .Z(Accumulator1[1]));
   OAI21_X1 i_3 (.A(n_158), .B1(p_0[1]), .B2(Accumulator[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_157), .B(n_2), .ZN(Accumulator1[2]));
   OAI21_X1 i_5 (.A(n_162), .B1(p_0[2]), .B2(Accumulator[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_156), .B(n_3), .Z(Accumulator1[3]));
   OAI21_X1 i_7 (.A(n_163), .B1(n_168), .B2(n_165), .ZN(n_3));
   XOR2_X1 i_8 (.A(n_154), .B(n_10), .Z(Accumulator1[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(Accumulator1[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(Accumulator1[6]));
   NOR2_X1 i_11 (.A1(n_151), .A2(n_142), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(Accumulator1[7]));
   OAI22_X1 i_13 (.A1(p_0[6]), .A2(Accumulator[6]), .B1(n_142), .B2(n_7), 
      .ZN(n_5));
   AOI21_X1 i_14 (.A(n_152), .B1(p_0[5]), .B2(Accumulator[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_152), .B1(n_146), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_149), .B1(n_154), .B2(n_147), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_147), .B1(p_0[4]), .B2(Accumulator[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_153), .A2(n_144), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_140), .B(n_18), .ZN(Accumulator1[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(Accumulator1[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(Accumulator1[10]));
   NOR2_X1 i_23 (.A1(n_137), .A2(n_128), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(Accumulator1[11]));
   OAI22_X1 i_25 (.A1(p_0[10]), .A2(Accumulator[10]), .B1(n_128), .B2(n_15), 
      .ZN(n_13));
   AOI21_X1 i_26 (.A(n_138), .B1(p_0[9]), .B2(Accumulator[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_138), .B1(n_132), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_135), .B1(n_140), .B2(n_133), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_135), .B1(p_0[8]), .B2(Accumulator[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_139), .A2(n_130), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_126), .B(n_26), .Z(Accumulator1[12]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(Accumulator1[13]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(Accumulator1[14]));
   NOR2_X1 i_35 (.A1(n_123), .A2(n_114), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(Accumulator1[15]));
   OAI22_X1 i_37 (.A1(p_0[14]), .A2(Accumulator[14]), .B1(n_114), .B2(n_23), 
      .ZN(n_21));
   AOI21_X1 i_38 (.A(n_124), .B1(p_0[13]), .B2(Accumulator[13]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_124), .B1(n_118), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_121), .B1(n_126), .B2(n_119), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_119), .B1(p_0[12]), .B2(Accumulator[12]), .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_125), .A2(n_116), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_112), .B(n_34), .Z(Accumulator1[16]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(Accumulator1[17]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(Accumulator1[18]));
   NOR2_X1 i_47 (.A1(n_109), .A2(n_100), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(Accumulator1[19]));
   OAI22_X1 i_49 (.A1(p_0[18]), .A2(Accumulator[18]), .B1(n_100), .B2(n_31), 
      .ZN(n_29));
   AOI21_X1 i_50 (.A(n_110), .B1(p_0[17]), .B2(Accumulator[17]), .ZN(n_30));
   AOI21_X1 i_51 (.A(n_110), .B1(n_104), .B2(n_32), .ZN(n_31));
   INV_X1 i_52 (.A(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_107), .B1(n_112), .B2(n_105), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_105), .B1(p_0[16]), .B2(Accumulator[16]), .ZN(n_34));
   NOR2_X1 i_55 (.A1(n_111), .A2(n_102), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_98), .B(n_42), .Z(Accumulator1[20]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(Accumulator1[21]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(Accumulator1[22]));
   NOR2_X1 i_59 (.A1(n_87), .A2(n_77), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(Accumulator1[23]));
   OAI21_X1 i_61 (.A(n_86), .B1(n_77), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_89), .A2(n_79), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_88), .B1(n_79), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_84), .B1(n_98), .B2(n_81), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_81), .B1(p_0[20]), .B2(Accumulator[20]), .ZN(n_42));
   AOI21_X1 i_67 (.A(n_91), .B1(p_0[23]), .B2(Accumulator[23]), .ZN(n_43));
   XNOR2_X1 i_68 (.A(n_52), .B(n_51), .ZN(Accumulator1[24]));
   OAI21_X1 i_79 (.A(n_74), .B1(p_0[24]), .B2(Accumulator[24]), .ZN(n_51));
   XNOR2_X1 i_82 (.A(n_66), .B(n_65), .ZN(Accumulator1[28]));
   AOI22_X1 i_83 (.A1(n_63), .A2(n_59), .B1(n_64), .B2(n_58), .ZN(
      Accumulator1[29]));
   OAI21_X1 i_91 (.A(n_60), .B1(n_170), .B2(n_167), .ZN(n_59));
   NAND2_X1 i_106 (.A1(p_0[24]), .A2(Accumulator[24]), .ZN(n_74));
   INV_X1 i_111 (.A(n_80), .ZN(n_79));
   NOR2_X1 i_116 (.A1(p_0[20]), .A2(Accumulator[20]), .ZN(n_84));
   NOR2_X1 i_119 (.A1(p_0[22]), .A2(Accumulator[22]), .ZN(n_87));
   NOR2_X1 i_121 (.A1(p_0[21]), .A2(Accumulator[21]), .ZN(n_89));
   NOR2_X1 i_131 (.A1(n_111), .A2(n_101), .ZN(n_99));
   INV_X1 i_132 (.A(n_101), .ZN(n_100));
   NAND2_X1 i_133 (.A1(p_0[18]), .A2(Accumulator[18]), .ZN(n_101));
   AND2_X1 i_134 (.A1(p_0[19]), .A2(Accumulator[19]), .ZN(n_102));
   AOI21_X1 i_135 (.A(n_108), .B1(n_105), .B2(n_104), .ZN(n_103));
   NAND2_X1 i_136 (.A1(p_0[17]), .A2(Accumulator[17]), .ZN(n_104));
   NAND2_X1 i_137 (.A1(p_0[16]), .A2(Accumulator[16]), .ZN(n_105));
   NOR3_X1 i_138 (.A1(n_108), .A2(n_107), .A3(n_112), .ZN(n_106));
   NOR2_X1 i_139 (.A1(p_0[16]), .A2(Accumulator[16]), .ZN(n_107));
   OR3_X1 i_140 (.A1(n_111), .A2(n_109), .A3(n_110), .ZN(n_108));
   NOR2_X1 i_141 (.A1(p_0[18]), .A2(Accumulator[18]), .ZN(n_109));
   NOR2_X1 i_142 (.A1(p_0[17]), .A2(Accumulator[17]), .ZN(n_110));
   NOR2_X1 i_143 (.A1(p_0[19]), .A2(Accumulator[19]), .ZN(n_111));
   NOR4_X1 i_144 (.A1(n_116), .A2(n_113), .A3(n_117), .A4(n_120), .ZN(n_112));
   NOR2_X1 i_145 (.A1(n_125), .A2(n_115), .ZN(n_113));
   INV_X1 i_146 (.A(n_115), .ZN(n_114));
   NAND2_X1 i_147 (.A1(p_0[14]), .A2(Accumulator[14]), .ZN(n_115));
   AND2_X1 i_148 (.A1(p_0[15]), .A2(Accumulator[15]), .ZN(n_116));
   AOI21_X1 i_149 (.A(n_122), .B1(n_119), .B2(n_118), .ZN(n_117));
   NAND2_X1 i_150 (.A1(p_0[13]), .A2(Accumulator[13]), .ZN(n_118));
   NAND2_X1 i_151 (.A1(p_0[12]), .A2(Accumulator[12]), .ZN(n_119));
   NOR3_X1 i_152 (.A1(n_122), .A2(n_121), .A3(n_126), .ZN(n_120));
   NOR2_X1 i_153 (.A1(p_0[12]), .A2(Accumulator[12]), .ZN(n_121));
   OR3_X1 i_154 (.A1(n_125), .A2(n_123), .A3(n_124), .ZN(n_122));
   NOR2_X1 i_155 (.A1(p_0[14]), .A2(Accumulator[14]), .ZN(n_123));
   NOR2_X1 i_156 (.A1(p_0[13]), .A2(Accumulator[13]), .ZN(n_124));
   NOR2_X1 i_157 (.A1(p_0[15]), .A2(Accumulator[15]), .ZN(n_125));
   NOR4_X1 i_158 (.A1(n_130), .A2(n_127), .A3(n_131), .A4(n_134), .ZN(n_126));
   NOR2_X1 i_159 (.A1(n_139), .A2(n_129), .ZN(n_127));
   INV_X1 i_160 (.A(n_129), .ZN(n_128));
   NAND2_X1 i_161 (.A1(p_0[10]), .A2(Accumulator[10]), .ZN(n_129));
   AND2_X1 i_162 (.A1(p_0[11]), .A2(Accumulator[11]), .ZN(n_130));
   AOI21_X1 i_163 (.A(n_136), .B1(n_133), .B2(n_132), .ZN(n_131));
   NAND2_X1 i_164 (.A1(p_0[9]), .A2(Accumulator[9]), .ZN(n_132));
   NAND2_X1 i_165 (.A1(p_0[8]), .A2(Accumulator[8]), .ZN(n_133));
   NOR3_X1 i_166 (.A1(n_136), .A2(n_135), .A3(n_140), .ZN(n_134));
   NOR2_X1 i_167 (.A1(p_0[8]), .A2(Accumulator[8]), .ZN(n_135));
   OR3_X1 i_168 (.A1(n_139), .A2(n_137), .A3(n_138), .ZN(n_136));
   NOR2_X1 i_169 (.A1(p_0[10]), .A2(Accumulator[10]), .ZN(n_137));
   NOR2_X1 i_170 (.A1(p_0[9]), .A2(Accumulator[9]), .ZN(n_138));
   NOR2_X1 i_171 (.A1(p_0[11]), .A2(Accumulator[11]), .ZN(n_139));
   NOR4_X1 i_172 (.A1(n_144), .A2(n_141), .A3(n_145), .A4(n_148), .ZN(n_140));
   NOR2_X1 i_173 (.A1(n_153), .A2(n_143), .ZN(n_141));
   INV_X1 i_174 (.A(n_143), .ZN(n_142));
   NAND2_X1 i_175 (.A1(p_0[6]), .A2(Accumulator[6]), .ZN(n_143));
   AND2_X1 i_176 (.A1(p_0[7]), .A2(Accumulator[7]), .ZN(n_144));
   AOI21_X1 i_177 (.A(n_150), .B1(n_147), .B2(n_146), .ZN(n_145));
   NAND2_X1 i_178 (.A1(p_0[5]), .A2(Accumulator[5]), .ZN(n_146));
   NAND2_X1 i_179 (.A1(p_0[4]), .A2(Accumulator[4]), .ZN(n_147));
   NOR3_X1 i_180 (.A1(n_150), .A2(n_149), .A3(n_154), .ZN(n_148));
   NOR2_X1 i_181 (.A1(p_0[4]), .A2(Accumulator[4]), .ZN(n_149));
   OR3_X1 i_182 (.A1(n_153), .A2(n_151), .A3(n_152), .ZN(n_150));
   NOR2_X1 i_183 (.A1(p_0[6]), .A2(Accumulator[6]), .ZN(n_151));
   NOR2_X1 i_184 (.A1(p_0[5]), .A2(Accumulator[5]), .ZN(n_152));
   NOR2_X1 i_185 (.A1(p_0[7]), .A2(Accumulator[7]), .ZN(n_153));
   NAND2_X1 i_186 (.A1(n_163), .A2(n_155), .ZN(n_154));
   OAI21_X1 i_187 (.A(n_156), .B1(n_168), .B2(n_165), .ZN(n_155));
   OAI22_X1 i_188 (.A1(p_0[2]), .A2(Accumulator[2]), .B1(n_161), .B2(n_157), 
      .ZN(n_156));
   AOI21_X1 i_189 (.A(n_160), .B1(n_159), .B2(n_158), .ZN(n_157));
   NAND2_X1 i_190 (.A1(p_0[1]), .A2(Accumulator[1]), .ZN(n_158));
   NAND2_X1 i_191 (.A1(p_0[0]), .A2(Accumulator[0]), .ZN(n_159));
   NOR2_X1 i_192 (.A1(p_0[1]), .A2(Accumulator[1]), .ZN(n_160));
   INV_X1 i_193 (.A(n_162), .ZN(n_161));
   NAND2_X1 i_194 (.A1(p_0[2]), .A2(Accumulator[2]), .ZN(n_162));
   NAND2_X1 i_195 (.A1(n_168), .A2(n_165), .ZN(n_163));
   INV_X1 i_197 (.A(Accumulator[3]), .ZN(n_165));
   INV_X1 i_198 (.A(Accumulator[27]), .ZN(n_166));
   INV_X1 i_199 (.A(Accumulator[29]), .ZN(n_167));
   INV_X1 i_200 (.A(p_0[3]), .ZN(n_168));
   INV_X1 i_201 (.A(p_0[27]), .ZN(n_169));
   INV_X1 i_202 (.A(p_0[29]), .ZN(n_170));
   INV_X1 i_69 (.A(n_59), .ZN(n_58));
   INV_X1 i_70 (.A(n_64), .ZN(n_63));
   INV_X1 i_71 (.A(n_44), .ZN(n_65));
   NAND2_X1 i_72 (.A1(n_45), .A2(n_185), .ZN(n_44));
   INV_X1 i_73 (.A(n_184), .ZN(n_45));
   INV_X1 i_74 (.A(n_89), .ZN(n_88));
   INV_X1 i_75 (.A(n_87), .ZN(n_86));
   XNOR2_X1 i_76 (.A(n_46), .B(n_53), .ZN(Accumulator1[25]));
   NAND2_X1 i_77 (.A1(n_55), .A2(n_95), .ZN(n_46));
   XNOR2_X1 i_78 (.A(n_49), .B(n_47), .ZN(Accumulator1[26]));
   NAND2_X1 i_80 (.A1(n_57), .A2(n_92), .ZN(n_47));
   XOR2_X1 i_81 (.A(n_61), .B(n_48), .Z(Accumulator1[27]));
   OAI21_X1 i_84 (.A(n_57), .B1(n_49), .B2(n_56), .ZN(n_48));
   NAND2_X1 i_85 (.A1(n_50), .A2(n_95), .ZN(n_49));
   NAND2_X1 i_86 (.A1(n_53), .A2(n_55), .ZN(n_50));
   OAI21_X1 i_87 (.A(n_96), .B1(n_74), .B2(n_54), .ZN(n_53));
   NOR2_X1 i_88 (.A1(p_0[24]), .A2(Accumulator[24]), .ZN(n_54));
   NAND2_X1 i_89 (.A1(n_181), .A2(n_180), .ZN(n_55));
   INV_X1 i_90 (.A(n_92), .ZN(n_56));
   INV_X1 i_92 (.A(n_179), .ZN(n_57));
   NAND2_X1 i_93 (.A1(n_182), .A2(n_62), .ZN(n_61));
   NAND2_X1 i_94 (.A1(p_0[27]), .A2(Accumulator[27]), .ZN(n_62));
   INV_X1 i_95 (.A(n_67), .ZN(Accumulator1[30]));
   XOR2_X1 i_96 (.A(n_70), .B(n_68), .Z(n_67));
   NAND2_X1 i_97 (.A1(n_82), .A2(n_69), .ZN(n_68));
   NAND2_X1 i_98 (.A1(p_0[29]), .A2(Accumulator[29]), .ZN(n_69));
   NAND2_X1 i_99 (.A1(n_187), .A2(n_78), .ZN(n_70));
   NAND2_X1 i_100 (.A1(n_71), .A2(n_73), .ZN(Accumulator1[31]));
   NAND2_X1 i_101 (.A1(n_72), .A2(p_0[31]), .ZN(n_71));
   NAND2_X1 i_102 (.A1(n_75), .A2(n_187), .ZN(n_72));
   NAND3_X1 i_103 (.A1(n_75), .A2(n_188), .A3(n_187), .ZN(n_73));
   NAND2_X1 i_104 (.A1(n_186), .A2(n_76), .ZN(n_75));
   AND2_X1 i_105 (.A1(n_82), .A2(n_78), .ZN(n_76));
   NAND2_X1 i_107 (.A1(p_0[30]), .A2(Accumulator[30]), .ZN(n_78));
   NAND2_X1 i_108 (.A1(n_60), .A2(n_64), .ZN(n_82));
   OAI21_X1 i_109 (.A(n_185), .B1(n_66), .B2(n_184), .ZN(n_64));
   INV_X1 i_110 (.A(n_83), .ZN(n_66));
   OAI211_X1 i_112 (.A(n_93), .B(n_85), .C1(n_177), .C2(n_96), .ZN(n_83));
   INV_X1 i_113 (.A(n_90), .ZN(n_85));
   OAI22_X1 i_114 (.A1(n_183), .A2(n_92), .B1(n_169), .B2(n_166), .ZN(n_90));
   NAND2_X1 i_115 (.A1(p_0[26]), .A2(Accumulator[26]), .ZN(n_92));
   NAND3_X1 i_117 (.A1(n_182), .A2(n_178), .A3(n_94), .ZN(n_93));
   NAND2_X1 i_118 (.A1(n_95), .A2(n_74), .ZN(n_94));
   NAND2_X1 i_120 (.A1(p_0[25]), .A2(Accumulator[25]), .ZN(n_95));
   OAI21_X1 i_122 (.A(n_52), .B1(p_0[24]), .B2(Accumulator[24]), .ZN(n_96));
   NAND4_X1 i_123 (.A1(n_174), .A2(n_172), .A3(n_171), .A4(n_97), .ZN(n_52));
   OAI21_X1 i_124 (.A(n_77), .B1(p_0[23]), .B2(Accumulator[23]), .ZN(n_97));
   INV_X1 i_125 (.A(n_164), .ZN(n_77));
   NAND2_X1 i_126 (.A1(p_0[22]), .A2(Accumulator[22]), .ZN(n_164));
   NAND2_X1 i_127 (.A1(p_0[23]), .A2(Accumulator[23]), .ZN(n_171));
   NAND2_X1 i_128 (.A1(n_176), .A2(n_173), .ZN(n_172));
   NAND2_X1 i_129 (.A1(n_80), .A2(n_81), .ZN(n_173));
   NAND2_X1 i_130 (.A1(p_0[21]), .A2(Accumulator[21]), .ZN(n_80));
   NAND2_X1 i_196 (.A1(p_0[20]), .A2(Accumulator[20]), .ZN(n_81));
   NAND2_X1 i_203 (.A1(n_176), .A2(n_175), .ZN(n_174));
   NOR2_X1 i_204 (.A1(n_98), .A2(n_84), .ZN(n_175));
   NOR4_X1 i_205 (.A1(n_106), .A2(n_103), .A3(n_102), .A4(n_99), .ZN(n_98));
   NOR3_X1 i_206 (.A1(n_91), .A2(n_87), .A3(n_89), .ZN(n_176));
   NOR2_X1 i_207 (.A1(p_0[23]), .A2(Accumulator[23]), .ZN(n_91));
   NAND2_X1 i_208 (.A1(n_182), .A2(n_178), .ZN(n_177));
   AOI21_X1 i_209 (.A(n_179), .B1(n_181), .B2(n_180), .ZN(n_178));
   NOR2_X1 i_210 (.A1(p_0[26]), .A2(Accumulator[26]), .ZN(n_179));
   INV_X1 i_211 (.A(Accumulator[25]), .ZN(n_180));
   INV_X1 i_212 (.A(p_0[25]), .ZN(n_181));
   INV_X1 i_213 (.A(n_183), .ZN(n_182));
   NOR2_X1 i_214 (.A1(p_0[27]), .A2(Accumulator[27]), .ZN(n_183));
   NOR2_X1 i_215 (.A1(p_0[28]), .A2(Accumulator[28]), .ZN(n_184));
   NAND2_X1 i_216 (.A1(p_0[28]), .A2(Accumulator[28]), .ZN(n_185));
   NAND2_X1 i_217 (.A1(n_59), .A2(n_60), .ZN(n_186));
   NAND2_X1 i_218 (.A1(n_170), .A2(n_167), .ZN(n_60));
   OR2_X1 i_219 (.A1(p_0[30]), .A2(Accumulator[30]), .ZN(n_187));
   INV_X1 i_220 (.A(p_0[31]), .ZN(n_188));
endmodule

module datapath__0_9(p_0, p_1);
   input [63:0]p_0;
   output [63:0]p_1;

   AOI21_X1 i_0 (.A(n_127), .B1(p_0[1]), .B2(p_0[0]), .ZN(p_1[1]));
   AOI21_X1 i_1 (.A(n_125), .B1(p_0[2]), .B2(n_126), .ZN(p_1[2]));
   AOI21_X1 i_2 (.A(n_123), .B1(p_0[3]), .B2(n_124), .ZN(p_1[3]));
   AOI21_X1 i_3 (.A(n_5), .B1(p_0[4]), .B2(n_122), .ZN(p_1[4]));
   AOI21_X1 i_4 (.A(n_3), .B1(p_0[5]), .B2(n_4), .ZN(p_1[5]));
   AOI21_X1 i_5 (.A(n_1), .B1(p_0[6]), .B2(n_2), .ZN(p_1[6]));
   AOI21_X1 i_6 (.A(n_120), .B1(p_0[7]), .B2(n_0), .ZN(p_1[7]));
   INV_X1 i_7 (.A(n_1), .ZN(n_0));
   NOR2_X1 i_8 (.A1(n_122), .A2(n_121), .ZN(n_1));
   INV_X1 i_9 (.A(n_3), .ZN(n_2));
   NOR2_X1 i_10 (.A1(p_0[5]), .A2(n_4), .ZN(n_3));
   INV_X1 i_11 (.A(n_5), .ZN(n_4));
   NOR2_X1 i_12 (.A1(p_0[4]), .A2(n_122), .ZN(n_5));
   AOI21_X1 i_13 (.A(n_11), .B1(p_0[8]), .B2(n_119), .ZN(p_1[8]));
   AOI21_X1 i_14 (.A(n_9), .B1(p_0[9]), .B2(n_10), .ZN(p_1[9]));
   AOI21_X1 i_15 (.A(n_7), .B1(p_0[10]), .B2(n_8), .ZN(p_1[10]));
   AOI21_X1 i_16 (.A(n_117), .B1(p_0[11]), .B2(n_6), .ZN(p_1[11]));
   INV_X1 i_17 (.A(n_7), .ZN(n_6));
   NOR2_X1 i_18 (.A1(n_119), .A2(n_118), .ZN(n_7));
   INV_X1 i_19 (.A(n_9), .ZN(n_8));
   NOR2_X1 i_20 (.A1(p_0[9]), .A2(n_10), .ZN(n_9));
   INV_X1 i_21 (.A(n_11), .ZN(n_10));
   NOR2_X1 i_22 (.A1(p_0[8]), .A2(n_119), .ZN(n_11));
   AOI21_X1 i_23 (.A(n_17), .B1(p_0[12]), .B2(n_116), .ZN(p_1[12]));
   AOI21_X1 i_24 (.A(n_15), .B1(p_0[13]), .B2(n_16), .ZN(p_1[13]));
   AOI21_X1 i_25 (.A(n_13), .B1(p_0[14]), .B2(n_14), .ZN(p_1[14]));
   AOI21_X1 i_26 (.A(n_114), .B1(p_0[15]), .B2(n_12), .ZN(p_1[15]));
   INV_X1 i_27 (.A(n_13), .ZN(n_12));
   NOR2_X1 i_28 (.A1(n_116), .A2(n_115), .ZN(n_13));
   INV_X1 i_29 (.A(n_15), .ZN(n_14));
   NOR2_X1 i_30 (.A1(p_0[13]), .A2(n_16), .ZN(n_15));
   INV_X1 i_31 (.A(n_17), .ZN(n_16));
   NOR2_X1 i_32 (.A1(p_0[12]), .A2(n_116), .ZN(n_17));
   AOI21_X1 i_33 (.A(n_112), .B1(p_0[16]), .B2(n_113), .ZN(p_1[16]));
   AOI21_X1 i_34 (.A(n_110), .B1(p_0[17]), .B2(n_111), .ZN(p_1[17]));
   AOI21_X1 i_35 (.A(n_108), .B1(p_0[18]), .B2(n_109), .ZN(p_1[18]));
   AOI21_X1 i_36 (.A(n_106), .B1(p_0[19]), .B2(n_107), .ZN(p_1[19]));
   AOI21_X1 i_37 (.A(n_104), .B1(p_0[20]), .B2(n_105), .ZN(p_1[20]));
   AOI21_X1 i_38 (.A(n_102), .B1(p_0[21]), .B2(n_103), .ZN(p_1[21]));
   AOI21_X1 i_39 (.A(n_100), .B1(p_0[22]), .B2(n_101), .ZN(p_1[22]));
   AOI21_X1 i_40 (.A(n_98), .B1(p_0[23]), .B2(n_99), .ZN(p_1[23]));
   AOI21_X1 i_41 (.A(n_96), .B1(p_0[24]), .B2(n_97), .ZN(p_1[24]));
   AOI21_X1 i_42 (.A(n_94), .B1(p_0[25]), .B2(n_95), .ZN(p_1[25]));
   AOI21_X1 i_43 (.A(n_92), .B1(p_0[26]), .B2(n_93), .ZN(p_1[26]));
   AOI21_X1 i_44 (.A(n_90), .B1(p_0[27]), .B2(n_91), .ZN(p_1[27]));
   AOI21_X1 i_45 (.A(n_88), .B1(p_0[28]), .B2(n_89), .ZN(p_1[28]));
   AOI21_X1 i_46 (.A(n_86), .B1(p_0[29]), .B2(n_87), .ZN(p_1[29]));
   AOI21_X1 i_47 (.A(n_84), .B1(p_0[30]), .B2(n_85), .ZN(p_1[30]));
   AOI21_X1 i_48 (.A(n_82), .B1(p_0[31]), .B2(n_83), .ZN(p_1[31]));
   AOI21_X1 i_49 (.A(n_23), .B1(p_0[32]), .B2(n_81), .ZN(p_1[32]));
   AOI21_X1 i_50 (.A(n_21), .B1(p_0[33]), .B2(n_22), .ZN(p_1[33]));
   AOI21_X1 i_51 (.A(n_19), .B1(p_0[34]), .B2(n_20), .ZN(p_1[34]));
   AOI21_X1 i_52 (.A(n_31), .B1(p_0[35]), .B2(n_18), .ZN(p_1[35]));
   INV_X1 i_53 (.A(n_19), .ZN(n_18));
   NOR2_X1 i_54 (.A1(p_0[34]), .A2(n_20), .ZN(n_19));
   INV_X1 i_55 (.A(n_21), .ZN(n_20));
   NOR2_X1 i_56 (.A1(p_0[33]), .A2(n_22), .ZN(n_21));
   INV_X1 i_57 (.A(n_23), .ZN(n_22));
   NOR2_X1 i_58 (.A1(p_0[32]), .A2(n_81), .ZN(n_23));
   AOI21_X1 i_59 (.A(n_29), .B1(p_0[36]), .B2(n_30), .ZN(p_1[36]));
   AOI21_X1 i_60 (.A(n_27), .B1(p_0[37]), .B2(n_28), .ZN(p_1[37]));
   AOI21_X1 i_61 (.A(n_25), .B1(p_0[38]), .B2(n_26), .ZN(p_1[38]));
   AOI21_X1 i_62 (.A(n_77), .B1(p_0[39]), .B2(n_24), .ZN(p_1[39]));
   INV_X1 i_63 (.A(n_25), .ZN(n_24));
   NOR2_X1 i_64 (.A1(p_0[38]), .A2(n_26), .ZN(n_25));
   INV_X1 i_65 (.A(n_27), .ZN(n_26));
   NOR2_X1 i_66 (.A1(p_0[37]), .A2(n_28), .ZN(n_27));
   INV_X1 i_67 (.A(n_29), .ZN(n_28));
   NOR2_X1 i_68 (.A1(p_0[36]), .A2(n_30), .ZN(n_29));
   INV_X1 i_69 (.A(n_31), .ZN(n_30));
   NOR2_X1 i_70 (.A1(n_81), .A2(n_79), .ZN(n_31));
   AOI21_X1 i_71 (.A(n_37), .B1(p_0[40]), .B2(n_76), .ZN(p_1[40]));
   AOI21_X1 i_72 (.A(n_35), .B1(p_0[41]), .B2(n_36), .ZN(p_1[41]));
   AOI21_X1 i_73 (.A(n_33), .B1(p_0[42]), .B2(n_34), .ZN(p_1[42]));
   AOI21_X1 i_74 (.A(n_75), .B1(p_0[43]), .B2(n_32), .ZN(p_1[43]));
   INV_X1 i_75 (.A(n_33), .ZN(n_32));
   NOR2_X1 i_76 (.A1(n_80), .A2(n_76), .ZN(n_33));
   INV_X1 i_77 (.A(n_35), .ZN(n_34));
   NOR2_X1 i_78 (.A1(p_0[41]), .A2(n_36), .ZN(n_35));
   INV_X1 i_79 (.A(n_37), .ZN(n_36));
   NOR2_X1 i_80 (.A1(p_0[40]), .A2(n_76), .ZN(n_37));
   AOI21_X1 i_81 (.A(n_73), .B1(p_0[44]), .B2(n_74), .ZN(p_1[44]));
   AOI21_X1 i_82 (.A(n_71), .B1(p_0[45]), .B2(n_72), .ZN(p_1[45]));
   AOI21_X1 i_83 (.A(n_69), .B1(p_0[46]), .B2(n_70), .ZN(p_1[46]));
   AOI21_X1 i_84 (.A(n_67), .B1(p_0[47]), .B2(n_68), .ZN(p_1[47]));
   AOI21_X1 i_85 (.A(n_43), .B1(p_0[48]), .B2(n_66), .ZN(p_1[48]));
   AOI21_X1 i_86 (.A(n_41), .B1(p_0[49]), .B2(n_42), .ZN(p_1[49]));
   AOI21_X1 i_95 (.A(n_45), .B1(p_0[52]), .B2(n_49), .ZN(p_1[52]));
   INV_X1 i_96 (.A(n_44), .ZN(p_1[53]));
   OAI21_X1 i_97 (.A(n_46), .B1(n_129), .B2(n_45), .ZN(n_44));
   NOR2_X1 i_98 (.A1(p_0[52]), .A2(n_49), .ZN(n_45));
   AOI21_X1 i_99 (.A(n_48), .B1(p_0[54]), .B2(n_46), .ZN(p_1[54]));
   OR3_X1 i_100 (.A1(p_0[53]), .A2(p_0[52]), .A3(n_49), .ZN(n_46));
   AOI21_X1 i_101 (.A(n_62), .B1(p_0[55]), .B2(n_47), .ZN(p_1[55]));
   INV_X1 i_102 (.A(n_48), .ZN(n_47));
   NOR2_X1 i_103 (.A1(n_63), .A2(n_49), .ZN(n_48));
   AOI21_X1 i_105 (.A(n_51), .B1(p_0[56]), .B2(n_61), .ZN(p_1[56]));
   AOI21_X1 i_109 (.A(n_54), .B1(p_0[58]), .B2(n_52), .ZN(p_1[58]));
   NOR2_X1 i_113 (.A1(n_65), .A2(n_61), .ZN(n_54));
   INV_X1 i_192 (.A(p_0[53]), .ZN(n_129));
   NAND3_X1 i_87 (.A1(n_162), .A2(n_60), .A3(n_161), .ZN(n_65));
   INV_X1 i_88 (.A(n_66), .ZN(n_67));
   INV_X1 i_89 (.A(n_88), .ZN(n_87));
   INV_X1 i_90 (.A(n_91), .ZN(n_92));
   INV_X1 i_91 (.A(n_96), .ZN(n_95));
   INV_X1 i_92 (.A(n_107), .ZN(n_108));
   INV_X1 i_93 (.A(n_112), .ZN(n_111));
   NAND2_X1 i_94 (.A1(n_172), .A2(n_173), .ZN(n_115));
   INV_X1 i_104 (.A(n_113), .ZN(n_114));
   INV_X1 i_106 (.A(n_117), .ZN(n_116));
   NAND2_X1 i_107 (.A1(n_185), .A2(n_58), .ZN(n_121));
   INV_X1 i_108 (.A(n_119), .ZN(n_120));
   INV_X1 i_110 (.A(n_123), .ZN(n_122));
   INV_X1 i_111 (.A(n_39), .ZN(n_38));
   OR3_X1 i_112 (.A1(p_0[50]), .A2(p_0[49]), .A3(p_0[48]), .ZN(n_39));
   INV_X1 i_114 (.A(p_0[51]), .ZN(n_40));
   OR2_X1 i_115 (.A1(n_80), .A2(p_0[43]), .ZN(n_50));
   OR3_X1 i_116 (.A1(p_0[42]), .A2(p_0[41]), .A3(p_0[40]), .ZN(n_80));
   OR3_X1 i_117 (.A1(n_79), .A2(p_0[36]), .A3(p_0[37]), .ZN(n_53));
   OR4_X1 i_118 (.A1(p_0[35]), .A2(p_0[34]), .A3(p_0[33]), .A4(p_0[32]), 
      .ZN(n_79));
   INV_X1 i_119 (.A(n_61), .ZN(n_62));
   INV_X1 i_120 (.A(n_93), .ZN(n_94));
   INV_X1 i_121 (.A(n_109), .ZN(n_110));
   OR2_X1 i_122 (.A1(n_63), .A2(n_64), .ZN(n_55));
   NAND2_X1 i_123 (.A1(n_38), .A2(n_40), .ZN(n_64));
   OR3_X1 i_124 (.A1(p_0[53]), .A2(p_0[54]), .A3(p_0[52]), .ZN(n_63));
   OR2_X1 i_125 (.A1(p_0[13]), .A2(p_0[14]), .ZN(n_56));
   OR2_X1 i_126 (.A1(p_0[10]), .A2(p_0[9]), .ZN(n_57));
   INV_X1 i_127 (.A(n_59), .ZN(n_58));
   NAND2_X1 i_128 (.A1(n_184), .A2(n_183), .ZN(n_59));
   INV_X1 i_129 (.A(p_0[58]), .ZN(n_60));
   NAND2_X1 i_130 (.A1(n_163), .A2(n_141), .ZN(n_52));
   INV_X1 i_131 (.A(n_140), .ZN(n_51));
   INV_X1 i_132 (.A(n_132), .ZN(n_41));
   INV_X1 i_133 (.A(n_42), .ZN(n_43));
   NAND2_X1 i_134 (.A1(n_138), .A2(n_134), .ZN(n_42));
   INV_X1 i_135 (.A(n_72), .ZN(n_73));
   NAND2_X1 i_136 (.A1(n_75), .A2(n_209), .ZN(n_72));
   INV_X1 i_137 (.A(n_81), .ZN(n_82));
   NAND2_X1 i_138 (.A1(n_84), .A2(n_207), .ZN(n_81));
   INV_X1 i_139 (.A(n_78), .ZN(n_88));
   NAND2_X1 i_140 (.A1(n_90), .A2(n_204), .ZN(n_78));
   NAND2_X1 i_141 (.A1(n_96), .A2(n_201), .ZN(n_93));
   INV_X1 i_142 (.A(n_99), .ZN(n_100));
   NAND2_X1 i_143 (.A1(n_102), .A2(n_198), .ZN(n_99));
   INV_X1 i_144 (.A(n_105), .ZN(n_106));
   NAND2_X1 i_145 (.A1(n_150), .A2(n_195), .ZN(n_105));
   INV_X1 i_146 (.A(n_128), .ZN(n_112));
   NAND2_X1 i_147 (.A1(n_151), .A2(n_192), .ZN(n_128));
   NAND2_X1 i_148 (.A1(n_179), .A2(n_178), .ZN(n_118));
   NAND2_X1 i_149 (.A1(n_123), .A2(n_181), .ZN(n_119));
   INV_X1 i_150 (.A(n_124), .ZN(n_125));
   NAND2_X1 i_151 (.A1(n_127), .A2(n_190), .ZN(n_124));
   INV_X1 i_152 (.A(n_126), .ZN(n_127));
   NAND2_X1 i_153 (.A1(n_189), .A2(n_188), .ZN(n_126));
   INV_X1 i_154 (.A(n_130), .ZN(p_1[50]));
   NAND2_X1 i_155 (.A1(n_131), .A2(n_133), .ZN(n_130));
   NAND2_X1 i_156 (.A1(n_132), .A2(p_0[50]), .ZN(n_131));
   NAND3_X1 i_157 (.A1(n_138), .A2(n_135), .A3(n_134), .ZN(n_132));
   AOI21_X1 i_158 (.A(n_137), .B1(n_133), .B2(p_0[51]), .ZN(p_1[51]));
   NAND4_X1 i_159 (.A1(n_138), .A2(n_136), .A3(n_135), .A4(n_134), .ZN(n_133));
   INV_X1 i_160 (.A(p_0[48]), .ZN(n_134));
   INV_X1 i_161 (.A(p_0[49]), .ZN(n_135));
   INV_X1 i_162 (.A(p_0[50]), .ZN(n_136));
   INV_X1 i_163 (.A(n_49), .ZN(n_137));
   NAND2_X1 i_164 (.A1(n_138), .A2(n_139), .ZN(n_49));
   INV_X1 i_165 (.A(n_66), .ZN(n_138));
   NAND2_X1 i_166 (.A1(n_69), .A2(n_212), .ZN(n_66));
   INV_X1 i_167 (.A(n_64), .ZN(n_139));
   AOI22_X1 i_168 (.A1(n_140), .A2(p_0[57]), .B1(n_163), .B2(n_141), .ZN(p_1[57]));
   NAND2_X1 i_169 (.A1(n_163), .A2(n_161), .ZN(n_140));
   INV_X1 i_170 (.A(n_160), .ZN(n_141));
   AOI21_X1 i_171 (.A(n_147), .B1(p_0[59]), .B2(n_142), .ZN(p_1[59]));
   INV_X1 i_172 (.A(n_54), .ZN(n_142));
   INV_X1 i_173 (.A(n_143), .ZN(p_1[60]));
   NAND2_X1 i_174 (.A1(n_145), .A2(n_144), .ZN(n_143));
   NAND2_X1 i_175 (.A1(n_148), .A2(p_0[60]), .ZN(n_144));
   NAND2_X1 i_176 (.A1(n_147), .A2(n_213), .ZN(n_145));
   NOR2_X1 i_177 (.A1(n_146), .A2(n_152), .ZN(p_1[61]));
   AOI21_X1 i_178 (.A(n_154), .B1(n_147), .B2(n_213), .ZN(n_146));
   INV_X1 i_179 (.A(n_148), .ZN(n_147));
   NAND4_X1 i_180 (.A1(n_69), .A2(n_212), .A3(n_164), .A4(n_158), .ZN(n_148));
   INV_X1 i_181 (.A(n_68), .ZN(n_69));
   NAND4_X1 i_182 (.A1(n_75), .A2(n_211), .A3(n_210), .A4(n_209), .ZN(n_68));
   INV_X1 i_183 (.A(n_74), .ZN(n_75));
   NAND4_X1 i_184 (.A1(n_84), .A2(n_207), .A3(n_208), .A4(n_166), .ZN(n_74));
   INV_X1 i_185 (.A(n_83), .ZN(n_84));
   NAND4_X1 i_186 (.A1(n_90), .A2(n_206), .A3(n_205), .A4(n_204), .ZN(n_83));
   INV_X1 i_187 (.A(n_89), .ZN(n_90));
   NAND4_X1 i_188 (.A1(n_96), .A2(n_203), .A3(n_202), .A4(n_201), .ZN(n_89));
   INV_X1 i_189 (.A(n_149), .ZN(n_96));
   NAND4_X1 i_190 (.A1(n_102), .A2(n_200), .A3(n_199), .A4(n_198), .ZN(n_149));
   INV_X1 i_191 (.A(n_101), .ZN(n_102));
   NAND4_X1 i_193 (.A1(n_150), .A2(n_197), .A3(n_196), .A4(n_195), .ZN(n_101));
   INV_X1 i_194 (.A(n_107), .ZN(n_150));
   NAND4_X1 i_195 (.A1(n_151), .A2(n_194), .A3(n_193), .A4(n_192), .ZN(n_107));
   INV_X1 i_196 (.A(n_113), .ZN(n_151));
   NAND4_X1 i_197 (.A1(n_123), .A2(n_181), .A3(n_176), .A4(n_170), .ZN(n_113));
   INV_X1 i_198 (.A(n_153), .ZN(n_152));
   AOI21_X1 i_199 (.A(n_155), .B1(n_153), .B2(p_0[62]), .ZN(p_1[62]));
   NAND4_X1 i_200 (.A1(n_163), .A2(n_154), .A3(n_213), .A4(n_158), .ZN(n_153));
   INV_X1 i_201 (.A(p_0[61]), .ZN(n_154));
   INV_X1 i_202 (.A(p_1[63]), .ZN(n_155));
   NAND4_X1 i_203 (.A1(n_163), .A2(n_213), .A3(n_158), .A4(n_156), .ZN(p_1[63]));
   INV_X1 i_204 (.A(n_157), .ZN(n_156));
   OR2_X1 i_205 (.A1(p_0[62]), .A2(p_0[61]), .ZN(n_157));
   INV_X1 i_206 (.A(n_159), .ZN(n_158));
   OR3_X1 i_207 (.A1(n_160), .A2(p_0[59]), .A3(p_0[58]), .ZN(n_159));
   NAND2_X1 i_208 (.A1(n_162), .A2(n_161), .ZN(n_160));
   INV_X1 i_209 (.A(p_0[56]), .ZN(n_161));
   INV_X1 i_210 (.A(p_0[57]), .ZN(n_162));
   INV_X1 i_211 (.A(n_61), .ZN(n_163));
   NAND4_X1 i_212 (.A1(n_71), .A2(n_212), .A3(n_211), .A4(n_164), .ZN(n_61));
   INV_X1 i_213 (.A(n_165), .ZN(n_164));
   OR2_X1 i_214 (.A1(p_0[55]), .A2(n_55), .ZN(n_165));
   INV_X1 i_215 (.A(n_70), .ZN(n_71));
   NAND4_X1 i_216 (.A1(n_77), .A2(n_210), .A3(n_209), .A4(n_208), .ZN(n_70));
   INV_X1 i_217 (.A(n_76), .ZN(n_77));
   NAND4_X1 i_218 (.A1(n_86), .A2(n_207), .A3(n_206), .A4(n_166), .ZN(n_76));
   INV_X1 i_219 (.A(n_167), .ZN(n_166));
   OR3_X1 i_220 (.A1(p_0[39]), .A2(p_0[38]), .A3(n_53), .ZN(n_167));
   INV_X1 i_221 (.A(n_85), .ZN(n_86));
   NAND4_X1 i_222 (.A1(n_168), .A2(n_205), .A3(n_204), .A4(n_203), .ZN(n_85));
   INV_X1 i_223 (.A(n_91), .ZN(n_168));
   NAND4_X1 i_224 (.A1(n_98), .A2(n_202), .A3(n_201), .A4(n_200), .ZN(n_91));
   INV_X1 i_225 (.A(n_97), .ZN(n_98));
   NAND4_X1 i_226 (.A1(n_104), .A2(n_199), .A3(n_198), .A4(n_197), .ZN(n_97));
   INV_X1 i_227 (.A(n_103), .ZN(n_104));
   NAND4_X1 i_228 (.A1(n_169), .A2(n_196), .A3(n_195), .A4(n_194), .ZN(n_103));
   INV_X1 i_229 (.A(n_109), .ZN(n_169));
   NAND4_X1 i_230 (.A1(n_117), .A2(n_193), .A3(n_192), .A4(n_170), .ZN(n_109));
   INV_X1 i_231 (.A(n_171), .ZN(n_170));
   NAND3_X1 i_232 (.A1(n_174), .A2(n_173), .A3(n_172), .ZN(n_171));
   INV_X1 i_233 (.A(n_56), .ZN(n_172));
   INV_X1 i_234 (.A(p_0[12]), .ZN(n_173));
   INV_X1 i_235 (.A(p_0[15]), .ZN(n_174));
   INV_X1 i_236 (.A(n_175), .ZN(n_117));
   NAND3_X1 i_237 (.A1(n_123), .A2(n_181), .A3(n_176), .ZN(n_175));
   INV_X1 i_238 (.A(n_177), .ZN(n_176));
   NAND3_X1 i_239 (.A1(n_180), .A2(n_179), .A3(n_178), .ZN(n_177));
   INV_X1 i_240 (.A(n_57), .ZN(n_178));
   INV_X1 i_241 (.A(p_0[8]), .ZN(n_179));
   INV_X1 i_242 (.A(p_0[11]), .ZN(n_180));
   INV_X1 i_243 (.A(n_182), .ZN(n_181));
   NAND4_X1 i_244 (.A1(n_186), .A2(n_185), .A3(n_184), .A4(n_183), .ZN(n_182));
   INV_X1 i_245 (.A(p_0[4]), .ZN(n_183));
   INV_X1 i_246 (.A(p_0[5]), .ZN(n_184));
   INV_X1 i_247 (.A(p_0[6]), .ZN(n_185));
   INV_X1 i_248 (.A(p_0[7]), .ZN(n_186));
   INV_X1 i_249 (.A(n_187), .ZN(n_123));
   NAND4_X1 i_250 (.A1(n_191), .A2(n_190), .A3(n_189), .A4(n_188), .ZN(n_187));
   INV_X1 i_251 (.A(p_0[0]), .ZN(n_188));
   INV_X1 i_252 (.A(p_0[1]), .ZN(n_189));
   INV_X1 i_253 (.A(p_0[2]), .ZN(n_190));
   INV_X1 i_254 (.A(p_0[3]), .ZN(n_191));
   INV_X1 i_255 (.A(p_0[16]), .ZN(n_192));
   INV_X1 i_256 (.A(p_0[17]), .ZN(n_193));
   INV_X1 i_257 (.A(p_0[18]), .ZN(n_194));
   INV_X1 i_258 (.A(p_0[19]), .ZN(n_195));
   INV_X1 i_259 (.A(p_0[20]), .ZN(n_196));
   INV_X1 i_260 (.A(p_0[21]), .ZN(n_197));
   INV_X1 i_261 (.A(p_0[22]), .ZN(n_198));
   INV_X1 i_262 (.A(p_0[23]), .ZN(n_199));
   INV_X1 i_263 (.A(p_0[24]), .ZN(n_200));
   INV_X1 i_264 (.A(p_0[25]), .ZN(n_201));
   INV_X1 i_265 (.A(p_0[26]), .ZN(n_202));
   INV_X1 i_266 (.A(p_0[27]), .ZN(n_203));
   INV_X1 i_267 (.A(p_0[28]), .ZN(n_204));
   INV_X1 i_268 (.A(p_0[29]), .ZN(n_205));
   INV_X1 i_269 (.A(p_0[30]), .ZN(n_206));
   INV_X1 i_270 (.A(p_0[31]), .ZN(n_207));
   INV_X1 i_271 (.A(n_50), .ZN(n_208));
   INV_X1 i_272 (.A(p_0[44]), .ZN(n_209));
   INV_X1 i_273 (.A(p_0[45]), .ZN(n_210));
   INV_X1 i_274 (.A(p_0[46]), .ZN(n_211));
   INV_X1 i_275 (.A(p_0[47]), .ZN(n_212));
   INV_X1 i_276 (.A(p_0[60]), .ZN(n_213));
endmodule

module seq_multiplier(clk, rst, a, b, c);
   input clk;
   input rst;
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_0_5;
   wire n_0_0_0;
   wire n_0_0_6;
   wire n_0_0_1;
   wire n_0_0_7;
   wire n_0_0_2;
   wire n_0_0_8;
   wire n_0_0_3;
   wire n_0_0_9;
   wire n_0_0_4;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_0_10;
   wire n_0_166;
   wire n_0_0_11;
   wire n_0_167;
   wire n_0_0_12;
   wire n_0_168;
   wire n_0_0_13;
   wire n_0_169;
   wire n_0_0_14;
   wire n_0_170;
   wire n_0_0_15;
   wire n_0_171;
   wire n_0_0_16;
   wire n_0_172;
   wire n_0_0_17;
   wire n_0_173;
   wire n_0_0_18;
   wire n_0_174;
   wire n_0_0_19;
   wire n_0_175;
   wire n_0_0_20;
   wire n_0_176;
   wire n_0_0_21;
   wire n_0_177;
   wire n_0_0_22;
   wire n_0_178;
   wire n_0_0_23;
   wire n_0_179;
   wire n_0_0_24;
   wire n_0_180;
   wire n_0_0_25;
   wire n_0_181;
   wire n_0_0_26;
   wire n_0_182;
   wire n_0_0_27;
   wire n_0_183;
   wire n_0_0_28;
   wire n_0_184;
   wire n_0_0_29;
   wire n_0_185;
   wire n_0_0_30;
   wire n_0_186;
   wire n_0_0_31;
   wire n_0_187;
   wire n_0_0_32;
   wire n_0_188;
   wire n_0_0_33;
   wire n_0_189;
   wire n_0_0_34;
   wire n_0_190;
   wire n_0_0_35;
   wire n_0_191;
   wire n_0_0_36;
   wire n_0_192;
   wire n_0_0_37;
   wire n_0_193;
   wire n_0_0_38;
   wire n_0_194;
   wire n_0_0_39;
   wire n_0_195;
   wire n_0_0_40;
   wire n_0_196;
   wire n_0_0_41;
   wire n_0_197;
   wire n_0_0_42;
   wire n_0_198;
   wire n_0_0_43;
   wire n_0_199;
   wire n_0_0_44;
   wire n_0_200;
   wire n_0_0_45;
   wire n_0_201;
   wire n_0_0_46;
   wire n_0_202;
   wire n_0_0_47;
   wire n_0_203;
   wire n_0_0_48;
   wire n_0_204;
   wire n_0_0_49;
   wire n_0_205;
   wire n_0_0_50;
   wire n_0_206;
   wire n_0_0_51;
   wire n_0_207;
   wire n_0_0_52;
   wire n_0_208;
   wire n_0_0_53;
   wire n_0_209;
   wire n_0_0_54;
   wire n_0_210;
   wire n_0_0_55;
   wire n_0_211;
   wire n_0_0_56;
   wire n_0_212;
   wire n_0_0_57;
   wire n_0_213;
   wire n_0_0_58;
   wire n_0_214;
   wire n_0_0_59;
   wire n_0_215;
   wire n_0_0_60;
   wire n_0_216;
   wire n_0_0_61;
   wire n_0_217;
   wire n_0_0_62;
   wire n_0_218;
   wire n_0_0_63;
   wire n_0_219;
   wire n_0_0_64;
   wire n_0_220;
   wire n_0_0_65;
   wire n_0_221;
   wire n_0_0_66;
   wire n_0_222;
   wire n_0_0_67;
   wire n_0_223;
   wire n_0_0_68;
   wire n_0_224;
   wire n_0_0_69;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_0_75;
   wire n_0_355;
   wire n_0_0_76;
   wire n_0_357;
   wire n_0_0_78;
   wire n_0_358;
   wire n_0_0_79;
   wire n_0_359;
   wire n_0_0_80;
   wire n_0_360;
   wire n_0_0_81;
   wire n_0_367;
   wire n_0_0_88;
   wire n_0_368;
   wire n_0_0_89;
   wire n_0_369;
   wire n_0_0_90;
   wire n_0_370;
   wire n_0_0_91;
   wire n_0_371;
   wire n_0_0_92;
   wire n_0_372;
   wire n_0_0_93;
   wire n_0_373;
   wire n_0_0_94;
   wire n_0_374;
   wire n_0_0_95;
   wire n_0_375;
   wire n_0_0_96;
   wire n_0_376;
   wire n_0_0_97;
   wire n_0_377;
   wire n_0_0_98;
   wire n_0_378;
   wire n_0_0_99;
   wire n_0_379;
   wire n_0_0_100;
   wire n_0_380;
   wire n_0_0_101;
   wire n_0_381;
   wire n_0_0_102;
   wire n_0_382;
   wire n_0_0_103;
   wire n_0_383;
   wire n_0_0_104;
   wire n_0_384;
   wire n_0_0_105;
   wire n_0_385;
   wire n_0_0_107;
   wire n_0_386;
   wire n_0_0_109;
   wire n_0_387;
   wire n_0_0_110;
   wire n_0_388;
   wire n_0_0_111;
   wire n_0_389;
   wire n_0_0_112;
   wire n_0_390;
   wire n_0_0_113;
   wire n_0_391;
   wire n_0_0_114;
   wire n_0_392;
   wire n_0_0_115;
   wire n_0_393;
   wire n_0_0_116;
   wire n_0_394;
   wire n_0_0_117;
   wire n_0_395;
   wire n_0_0_118;
   wire n_0_396;
   wire n_0_0_119;
   wire n_0_397;
   wire n_0_0_120;
   wire n_0_398;
   wire n_0_0_121;
   wire n_0_399;
   wire n_0_0_122;
   wire n_0_400;
   wire n_0_0_123;
   wire n_0_401;
   wire n_0_0_124;
   wire n_0_402;
   wire n_0_0_125;
   wire n_0_403;
   wire n_0_0_126;
   wire n_0_404;
   wire n_0_0_127;
   wire n_0_405;
   wire n_0_0_128;
   wire n_0_406;
   wire n_0_0_129;
   wire n_0_407;
   wire n_0_0_130;
   wire n_0_408;
   wire n_0_0_131;
   wire n_0_409;
   wire n_0_0_132;
   wire n_0_410;
   wire n_0_0_133;
   wire n_0_411;
   wire n_0_0_134;
   wire n_0_412;
   wire n_0_0_135;
   wire n_0_413;
   wire n_0_0_136;
   wire n_0_414;
   wire n_0_0_137;
   wire n_0_415;
   wire n_0_0_138;
   wire n_0_416;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_417;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_418;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_226;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_361;
   wire n_0_0_82;
   wire n_0_0_72;
   wire n_0_0_158;
   wire n_0_362;
   wire n_0_0_83;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_363;
   wire n_0_0_84;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_364;
   wire n_0_0_85;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_365;
   wire n_0_0_86;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_366;
   wire n_0_0_87;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_157;
   wire n_0_225;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_227;
   wire n_0_0_171;
   wire n_0_0_73;
   wire n_0_0_172;
   wire n_0_0_74;
   wire n_0_356;
   wire n_0_0_77;
   wire n_0_0_173;
   wire n_0_0_106;
   wire n_0_0_174;
   wire n_0_0_108;
   wire n_0_0_144;
   wire [6:0]counter;
   wire [31:0]A_r;
   wire [31:0]B_r;
   wire [31:0]Accumulator;
   wire negative;

   CLKGATETST_X1 clk_gate_c_reg (.CK(clk), .E(n_0_418), .SE(1'b0), .GCK(n_0_0));
   DFF_X1 \c_reg[63]  (.D(n_0_228), .CK(n_0_0), .Q(c[63]), .QN());
   DFF_X1 \c_reg[62]  (.D(n_0_227), .CK(n_0_0), .Q(c[62]), .QN());
   DFF_X1 \c_reg[61]  (.D(n_0_226), .CK(n_0_0), .Q(c[61]), .QN());
   DFF_X1 \c_reg[60]  (.D(n_0_225), .CK(n_0_0), .Q(c[60]), .QN());
   DFF_X1 \c_reg[59]  (.D(n_0_224), .CK(n_0_0), .Q(c[59]), .QN());
   DFF_X1 \c_reg[58]  (.D(n_0_223), .CK(n_0_0), .Q(c[58]), .QN());
   DFF_X1 \c_reg[57]  (.D(n_0_222), .CK(n_0_0), .Q(c[57]), .QN());
   DFF_X1 \c_reg[56]  (.D(n_0_221), .CK(n_0_0), .Q(c[56]), .QN());
   DFF_X1 \c_reg[55]  (.D(n_0_220), .CK(n_0_0), .Q(c[55]), .QN());
   DFF_X1 \c_reg[54]  (.D(n_0_219), .CK(n_0_0), .Q(c[54]), .QN());
   DFF_X1 \c_reg[53]  (.D(n_0_218), .CK(n_0_0), .Q(c[53]), .QN());
   DFF_X1 \c_reg[52]  (.D(n_0_217), .CK(n_0_0), .Q(c[52]), .QN());
   DFF_X1 \c_reg[51]  (.D(n_0_216), .CK(n_0_0), .Q(c[51]), .QN());
   DFF_X1 \c_reg[50]  (.D(n_0_215), .CK(n_0_0), .Q(c[50]), .QN());
   DFF_X1 \c_reg[49]  (.D(n_0_214), .CK(n_0_0), .Q(c[49]), .QN());
   DFF_X1 \c_reg[48]  (.D(n_0_213), .CK(n_0_0), .Q(c[48]), .QN());
   DFF_X1 \c_reg[47]  (.D(n_0_212), .CK(n_0_0), .Q(c[47]), .QN());
   DFF_X1 \c_reg[46]  (.D(n_0_211), .CK(n_0_0), .Q(c[46]), .QN());
   DFF_X1 \c_reg[45]  (.D(n_0_210), .CK(n_0_0), .Q(c[45]), .QN());
   DFF_X1 \c_reg[44]  (.D(n_0_209), .CK(n_0_0), .Q(c[44]), .QN());
   DFF_X1 \c_reg[43]  (.D(n_0_208), .CK(n_0_0), .Q(c[43]), .QN());
   DFF_X1 \c_reg[42]  (.D(n_0_207), .CK(n_0_0), .Q(c[42]), .QN());
   DFF_X1 \c_reg[41]  (.D(n_0_206), .CK(n_0_0), .Q(c[41]), .QN());
   DFF_X1 \c_reg[40]  (.D(n_0_205), .CK(n_0_0), .Q(c[40]), .QN());
   DFF_X1 \c_reg[39]  (.D(n_0_204), .CK(n_0_0), .Q(c[39]), .QN());
   DFF_X1 \c_reg[38]  (.D(n_0_203), .CK(n_0_0), .Q(c[38]), .QN());
   DFF_X1 \c_reg[37]  (.D(n_0_202), .CK(n_0_0), .Q(c[37]), .QN());
   DFF_X1 \c_reg[36]  (.D(n_0_201), .CK(n_0_0), .Q(c[36]), .QN());
   DFF_X1 \c_reg[35]  (.D(n_0_200), .CK(n_0_0), .Q(c[35]), .QN());
   DFF_X1 \c_reg[34]  (.D(n_0_199), .CK(n_0_0), .Q(c[34]), .QN());
   DFF_X1 \c_reg[33]  (.D(n_0_198), .CK(n_0_0), .Q(c[33]), .QN());
   DFF_X1 \c_reg[32]  (.D(n_0_197), .CK(n_0_0), .Q(c[32]), .QN());
   DFF_X1 \c_reg[31]  (.D(n_0_196), .CK(n_0_0), .Q(c[31]), .QN());
   DFF_X1 \c_reg[30]  (.D(n_0_195), .CK(n_0_0), .Q(c[30]), .QN());
   DFF_X1 \c_reg[29]  (.D(n_0_194), .CK(n_0_0), .Q(c[29]), .QN());
   DFF_X1 \c_reg[28]  (.D(n_0_193), .CK(n_0_0), .Q(c[28]), .QN());
   DFF_X1 \c_reg[27]  (.D(n_0_192), .CK(n_0_0), .Q(c[27]), .QN());
   DFF_X1 \c_reg[26]  (.D(n_0_191), .CK(n_0_0), .Q(c[26]), .QN());
   DFF_X1 \c_reg[25]  (.D(n_0_190), .CK(n_0_0), .Q(c[25]), .QN());
   DFF_X1 \c_reg[24]  (.D(n_0_189), .CK(n_0_0), .Q(c[24]), .QN());
   DFF_X1 \c_reg[23]  (.D(n_0_188), .CK(n_0_0), .Q(c[23]), .QN());
   DFF_X1 \c_reg[22]  (.D(n_0_187), .CK(n_0_0), .Q(c[22]), .QN());
   DFF_X1 \c_reg[21]  (.D(n_0_186), .CK(n_0_0), .Q(c[21]), .QN());
   DFF_X1 \c_reg[20]  (.D(n_0_185), .CK(n_0_0), .Q(c[20]), .QN());
   DFF_X1 \c_reg[19]  (.D(n_0_184), .CK(n_0_0), .Q(c[19]), .QN());
   DFF_X1 \c_reg[18]  (.D(n_0_183), .CK(n_0_0), .Q(c[18]), .QN());
   DFF_X1 \c_reg[17]  (.D(n_0_182), .CK(n_0_0), .Q(c[17]), .QN());
   DFF_X1 \c_reg[16]  (.D(n_0_181), .CK(n_0_0), .Q(c[16]), .QN());
   DFF_X1 \c_reg[15]  (.D(n_0_180), .CK(n_0_0), .Q(c[15]), .QN());
   DFF_X1 \c_reg[14]  (.D(n_0_179), .CK(n_0_0), .Q(c[14]), .QN());
   DFF_X1 \c_reg[13]  (.D(n_0_178), .CK(n_0_0), .Q(c[13]), .QN());
   DFF_X1 \c_reg[12]  (.D(n_0_177), .CK(n_0_0), .Q(c[12]), .QN());
   DFF_X1 \c_reg[11]  (.D(n_0_176), .CK(n_0_0), .Q(c[11]), .QN());
   DFF_X1 \c_reg[10]  (.D(n_0_175), .CK(n_0_0), .Q(c[10]), .QN());
   DFF_X1 \c_reg[9]  (.D(n_0_174), .CK(n_0_0), .Q(c[9]), .QN());
   DFF_X1 \c_reg[8]  (.D(n_0_173), .CK(n_0_0), .Q(c[8]), .QN());
   DFF_X1 \c_reg[7]  (.D(n_0_172), .CK(n_0_0), .Q(c[7]), .QN());
   DFF_X1 \c_reg[6]  (.D(n_0_171), .CK(n_0_0), .Q(c[6]), .QN());
   DFF_X1 \c_reg[5]  (.D(n_0_170), .CK(n_0_0), .Q(c[5]), .QN());
   DFF_X1 \c_reg[4]  (.D(n_0_169), .CK(n_0_0), .Q(c[4]), .QN());
   DFF_X1 \c_reg[3]  (.D(n_0_168), .CK(n_0_0), .Q(c[3]), .QN());
   DFF_X1 \c_reg[2]  (.D(n_0_167), .CK(n_0_0), .Q(c[2]), .QN());
   DFF_X1 \c_reg[1]  (.D(n_0_166), .CK(n_0_0), .Q(c[1]), .QN());
   DFF_X1 \c_reg[0]  (.D(n_0_260), .CK(n_0_0), .Q(c[0]), .QN());
   datapath i_0_1 (.a(a), .p_0({n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
      n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, 
      n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, 
      n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, uc_0}));
   datapath__0_2 i_0_4 (.b(b), .p_0({n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, 
      n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, 
      n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, 
      n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, uc_1}));
   datapath__0_6 i_0_8 (.p_0({n_0_354, n_0_353, n_0_352, n_0_351, n_0_350, 
      n_0_349, n_0_348, n_0_347, n_0_346, n_0_345, n_0_344, n_0_343, n_0_342, 
      n_0_341, n_0_340, n_0_339, n_0_338, n_0_337, n_0_336, n_0_335, n_0_334, 
      n_0_333, n_0_332, n_0_331, n_0_330, n_0_329, n_0_328, n_0_327, n_0_326, 
      n_0_325, n_0_324, n_0_323}), .Accumulator({uc_2, n_0_322, n_0_321, n_0_320, 
      n_0_319, n_0_318, n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, n_0_312, 
      n_0_311, n_0_310, n_0_309, n_0_308, n_0_307, n_0_306, n_0_305, n_0_304, 
      n_0_303, n_0_302, n_0_301, n_0_300, n_0_299, n_0_298, n_0_297, n_0_296, 
      n_0_295, n_0_294, n_0_293, n_0_292}), .Accumulator1({n_0_94, n_0_93, 
      n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, 
      n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, 
      n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, 
      n_0_65, n_0_64, n_0_63}));
   datapath__0_9 i_0_11 (.p_0({uc_3, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, 
      n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, 
      n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, 
      n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, 
      n_0_385, n_0_384, n_0_383, n_0_382, n_0_381, n_0_380, n_0_379, n_0_378, 
      n_0_377, n_0_376, n_0_375, n_0_374, n_0_373, n_0_372, n_0_371, n_0_370, 
      n_0_369, n_0_368, n_0_367, n_0_366, n_0_365, n_0_364, n_0_363, n_0_362, 
      n_0_361, n_0_360, n_0_359, n_0_358, n_0_357, n_0_356, n_0_355}), .p_1({
      n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, 
      n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, 
      n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, 
      n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, 
      n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, 
      n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, 
      n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, 
      n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, uc_4}));
   HA_X1 i_0_0_0 (.A(counter[1]), .B(counter[0]), .CO(n_0_0_0), .S(n_0_0_5));
   HA_X1 i_0_0_1 (.A(counter[2]), .B(n_0_0_0), .CO(n_0_0_1), .S(n_0_0_6));
   HA_X1 i_0_0_2 (.A(counter[3]), .B(n_0_0_1), .CO(n_0_0_2), .S(n_0_0_7));
   HA_X1 i_0_0_3 (.A(counter[4]), .B(n_0_0_2), .CO(n_0_0_3), .S(n_0_0_8));
   HA_X1 i_0_0_4 (.A(counter[5]), .B(n_0_0_3), .CO(n_0_0_4), .S(n_0_0_9));
   NOR2_X1 i_0_0_5 (.A1(rst), .A2(counter[0]), .ZN(n_0_158));
   AND2_X1 i_0_0_6 (.A1(n_0_0_5), .A2(n_0_0_147), .ZN(n_0_159));
   AND2_X1 i_0_0_7 (.A1(n_0_0_6), .A2(n_0_0_147), .ZN(n_0_160));
   AND2_X1 i_0_0_8 (.A1(n_0_0_7), .A2(n_0_0_147), .ZN(n_0_161));
   AND2_X1 i_0_0_9 (.A1(n_0_0_8), .A2(n_0_0_147), .ZN(n_0_162));
   AND2_X1 i_0_0_10 (.A1(n_0_0_9), .A2(n_0_0_147), .ZN(n_0_163));
   AOI221_X1 i_0_0_11 (.A(n_0_418), .B1(n_0_0_156), .B2(n_0_0_152), .C1(
      counter[6]), .C2(n_0_0_4), .ZN(n_0_164));
   AOI211_X1 i_0_0_12 (.A(n_0_0_10), .B(rst), .C1(n_0_0_153), .C2(n_0_0_144), 
      .ZN(n_0_165));
   AOI221_X1 i_0_0_13 (.A(n_0_0_144), .B1(a[31]), .B2(n_0_0_154), .C1(n_0_0_155), 
      .C2(b[31]), .ZN(n_0_0_10));
   INV_X1 i_0_0_14 (.A(n_0_0_11), .ZN(n_0_166));
   AOI22_X1 i_0_0_15 (.A1(n_0_356), .A2(n_0_0_73), .B1(n_0_95), .B2(n_0_0_74), 
      .ZN(n_0_0_11));
   INV_X1 i_0_0_16 (.A(n_0_0_12), .ZN(n_0_167));
   AOI22_X1 i_0_0_17 (.A1(n_0_357), .A2(n_0_0_73), .B1(n_0_96), .B2(n_0_0_74), 
      .ZN(n_0_0_12));
   INV_X1 i_0_0_18 (.A(n_0_0_13), .ZN(n_0_168));
   AOI22_X1 i_0_0_19 (.A1(n_0_358), .A2(n_0_0_73), .B1(n_0_97), .B2(n_0_0_74), 
      .ZN(n_0_0_13));
   INV_X1 i_0_0_20 (.A(n_0_0_14), .ZN(n_0_169));
   AOI22_X1 i_0_0_21 (.A1(n_0_359), .A2(n_0_0_73), .B1(n_0_98), .B2(n_0_0_74), 
      .ZN(n_0_0_14));
   INV_X1 i_0_0_22 (.A(n_0_0_15), .ZN(n_0_170));
   AOI22_X1 i_0_0_23 (.A1(n_0_360), .A2(n_0_0_73), .B1(n_0_99), .B2(n_0_0_74), 
      .ZN(n_0_0_15));
   INV_X1 i_0_0_24 (.A(n_0_0_16), .ZN(n_0_171));
   AOI22_X1 i_0_0_25 (.A1(n_0_361), .A2(n_0_0_73), .B1(n_0_100), .B2(n_0_0_74), 
      .ZN(n_0_0_16));
   INV_X1 i_0_0_26 (.A(n_0_0_17), .ZN(n_0_172));
   AOI22_X1 i_0_0_27 (.A1(n_0_362), .A2(n_0_0_73), .B1(n_0_101), .B2(n_0_0_74), 
      .ZN(n_0_0_17));
   INV_X1 i_0_0_28 (.A(n_0_0_18), .ZN(n_0_173));
   AOI22_X1 i_0_0_29 (.A1(n_0_363), .A2(n_0_0_73), .B1(n_0_102), .B2(n_0_0_74), 
      .ZN(n_0_0_18));
   INV_X1 i_0_0_30 (.A(n_0_0_19), .ZN(n_0_174));
   AOI22_X1 i_0_0_31 (.A1(n_0_364), .A2(n_0_0_73), .B1(n_0_103), .B2(n_0_0_74), 
      .ZN(n_0_0_19));
   INV_X1 i_0_0_32 (.A(n_0_0_20), .ZN(n_0_175));
   AOI22_X1 i_0_0_33 (.A1(n_0_365), .A2(n_0_0_73), .B1(n_0_104), .B2(n_0_0_74), 
      .ZN(n_0_0_20));
   INV_X1 i_0_0_34 (.A(n_0_0_21), .ZN(n_0_176));
   AOI22_X1 i_0_0_35 (.A1(n_0_366), .A2(n_0_0_73), .B1(n_0_105), .B2(n_0_0_74), 
      .ZN(n_0_0_21));
   INV_X1 i_0_0_36 (.A(n_0_0_22), .ZN(n_0_177));
   AOI22_X1 i_0_0_37 (.A1(n_0_367), .A2(n_0_0_73), .B1(n_0_106), .B2(n_0_0_74), 
      .ZN(n_0_0_22));
   INV_X1 i_0_0_38 (.A(n_0_0_23), .ZN(n_0_178));
   AOI22_X1 i_0_0_39 (.A1(n_0_368), .A2(n_0_0_73), .B1(n_0_107), .B2(n_0_0_74), 
      .ZN(n_0_0_23));
   INV_X1 i_0_0_40 (.A(n_0_0_24), .ZN(n_0_179));
   AOI22_X1 i_0_0_41 (.A1(n_0_369), .A2(n_0_0_73), .B1(n_0_108), .B2(n_0_0_74), 
      .ZN(n_0_0_24));
   INV_X1 i_0_0_42 (.A(n_0_0_25), .ZN(n_0_180));
   AOI22_X1 i_0_0_43 (.A1(n_0_370), .A2(n_0_0_73), .B1(n_0_109), .B2(n_0_0_74), 
      .ZN(n_0_0_25));
   INV_X1 i_0_0_44 (.A(n_0_0_26), .ZN(n_0_181));
   AOI22_X1 i_0_0_45 (.A1(n_0_371), .A2(n_0_0_73), .B1(n_0_110), .B2(n_0_0_74), 
      .ZN(n_0_0_26));
   INV_X1 i_0_0_46 (.A(n_0_0_27), .ZN(n_0_182));
   AOI22_X1 i_0_0_47 (.A1(n_0_372), .A2(n_0_0_73), .B1(n_0_111), .B2(n_0_0_74), 
      .ZN(n_0_0_27));
   INV_X1 i_0_0_48 (.A(n_0_0_28), .ZN(n_0_183));
   AOI22_X1 i_0_0_49 (.A1(n_0_373), .A2(n_0_0_73), .B1(n_0_112), .B2(n_0_0_74), 
      .ZN(n_0_0_28));
   INV_X1 i_0_0_50 (.A(n_0_0_29), .ZN(n_0_184));
   AOI22_X1 i_0_0_51 (.A1(n_0_374), .A2(n_0_0_73), .B1(n_0_113), .B2(n_0_0_74), 
      .ZN(n_0_0_29));
   INV_X1 i_0_0_52 (.A(n_0_0_30), .ZN(n_0_185));
   AOI22_X1 i_0_0_53 (.A1(n_0_375), .A2(n_0_0_73), .B1(n_0_114), .B2(n_0_0_74), 
      .ZN(n_0_0_30));
   INV_X1 i_0_0_54 (.A(n_0_0_31), .ZN(n_0_186));
   AOI22_X1 i_0_0_55 (.A1(n_0_376), .A2(n_0_0_73), .B1(n_0_115), .B2(n_0_0_74), 
      .ZN(n_0_0_31));
   INV_X1 i_0_0_56 (.A(n_0_0_32), .ZN(n_0_187));
   AOI22_X1 i_0_0_57 (.A1(n_0_377), .A2(n_0_0_73), .B1(n_0_116), .B2(n_0_0_74), 
      .ZN(n_0_0_32));
   INV_X1 i_0_0_58 (.A(n_0_0_33), .ZN(n_0_188));
   AOI22_X1 i_0_0_59 (.A1(n_0_378), .A2(n_0_0_73), .B1(n_0_117), .B2(n_0_0_74), 
      .ZN(n_0_0_33));
   INV_X1 i_0_0_60 (.A(n_0_0_34), .ZN(n_0_189));
   AOI22_X1 i_0_0_61 (.A1(n_0_379), .A2(n_0_0_73), .B1(n_0_118), .B2(n_0_0_74), 
      .ZN(n_0_0_34));
   INV_X1 i_0_0_62 (.A(n_0_0_35), .ZN(n_0_190));
   AOI22_X1 i_0_0_63 (.A1(n_0_380), .A2(n_0_0_73), .B1(n_0_119), .B2(n_0_0_74), 
      .ZN(n_0_0_35));
   INV_X1 i_0_0_64 (.A(n_0_0_36), .ZN(n_0_191));
   AOI22_X1 i_0_0_65 (.A1(n_0_381), .A2(n_0_0_73), .B1(n_0_120), .B2(n_0_0_74), 
      .ZN(n_0_0_36));
   INV_X1 i_0_0_66 (.A(n_0_0_37), .ZN(n_0_192));
   AOI22_X1 i_0_0_67 (.A1(n_0_382), .A2(n_0_0_73), .B1(n_0_121), .B2(n_0_0_74), 
      .ZN(n_0_0_37));
   INV_X1 i_0_0_68 (.A(n_0_0_38), .ZN(n_0_193));
   AOI22_X1 i_0_0_69 (.A1(n_0_383), .A2(n_0_0_73), .B1(n_0_122), .B2(n_0_0_74), 
      .ZN(n_0_0_38));
   INV_X1 i_0_0_70 (.A(n_0_0_39), .ZN(n_0_194));
   AOI22_X1 i_0_0_71 (.A1(n_0_384), .A2(n_0_0_73), .B1(n_0_123), .B2(n_0_0_74), 
      .ZN(n_0_0_39));
   INV_X1 i_0_0_72 (.A(n_0_0_40), .ZN(n_0_195));
   AOI22_X1 i_0_0_73 (.A1(n_0_124), .A2(n_0_0_74), .B1(n_0_385), .B2(n_0_0_73), 
      .ZN(n_0_0_40));
   INV_X1 i_0_0_74 (.A(n_0_0_41), .ZN(n_0_196));
   AOI22_X1 i_0_0_75 (.A1(n_0_125), .A2(n_0_0_74), .B1(n_0_63), .B2(n_0_0_73), 
      .ZN(n_0_0_41));
   INV_X1 i_0_0_76 (.A(n_0_0_42), .ZN(n_0_197));
   AOI22_X1 i_0_0_77 (.A1(n_0_126), .A2(n_0_0_74), .B1(n_0_64), .B2(n_0_0_73), 
      .ZN(n_0_0_42));
   INV_X1 i_0_0_78 (.A(n_0_0_43), .ZN(n_0_198));
   AOI22_X1 i_0_0_79 (.A1(n_0_127), .A2(n_0_0_74), .B1(n_0_65), .B2(n_0_0_73), 
      .ZN(n_0_0_43));
   INV_X1 i_0_0_80 (.A(n_0_0_44), .ZN(n_0_199));
   AOI22_X1 i_0_0_81 (.A1(n_0_128), .A2(n_0_0_74), .B1(n_0_66), .B2(n_0_0_73), 
      .ZN(n_0_0_44));
   INV_X1 i_0_0_82 (.A(n_0_0_45), .ZN(n_0_200));
   AOI22_X1 i_0_0_83 (.A1(n_0_129), .A2(n_0_0_74), .B1(n_0_67), .B2(n_0_0_73), 
      .ZN(n_0_0_45));
   INV_X1 i_0_0_84 (.A(n_0_0_46), .ZN(n_0_201));
   AOI22_X1 i_0_0_85 (.A1(n_0_130), .A2(n_0_0_74), .B1(n_0_68), .B2(n_0_0_73), 
      .ZN(n_0_0_46));
   INV_X1 i_0_0_86 (.A(n_0_0_47), .ZN(n_0_202));
   AOI22_X1 i_0_0_87 (.A1(n_0_131), .A2(n_0_0_74), .B1(n_0_69), .B2(n_0_0_73), 
      .ZN(n_0_0_47));
   INV_X1 i_0_0_88 (.A(n_0_0_48), .ZN(n_0_203));
   AOI22_X1 i_0_0_89 (.A1(n_0_132), .A2(n_0_0_74), .B1(n_0_70), .B2(n_0_0_73), 
      .ZN(n_0_0_48));
   INV_X1 i_0_0_90 (.A(n_0_0_49), .ZN(n_0_204));
   AOI22_X1 i_0_0_91 (.A1(n_0_133), .A2(n_0_0_74), .B1(n_0_71), .B2(n_0_0_73), 
      .ZN(n_0_0_49));
   INV_X1 i_0_0_92 (.A(n_0_0_50), .ZN(n_0_205));
   AOI22_X1 i_0_0_93 (.A1(n_0_134), .A2(n_0_0_74), .B1(n_0_72), .B2(n_0_0_73), 
      .ZN(n_0_0_50));
   INV_X1 i_0_0_94 (.A(n_0_0_51), .ZN(n_0_206));
   AOI22_X1 i_0_0_95 (.A1(n_0_135), .A2(n_0_0_74), .B1(n_0_73), .B2(n_0_0_73), 
      .ZN(n_0_0_51));
   INV_X1 i_0_0_96 (.A(n_0_0_52), .ZN(n_0_207));
   AOI22_X1 i_0_0_97 (.A1(n_0_136), .A2(n_0_0_74), .B1(n_0_74), .B2(n_0_0_73), 
      .ZN(n_0_0_52));
   INV_X1 i_0_0_98 (.A(n_0_0_53), .ZN(n_0_208));
   AOI22_X1 i_0_0_99 (.A1(n_0_137), .A2(n_0_0_74), .B1(n_0_75), .B2(n_0_0_73), 
      .ZN(n_0_0_53));
   INV_X1 i_0_0_100 (.A(n_0_0_54), .ZN(n_0_209));
   AOI22_X1 i_0_0_101 (.A1(n_0_138), .A2(n_0_0_74), .B1(n_0_76), .B2(n_0_0_73), 
      .ZN(n_0_0_54));
   INV_X1 i_0_0_102 (.A(n_0_0_55), .ZN(n_0_210));
   AOI22_X1 i_0_0_103 (.A1(n_0_139), .A2(n_0_0_74), .B1(n_0_77), .B2(n_0_0_73), 
      .ZN(n_0_0_55));
   INV_X1 i_0_0_104 (.A(n_0_0_56), .ZN(n_0_211));
   AOI22_X1 i_0_0_105 (.A1(n_0_140), .A2(n_0_0_74), .B1(n_0_78), .B2(n_0_0_73), 
      .ZN(n_0_0_56));
   INV_X1 i_0_0_106 (.A(n_0_0_57), .ZN(n_0_212));
   AOI22_X1 i_0_0_107 (.A1(n_0_141), .A2(n_0_0_74), .B1(n_0_79), .B2(n_0_0_73), 
      .ZN(n_0_0_57));
   INV_X1 i_0_0_108 (.A(n_0_0_58), .ZN(n_0_213));
   AOI22_X1 i_0_0_109 (.A1(n_0_142), .A2(n_0_0_74), .B1(n_0_80), .B2(n_0_0_73), 
      .ZN(n_0_0_58));
   INV_X1 i_0_0_110 (.A(n_0_0_59), .ZN(n_0_214));
   AOI22_X1 i_0_0_111 (.A1(n_0_143), .A2(n_0_0_74), .B1(n_0_81), .B2(n_0_0_73), 
      .ZN(n_0_0_59));
   INV_X1 i_0_0_112 (.A(n_0_0_60), .ZN(n_0_215));
   AOI22_X1 i_0_0_113 (.A1(n_0_144), .A2(n_0_0_74), .B1(n_0_82), .B2(n_0_0_73), 
      .ZN(n_0_0_60));
   INV_X1 i_0_0_114 (.A(n_0_0_61), .ZN(n_0_216));
   AOI22_X1 i_0_0_115 (.A1(n_0_145), .A2(n_0_0_74), .B1(n_0_83), .B2(n_0_0_73), 
      .ZN(n_0_0_61));
   INV_X1 i_0_0_116 (.A(n_0_0_62), .ZN(n_0_217));
   AOI22_X1 i_0_0_117 (.A1(n_0_146), .A2(n_0_0_74), .B1(n_0_84), .B2(n_0_0_73), 
      .ZN(n_0_0_62));
   INV_X1 i_0_0_118 (.A(n_0_0_63), .ZN(n_0_218));
   AOI22_X1 i_0_0_119 (.A1(n_0_147), .A2(n_0_0_74), .B1(n_0_85), .B2(n_0_0_73), 
      .ZN(n_0_0_63));
   INV_X1 i_0_0_120 (.A(n_0_0_64), .ZN(n_0_219));
   AOI22_X1 i_0_0_121 (.A1(n_0_148), .A2(n_0_0_74), .B1(n_0_86), .B2(n_0_0_73), 
      .ZN(n_0_0_64));
   INV_X1 i_0_0_122 (.A(n_0_0_65), .ZN(n_0_220));
   AOI22_X1 i_0_0_123 (.A1(n_0_149), .A2(n_0_0_74), .B1(n_0_87), .B2(n_0_0_73), 
      .ZN(n_0_0_65));
   INV_X1 i_0_0_124 (.A(n_0_0_66), .ZN(n_0_221));
   AOI22_X1 i_0_0_125 (.A1(n_0_150), .A2(n_0_0_74), .B1(n_0_88), .B2(n_0_0_73), 
      .ZN(n_0_0_66));
   INV_X1 i_0_0_126 (.A(n_0_0_67), .ZN(n_0_222));
   AOI22_X1 i_0_0_127 (.A1(n_0_151), .A2(n_0_0_74), .B1(n_0_89), .B2(n_0_0_73), 
      .ZN(n_0_0_67));
   INV_X1 i_0_0_128 (.A(n_0_0_68), .ZN(n_0_223));
   AOI22_X1 i_0_0_129 (.A1(n_0_152), .A2(n_0_0_74), .B1(n_0_90), .B2(n_0_0_73), 
      .ZN(n_0_0_68));
   INV_X1 i_0_0_130 (.A(n_0_0_69), .ZN(n_0_224));
   AOI22_X1 i_0_0_131 (.A1(n_0_153), .A2(n_0_0_74), .B1(n_0_91), .B2(n_0_0_73), 
      .ZN(n_0_0_69));
   AND2_X1 i_0_0_139 (.A1(n_0_157), .A2(n_0_0_74), .ZN(n_0_228));
   AND2_X1 i_0_0_141 (.A1(n_0_0_157), .A2(n_0_64), .ZN(n_0_229));
   AND2_X1 i_0_0_142 (.A1(n_0_0_157), .A2(n_0_65), .ZN(n_0_230));
   AND2_X1 i_0_0_143 (.A1(n_0_0_157), .A2(n_0_66), .ZN(n_0_231));
   AND2_X1 i_0_0_144 (.A1(n_0_0_157), .A2(n_0_67), .ZN(n_0_232));
   AND2_X1 i_0_0_145 (.A1(n_0_0_157), .A2(n_0_68), .ZN(n_0_233));
   AND2_X1 i_0_0_146 (.A1(n_0_0_157), .A2(n_0_69), .ZN(n_0_234));
   AND2_X1 i_0_0_147 (.A1(n_0_0_157), .A2(n_0_70), .ZN(n_0_235));
   AND2_X1 i_0_0_148 (.A1(n_0_0_157), .A2(n_0_71), .ZN(n_0_236));
   AND2_X1 i_0_0_149 (.A1(n_0_0_157), .A2(n_0_72), .ZN(n_0_237));
   AND2_X1 i_0_0_150 (.A1(n_0_0_157), .A2(n_0_73), .ZN(n_0_238));
   AND2_X1 i_0_0_151 (.A1(n_0_0_157), .A2(n_0_74), .ZN(n_0_239));
   AND2_X1 i_0_0_152 (.A1(n_0_0_157), .A2(n_0_75), .ZN(n_0_240));
   AND2_X1 i_0_0_153 (.A1(n_0_0_157), .A2(n_0_76), .ZN(n_0_241));
   AND2_X1 i_0_0_154 (.A1(n_0_0_157), .A2(n_0_77), .ZN(n_0_242));
   AND2_X1 i_0_0_155 (.A1(n_0_0_157), .A2(n_0_78), .ZN(n_0_243));
   AND2_X1 i_0_0_156 (.A1(n_0_0_157), .A2(n_0_79), .ZN(n_0_244));
   AND2_X1 i_0_0_157 (.A1(n_0_0_157), .A2(n_0_80), .ZN(n_0_245));
   AND2_X1 i_0_0_158 (.A1(n_0_0_157), .A2(n_0_81), .ZN(n_0_246));
   AND2_X1 i_0_0_159 (.A1(n_0_0_157), .A2(n_0_82), .ZN(n_0_247));
   AND2_X1 i_0_0_160 (.A1(n_0_0_157), .A2(n_0_83), .ZN(n_0_248));
   AND2_X1 i_0_0_161 (.A1(n_0_0_157), .A2(n_0_84), .ZN(n_0_249));
   AND2_X1 i_0_0_162 (.A1(n_0_0_157), .A2(n_0_85), .ZN(n_0_250));
   AND2_X1 i_0_0_163 (.A1(n_0_0_157), .A2(n_0_86), .ZN(n_0_251));
   AND2_X1 i_0_0_164 (.A1(n_0_0_157), .A2(n_0_87), .ZN(n_0_252));
   AND2_X1 i_0_0_165 (.A1(n_0_0_157), .A2(n_0_88), .ZN(n_0_253));
   AND2_X1 i_0_0_166 (.A1(n_0_0_157), .A2(n_0_89), .ZN(n_0_254));
   AND2_X1 i_0_0_167 (.A1(n_0_0_157), .A2(n_0_90), .ZN(n_0_255));
   AND2_X1 i_0_0_168 (.A1(n_0_0_157), .A2(n_0_91), .ZN(n_0_256));
   AND2_X1 i_0_0_169 (.A1(n_0_0_157), .A2(n_0_92), .ZN(n_0_257));
   AND2_X1 i_0_0_170 (.A1(n_0_0_157), .A2(n_0_93), .ZN(n_0_258));
   AND2_X1 i_0_0_171 (.A1(n_0_0_157), .A2(n_0_94), .ZN(n_0_259));
   NOR2_X1 i_0_0_172 (.A1(rst), .A2(n_0_0_76), .ZN(n_0_260));
   NOR2_X1 i_0_0_173 (.A1(rst), .A2(n_0_0_77), .ZN(n_0_261));
   NOR2_X1 i_0_0_174 (.A1(rst), .A2(n_0_0_78), .ZN(n_0_262));
   NOR2_X1 i_0_0_175 (.A1(rst), .A2(n_0_0_79), .ZN(n_0_263));
   NOR2_X1 i_0_0_176 (.A1(rst), .A2(n_0_0_80), .ZN(n_0_264));
   NOR2_X1 i_0_0_177 (.A1(rst), .A2(n_0_0_81), .ZN(n_0_265));
   NOR2_X1 i_0_0_178 (.A1(rst), .A2(n_0_0_82), .ZN(n_0_266));
   NOR2_X1 i_0_0_179 (.A1(rst), .A2(n_0_0_83), .ZN(n_0_267));
   NOR2_X1 i_0_0_180 (.A1(rst), .A2(n_0_0_84), .ZN(n_0_268));
   NOR2_X1 i_0_0_181 (.A1(rst), .A2(n_0_0_85), .ZN(n_0_269));
   NOR2_X1 i_0_0_182 (.A1(rst), .A2(n_0_0_86), .ZN(n_0_270));
   NOR2_X1 i_0_0_183 (.A1(rst), .A2(n_0_0_87), .ZN(n_0_271));
   NOR2_X1 i_0_0_184 (.A1(rst), .A2(n_0_0_88), .ZN(n_0_272));
   NOR2_X1 i_0_0_185 (.A1(rst), .A2(n_0_0_89), .ZN(n_0_273));
   NOR2_X1 i_0_0_186 (.A1(rst), .A2(n_0_0_90), .ZN(n_0_274));
   NOR2_X1 i_0_0_187 (.A1(rst), .A2(n_0_0_91), .ZN(n_0_275));
   NOR2_X1 i_0_0_188 (.A1(rst), .A2(n_0_0_92), .ZN(n_0_276));
   NOR2_X1 i_0_0_189 (.A1(rst), .A2(n_0_0_93), .ZN(n_0_277));
   NOR2_X1 i_0_0_190 (.A1(rst), .A2(n_0_0_94), .ZN(n_0_278));
   NOR2_X1 i_0_0_191 (.A1(rst), .A2(n_0_0_95), .ZN(n_0_279));
   NOR2_X1 i_0_0_192 (.A1(rst), .A2(n_0_0_96), .ZN(n_0_280));
   NOR2_X1 i_0_0_193 (.A1(rst), .A2(n_0_0_97), .ZN(n_0_281));
   NOR2_X1 i_0_0_194 (.A1(rst), .A2(n_0_0_98), .ZN(n_0_282));
   NOR2_X1 i_0_0_195 (.A1(rst), .A2(n_0_0_99), .ZN(n_0_283));
   NOR2_X1 i_0_0_196 (.A1(rst), .A2(n_0_0_100), .ZN(n_0_284));
   NOR2_X1 i_0_0_197 (.A1(rst), .A2(n_0_0_101), .ZN(n_0_285));
   NOR2_X1 i_0_0_198 (.A1(rst), .A2(n_0_0_102), .ZN(n_0_286));
   NOR2_X1 i_0_0_199 (.A1(rst), .A2(n_0_0_103), .ZN(n_0_287));
   NOR2_X1 i_0_0_200 (.A1(rst), .A2(n_0_0_104), .ZN(n_0_288));
   NOR2_X1 i_0_0_201 (.A1(rst), .A2(n_0_0_105), .ZN(n_0_289));
   NOR2_X1 i_0_0_202 (.A1(rst), .A2(n_0_0_107), .ZN(n_0_290));
   AND2_X1 i_0_0_203 (.A1(n_0_0_157), .A2(n_0_63), .ZN(n_0_291));
   AND2_X1 i_0_0_204 (.A1(Accumulator[0]), .A2(n_0_0_144), .ZN(n_0_292));
   AND2_X1 i_0_0_205 (.A1(Accumulator[1]), .A2(n_0_0_144), .ZN(n_0_293));
   AND2_X1 i_0_0_206 (.A1(Accumulator[2]), .A2(n_0_0_144), .ZN(n_0_294));
   AND2_X1 i_0_0_207 (.A1(Accumulator[3]), .A2(n_0_0_144), .ZN(n_0_295));
   AND2_X1 i_0_0_208 (.A1(Accumulator[4]), .A2(n_0_0_144), .ZN(n_0_296));
   AND2_X1 i_0_0_209 (.A1(Accumulator[5]), .A2(n_0_0_144), .ZN(n_0_297));
   AND2_X1 i_0_0_210 (.A1(Accumulator[6]), .A2(n_0_0_144), .ZN(n_0_298));
   AND2_X1 i_0_0_211 (.A1(Accumulator[7]), .A2(n_0_0_144), .ZN(n_0_299));
   AND2_X1 i_0_0_212 (.A1(Accumulator[8]), .A2(n_0_0_144), .ZN(n_0_300));
   AND2_X1 i_0_0_213 (.A1(Accumulator[9]), .A2(n_0_0_144), .ZN(n_0_301));
   AND2_X1 i_0_0_214 (.A1(Accumulator[10]), .A2(n_0_0_144), .ZN(n_0_302));
   AND2_X1 i_0_0_215 (.A1(Accumulator[11]), .A2(n_0_0_144), .ZN(n_0_303));
   AND2_X1 i_0_0_216 (.A1(Accumulator[12]), .A2(n_0_0_144), .ZN(n_0_304));
   AND2_X1 i_0_0_217 (.A1(Accumulator[13]), .A2(n_0_0_144), .ZN(n_0_305));
   AND2_X1 i_0_0_218 (.A1(Accumulator[14]), .A2(n_0_0_144), .ZN(n_0_306));
   AND2_X1 i_0_0_219 (.A1(Accumulator[15]), .A2(n_0_0_144), .ZN(n_0_307));
   AND2_X1 i_0_0_220 (.A1(Accumulator[16]), .A2(n_0_0_144), .ZN(n_0_308));
   AND2_X1 i_0_0_221 (.A1(Accumulator[17]), .A2(n_0_0_144), .ZN(n_0_309));
   AND2_X1 i_0_0_222 (.A1(Accumulator[18]), .A2(n_0_0_144), .ZN(n_0_310));
   AND2_X1 i_0_0_223 (.A1(Accumulator[19]), .A2(n_0_0_144), .ZN(n_0_311));
   AND2_X1 i_0_0_224 (.A1(Accumulator[20]), .A2(n_0_0_144), .ZN(n_0_312));
   AND2_X1 i_0_0_225 (.A1(Accumulator[21]), .A2(n_0_0_144), .ZN(n_0_313));
   AND2_X1 i_0_0_226 (.A1(Accumulator[22]), .A2(n_0_0_144), .ZN(n_0_314));
   AND2_X1 i_0_0_227 (.A1(Accumulator[23]), .A2(n_0_0_144), .ZN(n_0_315));
   AND2_X1 i_0_0_228 (.A1(Accumulator[24]), .A2(n_0_0_144), .ZN(n_0_316));
   AND2_X1 i_0_0_229 (.A1(Accumulator[25]), .A2(n_0_0_144), .ZN(n_0_317));
   AND2_X1 i_0_0_230 (.A1(Accumulator[26]), .A2(n_0_0_144), .ZN(n_0_318));
   AND2_X1 i_0_0_231 (.A1(Accumulator[27]), .A2(n_0_0_144), .ZN(n_0_319));
   AND2_X1 i_0_0_232 (.A1(Accumulator[28]), .A2(n_0_0_144), .ZN(n_0_320));
   AND2_X1 i_0_0_233 (.A1(Accumulator[29]), .A2(n_0_0_144), .ZN(n_0_321));
   AND2_X1 i_0_0_234 (.A1(Accumulator[30]), .A2(n_0_0_144), .ZN(n_0_322));
   NOR2_X1 i_0_0_235 (.A1(n_0_0_109), .A2(n_0_0_75), .ZN(n_0_323));
   NOR2_X1 i_0_0_236 (.A1(n_0_0_110), .A2(n_0_0_75), .ZN(n_0_324));
   NOR2_X1 i_0_0_237 (.A1(n_0_0_111), .A2(n_0_0_75), .ZN(n_0_325));
   NOR2_X1 i_0_0_238 (.A1(n_0_0_112), .A2(n_0_0_75), .ZN(n_0_326));
   NOR2_X1 i_0_0_239 (.A1(n_0_0_113), .A2(n_0_0_75), .ZN(n_0_327));
   NOR2_X1 i_0_0_240 (.A1(n_0_0_114), .A2(n_0_0_75), .ZN(n_0_328));
   NOR2_X1 i_0_0_241 (.A1(n_0_0_115), .A2(n_0_0_75), .ZN(n_0_329));
   NOR2_X1 i_0_0_242 (.A1(n_0_0_116), .A2(n_0_0_75), .ZN(n_0_330));
   NOR2_X1 i_0_0_243 (.A1(n_0_0_117), .A2(n_0_0_75), .ZN(n_0_331));
   NOR2_X1 i_0_0_244 (.A1(n_0_0_118), .A2(n_0_0_75), .ZN(n_0_332));
   NOR2_X1 i_0_0_245 (.A1(n_0_0_119), .A2(n_0_0_75), .ZN(n_0_333));
   NOR2_X1 i_0_0_246 (.A1(n_0_0_120), .A2(n_0_0_75), .ZN(n_0_334));
   NOR2_X1 i_0_0_247 (.A1(n_0_0_121), .A2(n_0_0_75), .ZN(n_0_335));
   NOR2_X1 i_0_0_248 (.A1(n_0_0_122), .A2(n_0_0_75), .ZN(n_0_336));
   NOR2_X1 i_0_0_249 (.A1(n_0_0_123), .A2(n_0_0_75), .ZN(n_0_337));
   NOR2_X1 i_0_0_250 (.A1(n_0_0_124), .A2(n_0_0_75), .ZN(n_0_338));
   NOR2_X1 i_0_0_251 (.A1(n_0_0_125), .A2(n_0_0_75), .ZN(n_0_339));
   NOR2_X1 i_0_0_252 (.A1(n_0_0_126), .A2(n_0_0_75), .ZN(n_0_340));
   NOR2_X1 i_0_0_253 (.A1(n_0_0_127), .A2(n_0_0_75), .ZN(n_0_341));
   NOR2_X1 i_0_0_254 (.A1(n_0_0_128), .A2(n_0_0_75), .ZN(n_0_342));
   NOR2_X1 i_0_0_255 (.A1(n_0_0_129), .A2(n_0_0_75), .ZN(n_0_343));
   NOR2_X1 i_0_0_256 (.A1(n_0_0_130), .A2(n_0_0_75), .ZN(n_0_344));
   NOR2_X1 i_0_0_257 (.A1(n_0_0_131), .A2(n_0_0_75), .ZN(n_0_345));
   NOR2_X1 i_0_0_258 (.A1(n_0_0_132), .A2(n_0_0_75), .ZN(n_0_346));
   NOR2_X1 i_0_0_259 (.A1(n_0_0_133), .A2(n_0_0_75), .ZN(n_0_347));
   NOR2_X1 i_0_0_260 (.A1(n_0_0_134), .A2(n_0_0_75), .ZN(n_0_348));
   NOR2_X1 i_0_0_261 (.A1(n_0_0_135), .A2(n_0_0_75), .ZN(n_0_349));
   NOR2_X1 i_0_0_262 (.A1(n_0_0_136), .A2(n_0_0_75), .ZN(n_0_350));
   NOR2_X1 i_0_0_263 (.A1(n_0_0_137), .A2(n_0_0_75), .ZN(n_0_351));
   NOR2_X1 i_0_0_264 (.A1(n_0_0_138), .A2(n_0_0_75), .ZN(n_0_352));
   NOR2_X1 i_0_0_265 (.A1(n_0_0_139), .A2(n_0_0_75), .ZN(n_0_353));
   NOR2_X1 i_0_0_266 (.A1(n_0_0_141), .A2(n_0_0_75), .ZN(n_0_354));
   AOI22_X1 i_0_0_267 (.A1(B_r[0]), .A2(n_0_0_144), .B1(b[0]), .B2(n_0_0_143), 
      .ZN(n_0_0_75));
   INV_X1 i_0_0_268 (.A(n_0_0_76), .ZN(n_0_355));
   AOI222_X1 i_0_0_269 (.A1(B_r[1]), .A2(n_0_0_144), .B1(n_0_32), .B2(n_0_0_108), 
      .C1(b[1]), .C2(n_0_0_106), .ZN(n_0_0_76));
   INV_X1 i_0_0_272 (.A(n_0_0_78), .ZN(n_0_357));
   AOI222_X1 i_0_0_273 (.A1(B_r[3]), .A2(n_0_0_144), .B1(n_0_34), .B2(n_0_0_108), 
      .C1(b[3]), .C2(n_0_0_106), .ZN(n_0_0_78));
   INV_X1 i_0_0_274 (.A(n_0_0_79), .ZN(n_0_358));
   AOI222_X1 i_0_0_275 (.A1(B_r[4]), .A2(n_0_0_144), .B1(n_0_35), .B2(n_0_0_108), 
      .C1(b[4]), .C2(n_0_0_106), .ZN(n_0_0_79));
   INV_X1 i_0_0_276 (.A(n_0_0_80), .ZN(n_0_359));
   AOI222_X1 i_0_0_277 (.A1(B_r[5]), .A2(n_0_0_144), .B1(n_0_36), .B2(n_0_0_108), 
      .C1(b[5]), .C2(n_0_0_106), .ZN(n_0_0_80));
   INV_X1 i_0_0_278 (.A(n_0_0_81), .ZN(n_0_360));
   AOI222_X1 i_0_0_279 (.A1(B_r[6]), .A2(n_0_0_144), .B1(n_0_37), .B2(n_0_0_108), 
      .C1(b[6]), .C2(n_0_0_106), .ZN(n_0_0_81));
   INV_X1 i_0_0_292 (.A(n_0_0_88), .ZN(n_0_367));
   AOI222_X1 i_0_0_293 (.A1(B_r[13]), .A2(n_0_0_144), .B1(n_0_44), .B2(n_0_0_108), 
      .C1(b[13]), .C2(n_0_0_106), .ZN(n_0_0_88));
   INV_X1 i_0_0_294 (.A(n_0_0_89), .ZN(n_0_368));
   AOI222_X1 i_0_0_295 (.A1(B_r[14]), .A2(n_0_0_144), .B1(n_0_45), .B2(n_0_0_108), 
      .C1(b[14]), .C2(n_0_0_106), .ZN(n_0_0_89));
   INV_X1 i_0_0_296 (.A(n_0_0_90), .ZN(n_0_369));
   AOI222_X1 i_0_0_297 (.A1(B_r[15]), .A2(n_0_0_144), .B1(n_0_46), .B2(n_0_0_108), 
      .C1(b[15]), .C2(n_0_0_106), .ZN(n_0_0_90));
   INV_X1 i_0_0_298 (.A(n_0_0_91), .ZN(n_0_370));
   AOI222_X1 i_0_0_299 (.A1(B_r[16]), .A2(n_0_0_144), .B1(n_0_47), .B2(n_0_0_108), 
      .C1(b[16]), .C2(n_0_0_106), .ZN(n_0_0_91));
   INV_X1 i_0_0_300 (.A(n_0_0_92), .ZN(n_0_371));
   AOI222_X1 i_0_0_301 (.A1(B_r[17]), .A2(n_0_0_144), .B1(n_0_48), .B2(n_0_0_108), 
      .C1(b[17]), .C2(n_0_0_106), .ZN(n_0_0_92));
   INV_X1 i_0_0_302 (.A(n_0_0_93), .ZN(n_0_372));
   AOI222_X1 i_0_0_303 (.A1(B_r[18]), .A2(n_0_0_144), .B1(n_0_49), .B2(n_0_0_108), 
      .C1(b[18]), .C2(n_0_0_106), .ZN(n_0_0_93));
   INV_X1 i_0_0_304 (.A(n_0_0_94), .ZN(n_0_373));
   AOI222_X1 i_0_0_305 (.A1(B_r[19]), .A2(n_0_0_144), .B1(n_0_50), .B2(n_0_0_108), 
      .C1(b[19]), .C2(n_0_0_106), .ZN(n_0_0_94));
   INV_X1 i_0_0_306 (.A(n_0_0_95), .ZN(n_0_374));
   AOI222_X1 i_0_0_307 (.A1(B_r[20]), .A2(n_0_0_144), .B1(n_0_51), .B2(n_0_0_108), 
      .C1(b[20]), .C2(n_0_0_106), .ZN(n_0_0_95));
   INV_X1 i_0_0_308 (.A(n_0_0_96), .ZN(n_0_375));
   AOI222_X1 i_0_0_309 (.A1(B_r[21]), .A2(n_0_0_144), .B1(n_0_52), .B2(n_0_0_108), 
      .C1(b[21]), .C2(n_0_0_106), .ZN(n_0_0_96));
   INV_X1 i_0_0_310 (.A(n_0_0_97), .ZN(n_0_376));
   AOI222_X1 i_0_0_311 (.A1(B_r[22]), .A2(n_0_0_144), .B1(n_0_53), .B2(n_0_0_108), 
      .C1(b[22]), .C2(n_0_0_106), .ZN(n_0_0_97));
   INV_X1 i_0_0_312 (.A(n_0_0_98), .ZN(n_0_377));
   AOI222_X1 i_0_0_313 (.A1(B_r[23]), .A2(n_0_0_144), .B1(n_0_54), .B2(n_0_0_108), 
      .C1(b[23]), .C2(n_0_0_106), .ZN(n_0_0_98));
   INV_X1 i_0_0_314 (.A(n_0_0_99), .ZN(n_0_378));
   AOI222_X1 i_0_0_315 (.A1(B_r[24]), .A2(n_0_0_144), .B1(n_0_55), .B2(n_0_0_108), 
      .C1(b[24]), .C2(n_0_0_106), .ZN(n_0_0_99));
   INV_X1 i_0_0_316 (.A(n_0_0_100), .ZN(n_0_379));
   AOI222_X1 i_0_0_317 (.A1(B_r[25]), .A2(n_0_0_144), .B1(n_0_56), .B2(n_0_0_108), 
      .C1(b[25]), .C2(n_0_0_106), .ZN(n_0_0_100));
   INV_X1 i_0_0_318 (.A(n_0_0_101), .ZN(n_0_380));
   AOI222_X1 i_0_0_319 (.A1(B_r[26]), .A2(n_0_0_144), .B1(n_0_57), .B2(n_0_0_108), 
      .C1(b[26]), .C2(n_0_0_106), .ZN(n_0_0_101));
   INV_X1 i_0_0_320 (.A(n_0_0_102), .ZN(n_0_381));
   AOI222_X1 i_0_0_321 (.A1(B_r[27]), .A2(n_0_0_144), .B1(n_0_58), .B2(n_0_0_108), 
      .C1(b[27]), .C2(n_0_0_106), .ZN(n_0_0_102));
   INV_X1 i_0_0_322 (.A(n_0_0_103), .ZN(n_0_382));
   AOI222_X1 i_0_0_323 (.A1(B_r[28]), .A2(n_0_0_144), .B1(n_0_59), .B2(n_0_0_108), 
      .C1(b[28]), .C2(n_0_0_106), .ZN(n_0_0_103));
   INV_X1 i_0_0_324 (.A(n_0_0_104), .ZN(n_0_383));
   AOI222_X1 i_0_0_325 (.A1(B_r[29]), .A2(n_0_0_144), .B1(n_0_60), .B2(n_0_0_108), 
      .C1(b[29]), .C2(n_0_0_106), .ZN(n_0_0_104));
   INV_X1 i_0_0_326 (.A(n_0_0_105), .ZN(n_0_384));
   AOI222_X1 i_0_0_327 (.A1(B_r[30]), .A2(n_0_0_144), .B1(n_0_61), .B2(n_0_0_108), 
      .C1(b[30]), .C2(n_0_0_106), .ZN(n_0_0_105));
   INV_X1 i_0_0_329 (.A(n_0_0_107), .ZN(n_0_385));
   AOI22_X1 i_0_0_330 (.A1(B_r[31]), .A2(n_0_0_144), .B1(n_0_62), .B2(n_0_0_108), 
      .ZN(n_0_0_107));
   NOR2_X1 i_0_0_332 (.A1(rst), .A2(n_0_0_109), .ZN(n_0_386));
   AOI22_X1 i_0_0_333 (.A1(A_r[0]), .A2(n_0_0_144), .B1(a[0]), .B2(n_0_0_143), 
      .ZN(n_0_0_109));
   NOR2_X1 i_0_0_334 (.A1(rst), .A2(n_0_0_110), .ZN(n_0_387));
   AOI222_X1 i_0_0_335 (.A1(A_r[1]), .A2(n_0_0_144), .B1(a[1]), .B2(n_0_0_140), 
      .C1(n_0_1), .C2(n_0_0_142), .ZN(n_0_0_110));
   NOR2_X1 i_0_0_336 (.A1(rst), .A2(n_0_0_111), .ZN(n_0_388));
   AOI222_X1 i_0_0_337 (.A1(A_r[2]), .A2(n_0_0_144), .B1(a[2]), .B2(n_0_0_140), 
      .C1(n_0_2), .C2(n_0_0_142), .ZN(n_0_0_111));
   NOR2_X1 i_0_0_338 (.A1(rst), .A2(n_0_0_112), .ZN(n_0_389));
   AOI222_X1 i_0_0_339 (.A1(A_r[3]), .A2(n_0_0_144), .B1(a[3]), .B2(n_0_0_140), 
      .C1(n_0_3), .C2(n_0_0_142), .ZN(n_0_0_112));
   NOR2_X1 i_0_0_340 (.A1(rst), .A2(n_0_0_113), .ZN(n_0_390));
   AOI222_X1 i_0_0_341 (.A1(A_r[4]), .A2(n_0_0_144), .B1(a[4]), .B2(n_0_0_140), 
      .C1(n_0_4), .C2(n_0_0_142), .ZN(n_0_0_113));
   NOR2_X1 i_0_0_342 (.A1(rst), .A2(n_0_0_114), .ZN(n_0_391));
   AOI222_X1 i_0_0_343 (.A1(A_r[5]), .A2(n_0_0_144), .B1(a[5]), .B2(n_0_0_140), 
      .C1(n_0_5), .C2(n_0_0_142), .ZN(n_0_0_114));
   NOR2_X1 i_0_0_344 (.A1(rst), .A2(n_0_0_115), .ZN(n_0_392));
   AOI222_X1 i_0_0_345 (.A1(A_r[6]), .A2(n_0_0_144), .B1(a[6]), .B2(n_0_0_140), 
      .C1(n_0_6), .C2(n_0_0_142), .ZN(n_0_0_115));
   NOR2_X1 i_0_0_346 (.A1(rst), .A2(n_0_0_116), .ZN(n_0_393));
   AOI222_X1 i_0_0_347 (.A1(A_r[7]), .A2(n_0_0_144), .B1(a[7]), .B2(n_0_0_140), 
      .C1(n_0_7), .C2(n_0_0_142), .ZN(n_0_0_116));
   NOR2_X1 i_0_0_348 (.A1(rst), .A2(n_0_0_117), .ZN(n_0_394));
   AOI222_X1 i_0_0_349 (.A1(A_r[8]), .A2(n_0_0_144), .B1(a[8]), .B2(n_0_0_140), 
      .C1(n_0_8), .C2(n_0_0_142), .ZN(n_0_0_117));
   NOR2_X1 i_0_0_350 (.A1(rst), .A2(n_0_0_118), .ZN(n_0_395));
   AOI222_X1 i_0_0_351 (.A1(A_r[9]), .A2(n_0_0_144), .B1(a[9]), .B2(n_0_0_140), 
      .C1(n_0_9), .C2(n_0_0_142), .ZN(n_0_0_118));
   NOR2_X1 i_0_0_352 (.A1(rst), .A2(n_0_0_119), .ZN(n_0_396));
   AOI222_X1 i_0_0_353 (.A1(A_r[10]), .A2(n_0_0_144), .B1(a[10]), .B2(n_0_0_140), 
      .C1(n_0_10), .C2(n_0_0_142), .ZN(n_0_0_119));
   NOR2_X1 i_0_0_354 (.A1(rst), .A2(n_0_0_120), .ZN(n_0_397));
   AOI222_X1 i_0_0_355 (.A1(A_r[11]), .A2(n_0_0_144), .B1(a[11]), .B2(n_0_0_140), 
      .C1(n_0_11), .C2(n_0_0_142), .ZN(n_0_0_120));
   NOR2_X1 i_0_0_356 (.A1(rst), .A2(n_0_0_121), .ZN(n_0_398));
   AOI222_X1 i_0_0_357 (.A1(A_r[12]), .A2(n_0_0_144), .B1(a[12]), .B2(n_0_0_140), 
      .C1(n_0_12), .C2(n_0_0_142), .ZN(n_0_0_121));
   NOR2_X1 i_0_0_358 (.A1(rst), .A2(n_0_0_122), .ZN(n_0_399));
   AOI222_X1 i_0_0_359 (.A1(A_r[13]), .A2(n_0_0_144), .B1(a[13]), .B2(n_0_0_140), 
      .C1(n_0_13), .C2(n_0_0_142), .ZN(n_0_0_122));
   NOR2_X1 i_0_0_360 (.A1(rst), .A2(n_0_0_123), .ZN(n_0_400));
   AOI222_X1 i_0_0_361 (.A1(A_r[14]), .A2(n_0_0_144), .B1(a[14]), .B2(n_0_0_140), 
      .C1(n_0_14), .C2(n_0_0_142), .ZN(n_0_0_123));
   NOR2_X1 i_0_0_362 (.A1(rst), .A2(n_0_0_124), .ZN(n_0_401));
   AOI222_X1 i_0_0_363 (.A1(A_r[15]), .A2(n_0_0_144), .B1(a[15]), .B2(n_0_0_140), 
      .C1(n_0_15), .C2(n_0_0_142), .ZN(n_0_0_124));
   NOR2_X1 i_0_0_364 (.A1(rst), .A2(n_0_0_125), .ZN(n_0_402));
   AOI222_X1 i_0_0_365 (.A1(A_r[16]), .A2(n_0_0_144), .B1(a[16]), .B2(n_0_0_140), 
      .C1(n_0_16), .C2(n_0_0_142), .ZN(n_0_0_125));
   NOR2_X1 i_0_0_366 (.A1(rst), .A2(n_0_0_126), .ZN(n_0_403));
   AOI222_X1 i_0_0_367 (.A1(A_r[17]), .A2(n_0_0_144), .B1(a[17]), .B2(n_0_0_140), 
      .C1(n_0_17), .C2(n_0_0_142), .ZN(n_0_0_126));
   NOR2_X1 i_0_0_368 (.A1(rst), .A2(n_0_0_127), .ZN(n_0_404));
   AOI222_X1 i_0_0_369 (.A1(A_r[18]), .A2(n_0_0_144), .B1(a[18]), .B2(n_0_0_140), 
      .C1(n_0_18), .C2(n_0_0_142), .ZN(n_0_0_127));
   NOR2_X1 i_0_0_370 (.A1(rst), .A2(n_0_0_128), .ZN(n_0_405));
   AOI222_X1 i_0_0_371 (.A1(A_r[19]), .A2(n_0_0_144), .B1(a[19]), .B2(n_0_0_140), 
      .C1(n_0_19), .C2(n_0_0_142), .ZN(n_0_0_128));
   NOR2_X1 i_0_0_372 (.A1(rst), .A2(n_0_0_129), .ZN(n_0_406));
   AOI222_X1 i_0_0_373 (.A1(A_r[20]), .A2(n_0_0_144), .B1(a[20]), .B2(n_0_0_140), 
      .C1(n_0_20), .C2(n_0_0_142), .ZN(n_0_0_129));
   NOR2_X1 i_0_0_374 (.A1(rst), .A2(n_0_0_130), .ZN(n_0_407));
   AOI222_X1 i_0_0_375 (.A1(A_r[21]), .A2(n_0_0_144), .B1(a[21]), .B2(n_0_0_140), 
      .C1(n_0_21), .C2(n_0_0_142), .ZN(n_0_0_130));
   NOR2_X1 i_0_0_376 (.A1(rst), .A2(n_0_0_131), .ZN(n_0_408));
   AOI222_X1 i_0_0_377 (.A1(A_r[22]), .A2(n_0_0_144), .B1(a[22]), .B2(n_0_0_140), 
      .C1(n_0_22), .C2(n_0_0_142), .ZN(n_0_0_131));
   NOR2_X1 i_0_0_378 (.A1(rst), .A2(n_0_0_132), .ZN(n_0_409));
   AOI222_X1 i_0_0_379 (.A1(A_r[23]), .A2(n_0_0_144), .B1(a[23]), .B2(n_0_0_140), 
      .C1(n_0_23), .C2(n_0_0_142), .ZN(n_0_0_132));
   NOR2_X1 i_0_0_380 (.A1(rst), .A2(n_0_0_133), .ZN(n_0_410));
   AOI222_X1 i_0_0_381 (.A1(A_r[24]), .A2(n_0_0_144), .B1(a[24]), .B2(n_0_0_140), 
      .C1(n_0_24), .C2(n_0_0_142), .ZN(n_0_0_133));
   NOR2_X1 i_0_0_382 (.A1(rst), .A2(n_0_0_134), .ZN(n_0_411));
   AOI222_X1 i_0_0_383 (.A1(A_r[25]), .A2(n_0_0_144), .B1(a[25]), .B2(n_0_0_140), 
      .C1(n_0_25), .C2(n_0_0_142), .ZN(n_0_0_134));
   NOR2_X1 i_0_0_384 (.A1(rst), .A2(n_0_0_135), .ZN(n_0_412));
   AOI222_X1 i_0_0_385 (.A1(A_r[26]), .A2(n_0_0_144), .B1(a[26]), .B2(n_0_0_140), 
      .C1(n_0_26), .C2(n_0_0_142), .ZN(n_0_0_135));
   NOR2_X1 i_0_0_386 (.A1(rst), .A2(n_0_0_136), .ZN(n_0_413));
   AOI222_X1 i_0_0_387 (.A1(A_r[27]), .A2(n_0_0_144), .B1(a[27]), .B2(n_0_0_140), 
      .C1(n_0_27), .C2(n_0_0_142), .ZN(n_0_0_136));
   NOR2_X1 i_0_0_388 (.A1(rst), .A2(n_0_0_137), .ZN(n_0_414));
   AOI222_X1 i_0_0_389 (.A1(A_r[28]), .A2(n_0_0_144), .B1(a[28]), .B2(n_0_0_140), 
      .C1(n_0_28), .C2(n_0_0_142), .ZN(n_0_0_137));
   NOR2_X1 i_0_0_390 (.A1(rst), .A2(n_0_0_138), .ZN(n_0_415));
   AOI222_X1 i_0_0_391 (.A1(A_r[29]), .A2(n_0_0_144), .B1(a[29]), .B2(n_0_0_140), 
      .C1(n_0_29), .C2(n_0_0_142), .ZN(n_0_0_138));
   NOR2_X1 i_0_0_392 (.A1(rst), .A2(n_0_0_139), .ZN(n_0_416));
   AOI222_X1 i_0_0_393 (.A1(A_r[30]), .A2(n_0_0_144), .B1(a[30]), .B2(n_0_0_140), 
      .C1(n_0_30), .C2(n_0_0_142), .ZN(n_0_0_139));
   NOR2_X1 i_0_0_394 (.A1(a[31]), .A2(n_0_0_144), .ZN(n_0_0_140));
   NOR2_X1 i_0_0_395 (.A1(rst), .A2(n_0_0_141), .ZN(n_0_417));
   AOI22_X1 i_0_0_396 (.A1(A_r[31]), .A2(n_0_0_144), .B1(n_0_31), .B2(n_0_0_142), 
      .ZN(n_0_0_141));
   NOR2_X1 i_0_0_397 (.A1(n_0_0_155), .A2(n_0_0_144), .ZN(n_0_0_142));
   INV_X1 i_0_0_398 (.A(n_0_0_144), .ZN(n_0_0_143));
   NOR4_X1 i_0_0_400 (.A1(counter[6]), .A2(counter[5]), .A3(counter[4]), 
      .A4(counter[3]), .ZN(n_0_0_145));
   NOR3_X1 i_0_0_401 (.A1(counter[2]), .A2(counter[1]), .A3(counter[0]), 
      .ZN(n_0_0_146));
   INV_X1 i_0_0_402 (.A(n_0_418), .ZN(n_0_0_147));
   NAND2_X1 i_0_0_403 (.A1(n_0_0_157), .A2(n_0_0_148), .ZN(n_0_418));
   INV_X1 i_0_0_404 (.A(n_0_0_149), .ZN(n_0_0_148));
   NOR4_X1 i_0_0_405 (.A1(counter[6]), .A2(counter[5]), .A3(n_0_0_150), .A4(
      n_0_0_151), .ZN(n_0_0_149));
   NAND2_X1 i_0_0_406 (.A1(counter[4]), .A2(counter[3]), .ZN(n_0_0_150));
   NAND3_X1 i_0_0_407 (.A1(counter[2]), .A2(counter[1]), .A3(counter[0]), 
      .ZN(n_0_0_151));
   INV_X1 i_0_0_408 (.A(n_0_0_4), .ZN(n_0_0_152));
   INV_X1 i_0_0_409 (.A(negative), .ZN(n_0_0_153));
   INV_X1 i_0_0_410 (.A(b[31]), .ZN(n_0_0_154));
   INV_X1 i_0_0_411 (.A(a[31]), .ZN(n_0_0_155));
   INV_X1 i_0_0_412 (.A(counter[6]), .ZN(n_0_0_156));
   NAND2_X1 i_0_0_132 (.A1(n_0_0_71), .A2(n_0_0_70), .ZN(n_0_226));
   NAND2_X1 i_0_0_133 (.A1(n_0_93), .A2(n_0_0_73), .ZN(n_0_0_70));
   NAND2_X1 i_0_0_134 (.A1(n_0_155), .A2(n_0_0_74), .ZN(n_0_0_71));
   INV_X1 i_0_0_135 (.A(n_0_0_82), .ZN(n_0_361));
   AND2_X1 i_0_0_136 (.A1(n_0_0_158), .A2(n_0_0_72), .ZN(n_0_0_82));
   AOI22_X1 i_0_0_137 (.A1(n_0_0_106), .A2(b[7]), .B1(B_r[7]), .B2(n_0_0_144), 
      .ZN(n_0_0_72));
   NAND2_X1 i_0_0_138 (.A1(n_0_38), .A2(n_0_0_108), .ZN(n_0_0_158));
   INV_X1 i_0_0_140 (.A(n_0_0_83), .ZN(n_0_362));
   AND2_X1 i_0_0_270 (.A1(n_0_0_160), .A2(n_0_0_159), .ZN(n_0_0_83));
   AOI22_X1 i_0_0_271 (.A1(n_0_0_106), .A2(b[8]), .B1(B_r[8]), .B2(n_0_0_144), 
      .ZN(n_0_0_159));
   NAND2_X1 i_0_0_280 (.A1(n_0_39), .A2(n_0_0_108), .ZN(n_0_0_160));
   INV_X1 i_0_0_281 (.A(n_0_0_84), .ZN(n_0_363));
   AND2_X1 i_0_0_282 (.A1(n_0_0_162), .A2(n_0_0_161), .ZN(n_0_0_84));
   AOI22_X1 i_0_0_283 (.A1(n_0_0_106), .A2(b[9]), .B1(B_r[9]), .B2(n_0_0_144), 
      .ZN(n_0_0_161));
   NAND2_X1 i_0_0_284 (.A1(n_0_40), .A2(n_0_0_108), .ZN(n_0_0_162));
   INV_X1 i_0_0_285 (.A(n_0_0_85), .ZN(n_0_364));
   AND2_X1 i_0_0_286 (.A1(n_0_0_164), .A2(n_0_0_163), .ZN(n_0_0_85));
   AOI22_X1 i_0_0_287 (.A1(n_0_0_106), .A2(b[10]), .B1(B_r[10]), .B2(n_0_0_144), 
      .ZN(n_0_0_163));
   NAND2_X1 i_0_0_288 (.A1(n_0_41), .A2(n_0_0_108), .ZN(n_0_0_164));
   INV_X1 i_0_0_289 (.A(n_0_0_86), .ZN(n_0_365));
   AND2_X1 i_0_0_290 (.A1(n_0_0_166), .A2(n_0_0_165), .ZN(n_0_0_86));
   AOI22_X1 i_0_0_291 (.A1(n_0_0_106), .A2(b[11]), .B1(B_r[11]), .B2(n_0_0_144), 
      .ZN(n_0_0_165));
   NAND2_X1 i_0_0_328 (.A1(n_0_42), .A2(n_0_0_108), .ZN(n_0_0_166));
   INV_X1 i_0_0_331 (.A(n_0_0_87), .ZN(n_0_366));
   AND2_X1 i_0_0_399 (.A1(n_0_0_168), .A2(n_0_0_167), .ZN(n_0_0_87));
   AOI22_X1 i_0_0_413 (.A1(n_0_0_106), .A2(b[12]), .B1(B_r[12]), .B2(n_0_0_144), 
      .ZN(n_0_0_167));
   NAND2_X1 i_0_0_414 (.A1(n_0_43), .A2(n_0_0_108), .ZN(n_0_0_168));
   INV_X1 i_0_0_415 (.A(rst), .ZN(n_0_0_157));
   NAND2_X1 i_0_0_416 (.A1(n_0_0_170), .A2(n_0_0_169), .ZN(n_0_225));
   NAND2_X1 i_0_0_417 (.A1(n_0_92), .A2(n_0_0_73), .ZN(n_0_0_169));
   NAND2_X1 i_0_0_418 (.A1(n_0_154), .A2(n_0_0_74), .ZN(n_0_0_170));
   NAND2_X1 i_0_0_419 (.A1(n_0_0_172), .A2(n_0_0_171), .ZN(n_0_227));
   NAND2_X1 i_0_0_420 (.A1(n_0_94), .A2(n_0_0_73), .ZN(n_0_0_171));
   AOI21_X1 i_0_0_421 (.A(rst), .B1(n_0_0_149), .B2(negative), .ZN(n_0_0_73));
   NAND2_X1 i_0_0_422 (.A1(n_0_156), .A2(n_0_0_74), .ZN(n_0_0_172));
   NOR3_X1 i_0_0_423 (.A1(n_0_0_148), .A2(rst), .A3(n_0_0_153), .ZN(n_0_0_74));
   INV_X1 i_0_0_424 (.A(n_0_0_77), .ZN(n_0_356));
   AND2_X1 i_0_0_425 (.A1(n_0_0_174), .A2(n_0_0_173), .ZN(n_0_0_77));
   AOI22_X1 i_0_0_426 (.A1(n_0_0_106), .A2(b[2]), .B1(B_r[2]), .B2(n_0_0_144), 
      .ZN(n_0_0_173));
   NOR2_X1 i_0_0_427 (.A1(b[31]), .A2(n_0_0_144), .ZN(n_0_0_106));
   NAND2_X1 i_0_0_428 (.A1(n_0_33), .A2(n_0_0_108), .ZN(n_0_0_174));
   NOR2_X1 i_0_0_429 (.A1(n_0_0_154), .A2(n_0_0_144), .ZN(n_0_0_108));
   NAND2_X1 i_0_0_430 (.A1(n_0_0_145), .A2(n_0_0_146), .ZN(n_0_0_144));
   DFF_X1 \counter_reg[6]  (.D(n_0_164), .CK(clk), .Q(counter[6]), .QN());
   DFF_X1 \counter_reg[5]  (.D(n_0_163), .CK(clk), .Q(counter[5]), .QN());
   DFF_X1 \counter_reg[4]  (.D(n_0_162), .CK(clk), .Q(counter[4]), .QN());
   DFF_X1 \counter_reg[3]  (.D(n_0_161), .CK(clk), .Q(counter[3]), .QN());
   DFF_X1 \counter_reg[2]  (.D(n_0_160), .CK(clk), .Q(counter[2]), .QN());
   DFF_X1 \counter_reg[1]  (.D(n_0_159), .CK(clk), .Q(counter[1]), .QN());
   DFF_X1 \counter_reg[0]  (.D(n_0_158), .CK(clk), .Q(counter[0]), .QN());
   DFF_X1 \A_r_reg[31]  (.D(n_0_417), .CK(clk), .Q(A_r[31]), .QN());
   DFF_X1 \A_r_reg[30]  (.D(n_0_416), .CK(clk), .Q(A_r[30]), .QN());
   DFF_X1 \A_r_reg[29]  (.D(n_0_415), .CK(clk), .Q(A_r[29]), .QN());
   DFF_X1 \A_r_reg[28]  (.D(n_0_414), .CK(clk), .Q(A_r[28]), .QN());
   DFF_X1 \A_r_reg[27]  (.D(n_0_413), .CK(clk), .Q(A_r[27]), .QN());
   DFF_X1 \A_r_reg[26]  (.D(n_0_412), .CK(clk), .Q(A_r[26]), .QN());
   DFF_X1 \A_r_reg[25]  (.D(n_0_411), .CK(clk), .Q(A_r[25]), .QN());
   DFF_X1 \A_r_reg[24]  (.D(n_0_410), .CK(clk), .Q(A_r[24]), .QN());
   DFF_X1 \A_r_reg[23]  (.D(n_0_409), .CK(clk), .Q(A_r[23]), .QN());
   DFF_X1 \A_r_reg[22]  (.D(n_0_408), .CK(clk), .Q(A_r[22]), .QN());
   DFF_X1 \A_r_reg[21]  (.D(n_0_407), .CK(clk), .Q(A_r[21]), .QN());
   DFF_X1 \A_r_reg[20]  (.D(n_0_406), .CK(clk), .Q(A_r[20]), .QN());
   DFF_X1 \A_r_reg[19]  (.D(n_0_405), .CK(clk), .Q(A_r[19]), .QN());
   DFF_X1 \A_r_reg[18]  (.D(n_0_404), .CK(clk), .Q(A_r[18]), .QN());
   DFF_X1 \A_r_reg[17]  (.D(n_0_403), .CK(clk), .Q(A_r[17]), .QN());
   DFF_X1 \A_r_reg[16]  (.D(n_0_402), .CK(clk), .Q(A_r[16]), .QN());
   DFF_X1 \A_r_reg[15]  (.D(n_0_401), .CK(clk), .Q(A_r[15]), .QN());
   DFF_X1 \A_r_reg[14]  (.D(n_0_400), .CK(clk), .Q(A_r[14]), .QN());
   DFF_X1 \A_r_reg[13]  (.D(n_0_399), .CK(clk), .Q(A_r[13]), .QN());
   DFF_X1 \A_r_reg[12]  (.D(n_0_398), .CK(clk), .Q(A_r[12]), .QN());
   DFF_X1 \A_r_reg[11]  (.D(n_0_397), .CK(clk), .Q(A_r[11]), .QN());
   DFF_X1 \A_r_reg[10]  (.D(n_0_396), .CK(clk), .Q(A_r[10]), .QN());
   DFF_X1 \A_r_reg[9]  (.D(n_0_395), .CK(clk), .Q(A_r[9]), .QN());
   DFF_X1 \A_r_reg[8]  (.D(n_0_394), .CK(clk), .Q(A_r[8]), .QN());
   DFF_X1 \A_r_reg[7]  (.D(n_0_393), .CK(clk), .Q(A_r[7]), .QN());
   DFF_X1 \A_r_reg[6]  (.D(n_0_392), .CK(clk), .Q(A_r[6]), .QN());
   DFF_X1 \A_r_reg[5]  (.D(n_0_391), .CK(clk), .Q(A_r[5]), .QN());
   DFF_X1 \A_r_reg[4]  (.D(n_0_390), .CK(clk), .Q(A_r[4]), .QN());
   DFF_X1 \A_r_reg[3]  (.D(n_0_389), .CK(clk), .Q(A_r[3]), .QN());
   DFF_X1 \A_r_reg[2]  (.D(n_0_388), .CK(clk), .Q(A_r[2]), .QN());
   DFF_X1 \A_r_reg[1]  (.D(n_0_387), .CK(clk), .Q(A_r[1]), .QN());
   DFF_X1 \A_r_reg[0]  (.D(n_0_386), .CK(clk), .Q(A_r[0]), .QN());
   DFF_X1 \B_r_reg[31]  (.D(n_0_291), .CK(clk), .Q(B_r[31]), .QN());
   DFF_X1 \B_r_reg[30]  (.D(n_0_290), .CK(clk), .Q(B_r[30]), .QN());
   DFF_X1 \B_r_reg[29]  (.D(n_0_289), .CK(clk), .Q(B_r[29]), .QN());
   DFF_X1 \B_r_reg[28]  (.D(n_0_288), .CK(clk), .Q(B_r[28]), .QN());
   DFF_X1 \B_r_reg[27]  (.D(n_0_287), .CK(clk), .Q(B_r[27]), .QN());
   DFF_X1 \B_r_reg[26]  (.D(n_0_286), .CK(clk), .Q(B_r[26]), .QN());
   DFF_X1 \B_r_reg[25]  (.D(n_0_285), .CK(clk), .Q(B_r[25]), .QN());
   DFF_X1 \B_r_reg[24]  (.D(n_0_284), .CK(clk), .Q(B_r[24]), .QN());
   DFF_X1 \B_r_reg[23]  (.D(n_0_283), .CK(clk), .Q(B_r[23]), .QN());
   DFF_X1 \B_r_reg[22]  (.D(n_0_282), .CK(clk), .Q(B_r[22]), .QN());
   DFF_X1 \B_r_reg[21]  (.D(n_0_281), .CK(clk), .Q(B_r[21]), .QN());
   DFF_X1 \B_r_reg[20]  (.D(n_0_280), .CK(clk), .Q(B_r[20]), .QN());
   DFF_X1 \B_r_reg[19]  (.D(n_0_279), .CK(clk), .Q(B_r[19]), .QN());
   DFF_X1 \B_r_reg[18]  (.D(n_0_278), .CK(clk), .Q(B_r[18]), .QN());
   DFF_X1 \B_r_reg[17]  (.D(n_0_277), .CK(clk), .Q(B_r[17]), .QN());
   DFF_X1 \B_r_reg[16]  (.D(n_0_276), .CK(clk), .Q(B_r[16]), .QN());
   DFF_X1 \B_r_reg[15]  (.D(n_0_275), .CK(clk), .Q(B_r[15]), .QN());
   DFF_X1 \B_r_reg[14]  (.D(n_0_274), .CK(clk), .Q(B_r[14]), .QN());
   DFF_X1 \B_r_reg[13]  (.D(n_0_273), .CK(clk), .Q(B_r[13]), .QN());
   DFF_X1 \B_r_reg[12]  (.D(n_0_272), .CK(clk), .Q(B_r[12]), .QN());
   DFF_X1 \B_r_reg[11]  (.D(n_0_271), .CK(clk), .Q(B_r[11]), .QN());
   DFF_X1 \B_r_reg[10]  (.D(n_0_270), .CK(clk), .Q(B_r[10]), .QN());
   DFF_X1 \B_r_reg[9]  (.D(n_0_269), .CK(clk), .Q(B_r[9]), .QN());
   DFF_X1 \B_r_reg[8]  (.D(n_0_268), .CK(clk), .Q(B_r[8]), .QN());
   DFF_X1 \B_r_reg[7]  (.D(n_0_267), .CK(clk), .Q(B_r[7]), .QN());
   DFF_X1 \B_r_reg[6]  (.D(n_0_266), .CK(clk), .Q(B_r[6]), .QN());
   DFF_X1 \B_r_reg[5]  (.D(n_0_265), .CK(clk), .Q(B_r[5]), .QN());
   DFF_X1 \B_r_reg[4]  (.D(n_0_264), .CK(clk), .Q(B_r[4]), .QN());
   DFF_X1 \B_r_reg[3]  (.D(n_0_263), .CK(clk), .Q(B_r[3]), .QN());
   DFF_X1 \B_r_reg[2]  (.D(n_0_262), .CK(clk), .Q(B_r[2]), .QN());
   DFF_X1 \B_r_reg[1]  (.D(n_0_261), .CK(clk), .Q(B_r[1]), .QN());
   DFF_X1 \B_r_reg[0]  (.D(n_0_260), .CK(clk), .Q(B_r[0]), .QN());
   DFF_X1 \Accumulator_reg[30]  (.D(n_0_259), .CK(clk), .Q(Accumulator[30]), 
      .QN());
   DFF_X1 \Accumulator_reg[29]  (.D(n_0_258), .CK(clk), .Q(Accumulator[29]), 
      .QN());
   DFF_X1 \Accumulator_reg[28]  (.D(n_0_257), .CK(clk), .Q(Accumulator[28]), 
      .QN());
   DFF_X1 \Accumulator_reg[27]  (.D(n_0_256), .CK(clk), .Q(Accumulator[27]), 
      .QN());
   DFF_X1 \Accumulator_reg[26]  (.D(n_0_255), .CK(clk), .Q(Accumulator[26]), 
      .QN());
   DFF_X1 \Accumulator_reg[25]  (.D(n_0_254), .CK(clk), .Q(Accumulator[25]), 
      .QN());
   DFF_X1 \Accumulator_reg[24]  (.D(n_0_253), .CK(clk), .Q(Accumulator[24]), 
      .QN());
   DFF_X1 \Accumulator_reg[23]  (.D(n_0_252), .CK(clk), .Q(Accumulator[23]), 
      .QN());
   DFF_X1 \Accumulator_reg[22]  (.D(n_0_251), .CK(clk), .Q(Accumulator[22]), 
      .QN());
   DFF_X1 \Accumulator_reg[21]  (.D(n_0_250), .CK(clk), .Q(Accumulator[21]), 
      .QN());
   DFF_X1 \Accumulator_reg[20]  (.D(n_0_249), .CK(clk), .Q(Accumulator[20]), 
      .QN());
   DFF_X1 \Accumulator_reg[19]  (.D(n_0_248), .CK(clk), .Q(Accumulator[19]), 
      .QN());
   DFF_X1 \Accumulator_reg[18]  (.D(n_0_247), .CK(clk), .Q(Accumulator[18]), 
      .QN());
   DFF_X1 \Accumulator_reg[17]  (.D(n_0_246), .CK(clk), .Q(Accumulator[17]), 
      .QN());
   DFF_X1 \Accumulator_reg[16]  (.D(n_0_245), .CK(clk), .Q(Accumulator[16]), 
      .QN());
   DFF_X1 \Accumulator_reg[15]  (.D(n_0_244), .CK(clk), .Q(Accumulator[15]), 
      .QN());
   DFF_X1 \Accumulator_reg[14]  (.D(n_0_243), .CK(clk), .Q(Accumulator[14]), 
      .QN());
   DFF_X1 \Accumulator_reg[13]  (.D(n_0_242), .CK(clk), .Q(Accumulator[13]), 
      .QN());
   DFF_X1 \Accumulator_reg[12]  (.D(n_0_241), .CK(clk), .Q(Accumulator[12]), 
      .QN());
   DFF_X1 \Accumulator_reg[11]  (.D(n_0_240), .CK(clk), .Q(Accumulator[11]), 
      .QN());
   DFF_X1 \Accumulator_reg[10]  (.D(n_0_239), .CK(clk), .Q(Accumulator[10]), 
      .QN());
   DFF_X1 \Accumulator_reg[9]  (.D(n_0_238), .CK(clk), .Q(Accumulator[9]), .QN());
   DFF_X1 \Accumulator_reg[8]  (.D(n_0_237), .CK(clk), .Q(Accumulator[8]), .QN());
   DFF_X1 \Accumulator_reg[7]  (.D(n_0_236), .CK(clk), .Q(Accumulator[7]), .QN());
   DFF_X1 \Accumulator_reg[6]  (.D(n_0_235), .CK(clk), .Q(Accumulator[6]), .QN());
   DFF_X1 \Accumulator_reg[5]  (.D(n_0_234), .CK(clk), .Q(Accumulator[5]), .QN());
   DFF_X1 \Accumulator_reg[4]  (.D(n_0_233), .CK(clk), .Q(Accumulator[4]), .QN());
   DFF_X1 \Accumulator_reg[3]  (.D(n_0_232), .CK(clk), .Q(Accumulator[3]), .QN());
   DFF_X1 \Accumulator_reg[2]  (.D(n_0_231), .CK(clk), .Q(Accumulator[2]), .QN());
   DFF_X1 \Accumulator_reg[1]  (.D(n_0_230), .CK(clk), .Q(Accumulator[1]), .QN());
   DFF_X1 \Accumulator_reg[0]  (.D(n_0_229), .CK(clk), .Q(Accumulator[0]), .QN());
   DFF_X1 negative_reg (.D(n_0_165), .CK(clk), .Q(negative), .QN());
endmodule
