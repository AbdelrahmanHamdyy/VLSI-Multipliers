/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu Dec 22 23:56:51 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1210537045 */

module buffer__0_68(clk, rst, en, D, Q);
   input clk;
   input rst;
   input en;
   input [31:0]D;
   output [31:0]Q;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[31]  (.D(n_33), .CK(n_0), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_32), .CK(n_0), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_31), .CK(n_0), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_30), .CK(n_0), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_29), .CK(n_0), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_28), .CK(n_0), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_27), .CK(n_0), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_26), .CK(n_0), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_25), .CK(n_0), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_24), .CK(n_0), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_23), .CK(n_0), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_22), .CK(n_0), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_21), .CK(n_0), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_20), .CK(n_0), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_19), .CK(n_0), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_18), .CK(n_0), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_17), .CK(n_0), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_16), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_15), .CK(n_0), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_14), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_13), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_12), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_11), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_10), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_9), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_8), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_7), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_6), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_5), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_4), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_3), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_2), .CK(n_0), .Q(Q[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(rst), .ZN(n_1));
   INV_X1 i_0_1 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(D[31]), .ZN(n_33));
endmodule

module buffer(clk, rst, en, D, Q);
   input clk;
   input rst;
   input en;
   input [31:0]D;
   output [31:0]Q;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[31]  (.D(n_33), .CK(n_0), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_32), .CK(n_0), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_31), .CK(n_0), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_30), .CK(n_0), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_29), .CK(n_0), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_28), .CK(n_0), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_27), .CK(n_0), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_26), .CK(n_0), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_25), .CK(n_0), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_24), .CK(n_0), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_23), .CK(n_0), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_22), .CK(n_0), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_21), .CK(n_0), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_20), .CK(n_0), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_19), .CK(n_0), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_18), .CK(n_0), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_17), .CK(n_0), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_16), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_15), .CK(n_0), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_14), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_13), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_12), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_11), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_10), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_9), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_8), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_7), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_6), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_5), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_4), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_3), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_2), .CK(n_0), .Q(Q[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(rst), .ZN(n_1));
   INV_X1 i_0_1 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(D[31]), .ZN(n_33));
endmodule

module datapath(b, a, p_0);
   input [31:0]b;
   input [31:0]a;
   output [63:0]p_0;

   HA_X1 i_0 (.A(n_2818), .B(n_3231), .CO(n_1), .S(n_0));
   FA_X1 i_1 (.A(n_2786), .B(n_2817), .CI(n_2848), .CO(n_3), .S(n_2));
   HA_X1 i_2 (.A(n_2877), .B(n_1), .CO(n_5), .S(n_4));
   FA_X1 i_3 (.A(n_2754), .B(n_2785), .CI(n_2816), .CO(n_7), .S(n_6));
   FA_X1 i_4 (.A(n_2847), .B(n_2876), .CI(n_5), .CO(n_9), .S(n_8));
   HA_X1 i_5 (.A(n_3), .B(n_8), .CO(n_11), .S(n_10));
   FA_X1 i_6 (.A(n_2722), .B(n_2753), .CI(n_2784), .CO(n_13), .S(n_12));
   FA_X1 i_7 (.A(n_2815), .B(n_2846), .CI(n_2875), .CO(n_15), .S(n_14));
   FA_X1 i_8 (.A(n_7), .B(n_9), .CI(n_14), .CO(n_17), .S(n_16));
   HA_X1 i_9 (.A(n_12), .B(n_11), .CO(n_19), .S(n_18));
   FA_X1 i_10 (.A(n_2690), .B(n_2721), .CI(n_2752), .CO(n_21), .S(n_20));
   FA_X1 i_11 (.A(n_2783), .B(n_2814), .CI(n_2845), .CO(n_23), .S(n_22));
   FA_X1 i_12 (.A(n_2874), .B(n_15), .CI(n_13), .CO(n_25), .S(n_24));
   FA_X1 i_13 (.A(n_22), .B(n_20), .CI(n_24), .CO(n_27), .S(n_26));
   HA_X1 i_14 (.A(n_19), .B(n_17), .CO(n_29), .S(n_28));
   FA_X1 i_15 (.A(n_2658), .B(n_2689), .CI(n_2720), .CO(n_31), .S(n_30));
   FA_X1 i_16 (.A(n_2751), .B(n_2782), .CI(n_2813), .CO(n_33), .S(n_32));
   FA_X1 i_17 (.A(n_2844), .B(n_2873), .CI(n_23), .CO(n_35), .S(n_34));
   FA_X1 i_18 (.A(n_21), .B(n_25), .CI(n_34), .CO(n_37), .S(n_36));
   FA_X1 i_19 (.A(n_32), .B(n_30), .CI(n_29), .CO(n_39), .S(n_38));
   HA_X1 i_20 (.A(n_36), .B(n_27), .CO(n_41), .S(n_40));
   FA_X1 i_21 (.A(n_2626), .B(n_2657), .CI(n_2688), .CO(n_43), .S(n_42));
   FA_X1 i_22 (.A(n_2719), .B(n_2750), .CI(n_2781), .CO(n_45), .S(n_44));
   FA_X1 i_23 (.A(n_2812), .B(n_2843), .CI(n_2872), .CO(n_47), .S(n_46));
   FA_X1 i_24 (.A(n_33), .B(n_31), .CI(n_35), .CO(n_49), .S(n_48));
   FA_X1 i_25 (.A(n_46), .B(n_44), .CI(n_42), .CO(n_51), .S(n_50));
   FA_X1 i_26 (.A(n_48), .B(n_37), .CI(n_41), .CO(n_53), .S(n_52));
   HA_X1 i_27 (.A(n_39), .B(n_50), .CO(n_55), .S(n_54));
   FA_X1 i_28 (.A(n_2594), .B(n_2625), .CI(n_2656), .CO(n_57), .S(n_56));
   FA_X1 i_29 (.A(n_2687), .B(n_2718), .CI(n_2749), .CO(n_59), .S(n_58));
   FA_X1 i_30 (.A(n_2780), .B(n_2811), .CI(n_2842), .CO(n_61), .S(n_60));
   FA_X1 i_31 (.A(n_2871), .B(n_47), .CI(n_45), .CO(n_63), .S(n_62));
   FA_X1 i_32 (.A(n_43), .B(n_60), .CI(n_58), .CO(n_65), .S(n_64));
   FA_X1 i_33 (.A(n_56), .B(n_49), .CI(n_62), .CO(n_67), .S(n_66));
   FA_X1 i_34 (.A(n_51), .B(n_64), .CI(n_66), .CO(n_69), .S(n_68));
   HA_X1 i_35 (.A(n_55), .B(n_53), .CO(n_71), .S(n_70));
   FA_X1 i_36 (.A(n_2562), .B(n_2593), .CI(n_2624), .CO(n_73), .S(n_72));
   FA_X1 i_37 (.A(n_2655), .B(n_2686), .CI(n_2717), .CO(n_75), .S(n_74));
   FA_X1 i_38 (.A(n_2748), .B(n_2779), .CI(n_2810), .CO(n_77), .S(n_76));
   FA_X1 i_39 (.A(n_2841), .B(n_2870), .CI(n_61), .CO(n_79), .S(n_78));
   FA_X1 i_40 (.A(n_59), .B(n_57), .CI(n_63), .CO(n_81), .S(n_80));
   FA_X1 i_41 (.A(n_78), .B(n_76), .CI(n_74), .CO(n_83), .S(n_82));
   FA_X1 i_42 (.A(n_72), .B(n_80), .CI(n_65), .CO(n_85), .S(n_84));
   FA_X1 i_43 (.A(n_67), .B(n_82), .CI(n_84), .CO(n_87), .S(n_86));
   HA_X1 i_44 (.A(n_71), .B(n_69), .CO(n_89), .S(n_88));
   FA_X1 i_45 (.A(n_2530), .B(n_2561), .CI(n_2592), .CO(n_91), .S(n_90));
   FA_X1 i_46 (.A(n_2623), .B(n_2654), .CI(n_2685), .CO(n_93), .S(n_92));
   FA_X1 i_47 (.A(n_2716), .B(n_2747), .CI(n_2778), .CO(n_95), .S(n_94));
   FA_X1 i_48 (.A(n_2809), .B(n_2840), .CI(n_2869), .CO(n_97), .S(n_96));
   FA_X1 i_49 (.A(n_77), .B(n_75), .CI(n_73), .CO(n_99), .S(n_98));
   FA_X1 i_50 (.A(n_79), .B(n_96), .CI(n_94), .CO(n_101), .S(n_100));
   FA_X1 i_51 (.A(n_92), .B(n_90), .CI(n_81), .CO(n_103), .S(n_102));
   FA_X1 i_52 (.A(n_98), .B(n_83), .CI(n_85), .CO(n_105), .S(n_104));
   FA_X1 i_53 (.A(n_102), .B(n_100), .CI(n_104), .CO(n_107), .S(n_106));
   HA_X1 i_54 (.A(n_89), .B(n_87), .CO(n_109), .S(n_108));
   FA_X1 i_55 (.A(n_2498), .B(n_2529), .CI(n_2560), .CO(n_111), .S(n_110));
   FA_X1 i_56 (.A(n_2591), .B(n_2622), .CI(n_2653), .CO(n_113), .S(n_112));
   FA_X1 i_57 (.A(n_2684), .B(n_2715), .CI(n_2746), .CO(n_115), .S(n_114));
   FA_X1 i_58 (.A(n_2777), .B(n_2808), .CI(n_2839), .CO(n_117), .S(n_116));
   FA_X1 i_59 (.A(n_2868), .B(n_97), .CI(n_95), .CO(n_119), .S(n_118));
   FA_X1 i_60 (.A(n_93), .B(n_91), .CI(n_99), .CO(n_121), .S(n_120));
   FA_X1 i_61 (.A(n_116), .B(n_114), .CI(n_112), .CO(n_123), .S(n_122));
   FA_X1 i_62 (.A(n_110), .B(n_120), .CI(n_118), .CO(n_125), .S(n_124));
   FA_X1 i_63 (.A(n_101), .B(n_103), .CI(n_122), .CO(n_127), .S(n_126));
   FA_X1 i_64 (.A(n_105), .B(n_124), .CI(n_126), .CO(n_129), .S(n_128));
   HA_X1 i_65 (.A(n_107), .B(n_109), .CO(n_131), .S(n_130));
   FA_X1 i_66 (.A(n_2466), .B(n_2497), .CI(n_2528), .CO(n_133), .S(n_132));
   FA_X1 i_67 (.A(n_2559), .B(n_2590), .CI(n_2621), .CO(n_135), .S(n_134));
   FA_X1 i_68 (.A(n_2652), .B(n_2683), .CI(n_2714), .CO(n_137), .S(n_136));
   FA_X1 i_69 (.A(n_2745), .B(n_2776), .CI(n_2807), .CO(n_139), .S(n_138));
   FA_X1 i_70 (.A(n_2838), .B(n_2867), .CI(n_117), .CO(n_141), .S(n_140));
   FA_X1 i_71 (.A(n_115), .B(n_113), .CI(n_111), .CO(n_143), .S(n_142));
   FA_X1 i_72 (.A(n_119), .B(n_140), .CI(n_138), .CO(n_145), .S(n_144));
   FA_X1 i_73 (.A(n_136), .B(n_134), .CI(n_132), .CO(n_147), .S(n_146));
   FA_X1 i_74 (.A(n_121), .B(n_142), .CI(n_123), .CO(n_149), .S(n_148));
   FA_X1 i_75 (.A(n_125), .B(n_146), .CI(n_144), .CO(n_151), .S(n_150));
   FA_X1 i_76 (.A(n_148), .B(n_127), .CI(n_129), .CO(n_153), .S(n_152));
   HA_X1 i_77 (.A(n_150), .B(n_131), .CO(n_155), .S(n_154));
   FA_X1 i_78 (.A(n_2434), .B(n_2465), .CI(n_2496), .CO(n_157), .S(n_156));
   FA_X1 i_79 (.A(n_2527), .B(n_2558), .CI(n_2589), .CO(n_159), .S(n_158));
   FA_X1 i_80 (.A(n_2620), .B(n_2651), .CI(n_2682), .CO(n_161), .S(n_160));
   FA_X1 i_81 (.A(n_2713), .B(n_2744), .CI(n_2775), .CO(n_163), .S(n_162));
   FA_X1 i_82 (.A(n_2806), .B(n_2837), .CI(n_2866), .CO(n_165), .S(n_164));
   FA_X1 i_83 (.A(n_139), .B(n_137), .CI(n_135), .CO(n_167), .S(n_166));
   FA_X1 i_84 (.A(n_133), .B(n_143), .CI(n_141), .CO(n_169), .S(n_168));
   FA_X1 i_85 (.A(n_164), .B(n_162), .CI(n_160), .CO(n_171), .S(n_170));
   FA_X1 i_86 (.A(n_158), .B(n_156), .CI(n_166), .CO(n_173), .S(n_172));
   FA_X1 i_87 (.A(n_147), .B(n_145), .CI(n_168), .CO(n_175), .S(n_174));
   FA_X1 i_88 (.A(n_149), .B(n_172), .CI(n_170), .CO(n_177), .S(n_176));
   FA_X1 i_89 (.A(n_174), .B(n_151), .CI(n_176), .CO(n_179), .S(n_178));
   HA_X1 i_90 (.A(n_153), .B(n_155), .CO(n_181), .S(n_180));
   FA_X1 i_91 (.A(n_2402), .B(n_2433), .CI(n_2464), .CO(n_183), .S(n_182));
   FA_X1 i_92 (.A(n_2495), .B(n_2526), .CI(n_2557), .CO(n_185), .S(n_184));
   FA_X1 i_93 (.A(n_2588), .B(n_2619), .CI(n_2650), .CO(n_187), .S(n_186));
   FA_X1 i_94 (.A(n_2681), .B(n_2712), .CI(n_2743), .CO(n_189), .S(n_188));
   FA_X1 i_95 (.A(n_2774), .B(n_2805), .CI(n_2836), .CO(n_191), .S(n_190));
   FA_X1 i_96 (.A(n_2865), .B(n_165), .CI(n_163), .CO(n_193), .S(n_192));
   FA_X1 i_97 (.A(n_161), .B(n_159), .CI(n_157), .CO(n_195), .S(n_194));
   FA_X1 i_98 (.A(n_167), .B(n_190), .CI(n_188), .CO(n_197), .S(n_196));
   FA_X1 i_99 (.A(n_186), .B(n_184), .CI(n_182), .CO(n_199), .S(n_198));
   FA_X1 i_100 (.A(n_169), .B(n_194), .CI(n_192), .CO(n_201), .S(n_200));
   FA_X1 i_101 (.A(n_171), .B(n_173), .CI(n_198), .CO(n_203), .S(n_202));
   FA_X1 i_102 (.A(n_196), .B(n_175), .CI(n_200), .CO(n_205), .S(n_204));
   FA_X1 i_103 (.A(n_177), .B(n_202), .CI(n_204), .CO(n_207), .S(n_206));
   HA_X1 i_104 (.A(n_179), .B(n_181), .CO(n_209), .S(n_208));
   FA_X1 i_105 (.A(n_2370), .B(n_2401), .CI(n_2432), .CO(n_211), .S(n_210));
   FA_X1 i_106 (.A(n_2463), .B(n_2494), .CI(n_2525), .CO(n_213), .S(n_212));
   FA_X1 i_107 (.A(n_2556), .B(n_2587), .CI(n_2618), .CO(n_215), .S(n_214));
   FA_X1 i_108 (.A(n_2649), .B(n_2680), .CI(n_2711), .CO(n_217), .S(n_216));
   FA_X1 i_109 (.A(n_2742), .B(n_2773), .CI(n_2804), .CO(n_219), .S(n_218));
   FA_X1 i_110 (.A(n_2835), .B(n_2864), .CI(n_191), .CO(n_221), .S(n_220));
   FA_X1 i_111 (.A(n_189), .B(n_187), .CI(n_185), .CO(n_223), .S(n_222));
   FA_X1 i_112 (.A(n_183), .B(n_195), .CI(n_193), .CO(n_225), .S(n_224));
   FA_X1 i_113 (.A(n_220), .B(n_218), .CI(n_216), .CO(n_227), .S(n_226));
   FA_X1 i_114 (.A(n_214), .B(n_212), .CI(n_210), .CO(n_229), .S(n_228));
   FA_X1 i_115 (.A(n_222), .B(n_199), .CI(n_197), .CO(n_231), .S(n_230));
   FA_X1 i_116 (.A(n_224), .B(n_201), .CI(n_228), .CO(n_233), .S(n_232));
   FA_X1 i_117 (.A(n_226), .B(n_230), .CI(n_203), .CO(n_235), .S(n_234));
   FA_X1 i_118 (.A(n_232), .B(n_205), .CI(n_234), .CO(n_237), .S(n_236));
   HA_X1 i_119 (.A(n_207), .B(n_209), .CO(n_239), .S(n_238));
   FA_X1 i_120 (.A(n_2338), .B(n_2369), .CI(n_2400), .CO(n_241), .S(n_240));
   FA_X1 i_121 (.A(n_2431), .B(n_2462), .CI(n_2493), .CO(n_243), .S(n_242));
   FA_X1 i_122 (.A(n_2524), .B(n_2555), .CI(n_2586), .CO(n_245), .S(n_244));
   FA_X1 i_123 (.A(n_2617), .B(n_2648), .CI(n_2679), .CO(n_247), .S(n_246));
   FA_X1 i_124 (.A(n_2710), .B(n_2741), .CI(n_2772), .CO(n_249), .S(n_248));
   FA_X1 i_125 (.A(n_2803), .B(n_2834), .CI(n_2863), .CO(n_251), .S(n_250));
   FA_X1 i_126 (.A(n_219), .B(n_217), .CI(n_215), .CO(n_253), .S(n_252));
   FA_X1 i_127 (.A(n_213), .B(n_211), .CI(n_223), .CO(n_255), .S(n_254));
   FA_X1 i_128 (.A(n_221), .B(n_250), .CI(n_248), .CO(n_257), .S(n_256));
   FA_X1 i_129 (.A(n_246), .B(n_244), .CI(n_242), .CO(n_259), .S(n_258));
   FA_X1 i_130 (.A(n_240), .B(n_225), .CI(n_254), .CO(n_261), .S(n_260));
   FA_X1 i_131 (.A(n_252), .B(n_229), .CI(n_227), .CO(n_263), .S(n_262));
   FA_X1 i_132 (.A(n_231), .B(n_258), .CI(n_256), .CO(n_265), .S(n_264));
   FA_X1 i_133 (.A(n_260), .B(n_262), .CI(n_233), .CO(n_267), .S(n_266));
   FA_X1 i_134 (.A(n_235), .B(n_264), .CI(n_266), .CO(n_269), .S(n_268));
   HA_X1 i_135 (.A(n_237), .B(n_239), .CO(n_271), .S(n_270));
   FA_X1 i_136 (.A(n_2306), .B(n_2337), .CI(n_2368), .CO(n_273), .S(n_272));
   FA_X1 i_137 (.A(n_2399), .B(n_2430), .CI(n_2461), .CO(n_275), .S(n_274));
   FA_X1 i_138 (.A(n_2492), .B(n_2523), .CI(n_2554), .CO(n_277), .S(n_276));
   FA_X1 i_139 (.A(n_2585), .B(n_2616), .CI(n_2647), .CO(n_279), .S(n_278));
   FA_X1 i_140 (.A(n_2678), .B(n_2709), .CI(n_2740), .CO(n_281), .S(n_280));
   FA_X1 i_141 (.A(n_2771), .B(n_2802), .CI(n_2833), .CO(n_283), .S(n_282));
   FA_X1 i_142 (.A(n_2862), .B(n_251), .CI(n_249), .CO(n_285), .S(n_284));
   FA_X1 i_143 (.A(n_247), .B(n_245), .CI(n_243), .CO(n_287), .S(n_286));
   FA_X1 i_144 (.A(n_241), .B(n_253), .CI(n_282), .CO(n_289), .S(n_288));
   FA_X1 i_145 (.A(n_280), .B(n_278), .CI(n_276), .CO(n_291), .S(n_290));
   FA_X1 i_146 (.A(n_274), .B(n_272), .CI(n_255), .CO(n_293), .S(n_292));
   FA_X1 i_147 (.A(n_286), .B(n_284), .CI(n_259), .CO(n_295), .S(n_294));
   FA_X1 i_148 (.A(n_257), .B(n_288), .CI(n_263), .CO(n_297), .S(n_296));
   FA_X1 i_149 (.A(n_261), .B(n_292), .CI(n_290), .CO(n_299), .S(n_298));
   FA_X1 i_150 (.A(n_294), .B(n_265), .CI(n_296), .CO(n_301), .S(n_300));
   FA_X1 i_151 (.A(n_267), .B(n_298), .CI(n_300), .CO(n_303), .S(n_302));
   HA_X1 i_152 (.A(n_269), .B(n_302), .CO(n_305), .S(n_304));
   FA_X1 i_153 (.A(n_2274), .B(n_2305), .CI(n_2336), .CO(n_307), .S(n_306));
   FA_X1 i_154 (.A(n_2367), .B(n_2398), .CI(n_2429), .CO(n_309), .S(n_308));
   FA_X1 i_155 (.A(n_2460), .B(n_2491), .CI(n_2522), .CO(n_311), .S(n_310));
   FA_X1 i_156 (.A(n_2553), .B(n_2584), .CI(n_2615), .CO(n_313), .S(n_312));
   FA_X1 i_157 (.A(n_2646), .B(n_2677), .CI(n_2708), .CO(n_315), .S(n_314));
   FA_X1 i_158 (.A(n_2739), .B(n_2770), .CI(n_2801), .CO(n_317), .S(n_316));
   FA_X1 i_159 (.A(n_2832), .B(n_2861), .CI(n_283), .CO(n_319), .S(n_318));
   FA_X1 i_160 (.A(n_281), .B(n_279), .CI(n_277), .CO(n_321), .S(n_320));
   FA_X1 i_161 (.A(n_275), .B(n_273), .CI(n_287), .CO(n_323), .S(n_322));
   FA_X1 i_162 (.A(n_285), .B(n_318), .CI(n_316), .CO(n_325), .S(n_324));
   FA_X1 i_163 (.A(n_314), .B(n_312), .CI(n_310), .CO(n_327), .S(n_326));
   FA_X1 i_164 (.A(n_308), .B(n_306), .CI(n_322), .CO(n_329), .S(n_328));
   FA_X1 i_165 (.A(n_320), .B(n_291), .CI(n_289), .CO(n_331), .S(n_330));
   FA_X1 i_166 (.A(n_293), .B(n_295), .CI(n_328), .CO(n_333), .S(n_332));
   FA_X1 i_167 (.A(n_326), .B(n_324), .CI(n_297), .CO(n_335), .S(n_334));
   FA_X1 i_168 (.A(n_330), .B(n_299), .CI(n_332), .CO(n_337), .S(n_336));
   FA_X1 i_169 (.A(n_334), .B(n_301), .CI(n_336), .CO(n_339), .S(n_338));
   HA_X1 i_170 (.A(n_303), .B(n_338), .CO(n_341), .S(n_340));
   FA_X1 i_171 (.A(n_2242), .B(n_2273), .CI(n_2304), .CO(n_343), .S(n_342));
   FA_X1 i_172 (.A(n_2335), .B(n_2366), .CI(n_2397), .CO(n_345), .S(n_344));
   FA_X1 i_173 (.A(n_2428), .B(n_2459), .CI(n_2490), .CO(n_347), .S(n_346));
   FA_X1 i_174 (.A(n_2521), .B(n_2552), .CI(n_2583), .CO(n_349), .S(n_348));
   FA_X1 i_175 (.A(n_2614), .B(n_2645), .CI(n_2676), .CO(n_351), .S(n_350));
   FA_X1 i_176 (.A(n_2707), .B(n_2738), .CI(n_2769), .CO(n_353), .S(n_352));
   FA_X1 i_177 (.A(n_2800), .B(n_2831), .CI(n_2860), .CO(n_355), .S(n_354));
   FA_X1 i_178 (.A(n_317), .B(n_315), .CI(n_313), .CO(n_357), .S(n_356));
   FA_X1 i_179 (.A(n_311), .B(n_309), .CI(n_307), .CO(n_359), .S(n_358));
   FA_X1 i_180 (.A(n_321), .B(n_319), .CI(n_354), .CO(n_361), .S(n_360));
   FA_X1 i_181 (.A(n_352), .B(n_350), .CI(n_348), .CO(n_363), .S(n_362));
   FA_X1 i_182 (.A(n_346), .B(n_344), .CI(n_342), .CO(n_365), .S(n_364));
   FA_X1 i_183 (.A(n_323), .B(n_358), .CI(n_356), .CO(n_367), .S(n_366));
   FA_X1 i_184 (.A(n_327), .B(n_325), .CI(n_360), .CO(n_369), .S(n_368));
   FA_X1 i_185 (.A(n_331), .B(n_329), .CI(n_364), .CO(n_371), .S(n_370));
   FA_X1 i_186 (.A(n_362), .B(n_368), .CI(n_366), .CO(n_373), .S(n_372));
   FA_X1 i_187 (.A(n_333), .B(n_335), .CI(n_370), .CO(n_375), .S(n_374));
   FA_X1 i_188 (.A(n_337), .B(n_372), .CI(n_374), .CO(n_377), .S(n_376));
   HA_X1 i_189 (.A(n_339), .B(n_341), .CO(n_379), .S(n_378));
   FA_X1 i_190 (.A(n_2210), .B(n_2241), .CI(n_2272), .CO(n_381), .S(n_380));
   FA_X1 i_191 (.A(n_2303), .B(n_2334), .CI(n_2365), .CO(n_383), .S(n_382));
   FA_X1 i_192 (.A(n_2396), .B(n_2427), .CI(n_2458), .CO(n_385), .S(n_384));
   FA_X1 i_193 (.A(n_2489), .B(n_2520), .CI(n_2551), .CO(n_387), .S(n_386));
   FA_X1 i_194 (.A(n_2582), .B(n_2613), .CI(n_2644), .CO(n_389), .S(n_388));
   FA_X1 i_195 (.A(n_2675), .B(n_2706), .CI(n_2737), .CO(n_391), .S(n_390));
   FA_X1 i_196 (.A(n_2768), .B(n_2799), .CI(n_2830), .CO(n_393), .S(n_392));
   FA_X1 i_197 (.A(n_2859), .B(n_355), .CI(n_353), .CO(n_395), .S(n_394));
   FA_X1 i_198 (.A(n_351), .B(n_349), .CI(n_347), .CO(n_397), .S(n_396));
   FA_X1 i_199 (.A(n_345), .B(n_343), .CI(n_359), .CO(n_399), .S(n_398));
   FA_X1 i_200 (.A(n_357), .B(n_392), .CI(n_390), .CO(n_401), .S(n_400));
   FA_X1 i_201 (.A(n_388), .B(n_386), .CI(n_384), .CO(n_403), .S(n_402));
   FA_X1 i_202 (.A(n_382), .B(n_380), .CI(n_398), .CO(n_405), .S(n_404));
   FA_X1 i_203 (.A(n_396), .B(n_394), .CI(n_365), .CO(n_407), .S(n_406));
   FA_X1 i_204 (.A(n_363), .B(n_361), .CI(n_367), .CO(n_409), .S(n_408));
   FA_X1 i_205 (.A(n_404), .B(n_402), .CI(n_400), .CO(n_411), .S(n_410));
   FA_X1 i_206 (.A(n_369), .B(n_408), .CI(n_406), .CO(n_413), .S(n_412));
   FA_X1 i_207 (.A(n_371), .B(n_373), .CI(n_410), .CO(n_415), .S(n_414));
   FA_X1 i_208 (.A(n_375), .B(n_412), .CI(n_414), .CO(n_417), .S(n_416));
   HA_X1 i_209 (.A(n_377), .B(n_416), .CO(n_419), .S(n_418));
   FA_X1 i_210 (.A(n_2178), .B(n_2209), .CI(n_2240), .CO(n_421), .S(n_420));
   FA_X1 i_211 (.A(n_2271), .B(n_2302), .CI(n_2333), .CO(n_423), .S(n_422));
   FA_X1 i_212 (.A(n_2364), .B(n_2395), .CI(n_2426), .CO(n_425), .S(n_424));
   FA_X1 i_213 (.A(n_2457), .B(n_2488), .CI(n_2519), .CO(n_427), .S(n_426));
   FA_X1 i_214 (.A(n_2550), .B(n_2581), .CI(n_2612), .CO(n_429), .S(n_428));
   FA_X1 i_215 (.A(n_2643), .B(n_2674), .CI(n_2705), .CO(n_431), .S(n_430));
   FA_X1 i_216 (.A(n_2736), .B(n_2767), .CI(n_2798), .CO(n_433), .S(n_432));
   FA_X1 i_217 (.A(n_2829), .B(n_2858), .CI(n_393), .CO(n_435), .S(n_434));
   FA_X1 i_218 (.A(n_391), .B(n_389), .CI(n_387), .CO(n_437), .S(n_436));
   FA_X1 i_219 (.A(n_385), .B(n_383), .CI(n_381), .CO(n_439), .S(n_438));
   FA_X1 i_220 (.A(n_397), .B(n_395), .CI(n_434), .CO(n_441), .S(n_440));
   FA_X1 i_221 (.A(n_432), .B(n_430), .CI(n_428), .CO(n_443), .S(n_442));
   FA_X1 i_222 (.A(n_426), .B(n_424), .CI(n_422), .CO(n_445), .S(n_444));
   FA_X1 i_223 (.A(n_420), .B(n_399), .CI(n_438), .CO(n_447), .S(n_446));
   FA_X1 i_224 (.A(n_436), .B(n_403), .CI(n_401), .CO(n_449), .S(n_448));
   FA_X1 i_225 (.A(n_440), .B(n_407), .CI(n_405), .CO(n_451), .S(n_450));
   FA_X1 i_226 (.A(n_444), .B(n_442), .CI(n_446), .CO(n_453), .S(n_452));
   FA_X1 i_227 (.A(n_409), .B(n_448), .CI(n_411), .CO(n_455), .S(n_454));
   FA_X1 i_228 (.A(n_450), .B(n_413), .CI(n_452), .CO(n_457), .S(n_456));
   FA_X1 i_229 (.A(n_454), .B(n_415), .CI(n_456), .CO(n_459), .S(n_458));
   HA_X1 i_230 (.A(n_417), .B(n_458), .CO(n_461), .S(n_460));
   FA_X1 i_231 (.A(n_2146), .B(n_2177), .CI(n_2208), .CO(n_463), .S(n_462));
   FA_X1 i_232 (.A(n_2239), .B(n_2270), .CI(n_2301), .CO(n_465), .S(n_464));
   FA_X1 i_233 (.A(n_2332), .B(n_2363), .CI(n_2394), .CO(n_467), .S(n_466));
   FA_X1 i_234 (.A(n_2425), .B(n_2456), .CI(n_2487), .CO(n_469), .S(n_468));
   FA_X1 i_235 (.A(n_2518), .B(n_2549), .CI(n_2580), .CO(n_471), .S(n_470));
   FA_X1 i_236 (.A(n_2611), .B(n_2642), .CI(n_2673), .CO(n_473), .S(n_472));
   FA_X1 i_237 (.A(n_2704), .B(n_2735), .CI(n_2766), .CO(n_475), .S(n_474));
   FA_X1 i_238 (.A(n_2797), .B(n_2828), .CI(n_2857), .CO(n_477), .S(n_476));
   FA_X1 i_239 (.A(n_433), .B(n_431), .CI(n_429), .CO(n_479), .S(n_478));
   FA_X1 i_240 (.A(n_427), .B(n_425), .CI(n_423), .CO(n_481), .S(n_480));
   FA_X1 i_241 (.A(n_421), .B(n_439), .CI(n_437), .CO(n_483), .S(n_482));
   FA_X1 i_242 (.A(n_435), .B(n_476), .CI(n_474), .CO(n_485), .S(n_484));
   FA_X1 i_243 (.A(n_472), .B(n_470), .CI(n_468), .CO(n_487), .S(n_486));
   FA_X1 i_244 (.A(n_466), .B(n_464), .CI(n_462), .CO(n_489), .S(n_488));
   FA_X1 i_245 (.A(n_480), .B(n_478), .CI(n_445), .CO(n_491), .S(n_490));
   FA_X1 i_246 (.A(n_443), .B(n_441), .CI(n_482), .CO(n_493), .S(n_492));
   FA_X1 i_247 (.A(n_449), .B(n_447), .CI(n_488), .CO(n_495), .S(n_494));
   FA_X1 i_248 (.A(n_486), .B(n_484), .CI(n_451), .CO(n_497), .S(n_496));
   FA_X1 i_249 (.A(n_492), .B(n_490), .CI(n_453), .CO(n_499), .S(n_498));
   FA_X1 i_250 (.A(n_494), .B(n_455), .CI(n_496), .CO(n_501), .S(n_500));
   FA_X1 i_251 (.A(n_498), .B(n_457), .CI(n_500), .CO(n_503), .S(n_502));
   HA_X1 i_252 (.A(n_459), .B(n_502), .CO(n_505), .S(n_504));
   FA_X1 i_253 (.A(n_2114), .B(n_2145), .CI(n_2176), .CO(n_507), .S(n_506));
   FA_X1 i_254 (.A(n_2207), .B(n_2238), .CI(n_2269), .CO(n_509), .S(n_508));
   FA_X1 i_255 (.A(n_2300), .B(n_2331), .CI(n_2362), .CO(n_511), .S(n_510));
   FA_X1 i_256 (.A(n_2393), .B(n_2424), .CI(n_2455), .CO(n_513), .S(n_512));
   FA_X1 i_257 (.A(n_2486), .B(n_2517), .CI(n_2548), .CO(n_515), .S(n_514));
   FA_X1 i_258 (.A(n_2579), .B(n_2610), .CI(n_2641), .CO(n_517), .S(n_516));
   FA_X1 i_259 (.A(n_2672), .B(n_2703), .CI(n_2734), .CO(n_519), .S(n_518));
   FA_X1 i_260 (.A(n_2765), .B(n_2796), .CI(n_2827), .CO(n_521), .S(n_520));
   FA_X1 i_261 (.A(n_2856), .B(n_477), .CI(n_475), .CO(n_523), .S(n_522));
   FA_X1 i_262 (.A(n_473), .B(n_471), .CI(n_469), .CO(n_525), .S(n_524));
   FA_X1 i_263 (.A(n_467), .B(n_465), .CI(n_463), .CO(n_527), .S(n_526));
   FA_X1 i_264 (.A(n_481), .B(n_479), .CI(n_520), .CO(n_529), .S(n_528));
   FA_X1 i_265 (.A(n_518), .B(n_516), .CI(n_514), .CO(n_531), .S(n_530));
   FA_X1 i_266 (.A(n_512), .B(n_510), .CI(n_508), .CO(n_533), .S(n_532));
   FA_X1 i_267 (.A(n_506), .B(n_483), .CI(n_526), .CO(n_535), .S(n_534));
   FA_X1 i_268 (.A(n_524), .B(n_522), .CI(n_489), .CO(n_537), .S(n_536));
   FA_X1 i_269 (.A(n_487), .B(n_485), .CI(n_528), .CO(n_539), .S(n_538));
   FA_X1 i_270 (.A(n_491), .B(n_532), .CI(n_530), .CO(n_541), .S(n_540));
   FA_X1 i_271 (.A(n_534), .B(n_493), .CI(n_538), .CO(n_543), .S(n_542));
   FA_X1 i_272 (.A(n_536), .B(n_495), .CI(n_497), .CO(n_545), .S(n_544));
   FA_X1 i_273 (.A(n_499), .B(n_540), .CI(n_542), .CO(n_547), .S(n_546));
   FA_X1 i_274 (.A(n_544), .B(n_501), .CI(n_546), .CO(n_549), .S(n_548));
   HA_X1 i_275 (.A(n_503), .B(n_548), .CO(n_551), .S(n_550));
   FA_X1 i_276 (.A(n_2082), .B(n_2113), .CI(n_2144), .CO(n_553), .S(n_552));
   FA_X1 i_277 (.A(n_2175), .B(n_2206), .CI(n_2237), .CO(n_555), .S(n_554));
   FA_X1 i_278 (.A(n_2268), .B(n_2299), .CI(n_2330), .CO(n_557), .S(n_556));
   FA_X1 i_279 (.A(n_2361), .B(n_2392), .CI(n_2423), .CO(n_559), .S(n_558));
   FA_X1 i_280 (.A(n_2454), .B(n_2485), .CI(n_2516), .CO(n_561), .S(n_560));
   FA_X1 i_281 (.A(n_2547), .B(n_2578), .CI(n_2609), .CO(n_563), .S(n_562));
   FA_X1 i_282 (.A(n_2640), .B(n_2671), .CI(n_2702), .CO(n_565), .S(n_564));
   FA_X1 i_283 (.A(n_2733), .B(n_2764), .CI(n_2795), .CO(n_567), .S(n_566));
   FA_X1 i_284 (.A(n_2826), .B(n_2855), .CI(n_521), .CO(n_569), .S(n_568));
   FA_X1 i_285 (.A(n_519), .B(n_517), .CI(n_515), .CO(n_571), .S(n_570));
   FA_X1 i_286 (.A(n_513), .B(n_511), .CI(n_509), .CO(n_573), .S(n_572));
   FA_X1 i_287 (.A(n_507), .B(n_527), .CI(n_525), .CO(n_575), .S(n_574));
   FA_X1 i_288 (.A(n_523), .B(n_568), .CI(n_566), .CO(n_577), .S(n_576));
   FA_X1 i_289 (.A(n_564), .B(n_562), .CI(n_560), .CO(n_579), .S(n_578));
   FA_X1 i_290 (.A(n_558), .B(n_556), .CI(n_554), .CO(n_581), .S(n_580));
   FA_X1 i_291 (.A(n_552), .B(n_572), .CI(n_570), .CO(n_583), .S(n_582));
   FA_X1 i_292 (.A(n_533), .B(n_531), .CI(n_529), .CO(n_585), .S(n_584));
   FA_X1 i_293 (.A(n_574), .B(n_537), .CI(n_535), .CO(n_587), .S(n_586));
   FA_X1 i_294 (.A(n_580), .B(n_578), .CI(n_576), .CO(n_589), .S(n_588));
   FA_X1 i_295 (.A(n_539), .B(n_584), .CI(n_582), .CO(n_591), .S(n_590));
   FA_X1 i_296 (.A(n_541), .B(n_586), .CI(n_543), .CO(n_593), .S(n_592));
   FA_X1 i_297 (.A(n_545), .B(n_588), .CI(n_590), .CO(n_595), .S(n_594));
   FA_X1 i_298 (.A(n_547), .B(n_592), .CI(n_594), .CO(n_597), .S(n_596));
   HA_X1 i_299 (.A(n_549), .B(n_551), .CO(n_599), .S(n_598));
   FA_X1 i_300 (.A(n_2050), .B(n_2081), .CI(n_2112), .CO(n_601), .S(n_600));
   FA_X1 i_301 (.A(n_2143), .B(n_2174), .CI(n_2205), .CO(n_603), .S(n_602));
   FA_X1 i_302 (.A(n_2236), .B(n_2267), .CI(n_2298), .CO(n_605), .S(n_604));
   FA_X1 i_303 (.A(n_2329), .B(n_2360), .CI(n_2391), .CO(n_607), .S(n_606));
   FA_X1 i_304 (.A(n_2422), .B(n_2453), .CI(n_2484), .CO(n_609), .S(n_608));
   FA_X1 i_305 (.A(n_2515), .B(n_2546), .CI(n_2577), .CO(n_611), .S(n_610));
   FA_X1 i_306 (.A(n_2608), .B(n_2639), .CI(n_2670), .CO(n_613), .S(n_612));
   FA_X1 i_307 (.A(n_2701), .B(n_2732), .CI(n_2763), .CO(n_615), .S(n_614));
   FA_X1 i_308 (.A(n_2794), .B(n_2825), .CI(n_2854), .CO(n_617), .S(n_616));
   FA_X1 i_309 (.A(n_567), .B(n_565), .CI(n_563), .CO(n_619), .S(n_618));
   FA_X1 i_310 (.A(n_561), .B(n_559), .CI(n_557), .CO(n_621), .S(n_620));
   FA_X1 i_311 (.A(n_555), .B(n_553), .CI(n_573), .CO(n_623), .S(n_622));
   FA_X1 i_312 (.A(n_571), .B(n_569), .CI(n_616), .CO(n_625), .S(n_624));
   FA_X1 i_313 (.A(n_614), .B(n_612), .CI(n_610), .CO(n_627), .S(n_626));
   FA_X1 i_314 (.A(n_608), .B(n_606), .CI(n_604), .CO(n_629), .S(n_628));
   FA_X1 i_315 (.A(n_602), .B(n_600), .CI(n_575), .CO(n_631), .S(n_630));
   FA_X1 i_316 (.A(n_622), .B(n_620), .CI(n_618), .CO(n_633), .S(n_632));
   FA_X1 i_317 (.A(n_581), .B(n_579), .CI(n_577), .CO(n_635), .S(n_634));
   FA_X1 i_318 (.A(n_624), .B(n_585), .CI(n_583), .CO(n_637), .S(n_636));
   FA_X1 i_319 (.A(n_630), .B(n_628), .CI(n_626), .CO(n_639), .S(n_638));
   FA_X1 i_320 (.A(n_587), .B(n_634), .CI(n_632), .CO(n_641), .S(n_640));
   FA_X1 i_321 (.A(n_589), .B(n_636), .CI(n_591), .CO(n_643), .S(n_642));
   FA_X1 i_322 (.A(n_638), .B(n_593), .CI(n_640), .CO(n_645), .S(n_644));
   FA_X1 i_323 (.A(n_642), .B(n_595), .CI(n_644), .CO(n_647), .S(n_646));
   HA_X1 i_324 (.A(n_597), .B(n_646), .CO(n_649), .S(n_648));
   FA_X1 i_325 (.A(n_2018), .B(n_2049), .CI(n_2080), .CO(n_651), .S(n_650));
   FA_X1 i_326 (.A(n_2111), .B(n_2142), .CI(n_2173), .CO(n_653), .S(n_652));
   FA_X1 i_327 (.A(n_2204), .B(n_2235), .CI(n_2266), .CO(n_655), .S(n_654));
   FA_X1 i_328 (.A(n_2297), .B(n_2328), .CI(n_2359), .CO(n_657), .S(n_656));
   FA_X1 i_329 (.A(n_2390), .B(n_2421), .CI(n_2452), .CO(n_659), .S(n_658));
   FA_X1 i_330 (.A(n_2483), .B(n_2514), .CI(n_2545), .CO(n_661), .S(n_660));
   FA_X1 i_331 (.A(n_2576), .B(n_2607), .CI(n_2638), .CO(n_663), .S(n_662));
   FA_X1 i_332 (.A(n_2669), .B(n_2700), .CI(n_2731), .CO(n_665), .S(n_664));
   FA_X1 i_333 (.A(n_2762), .B(n_2793), .CI(n_2824), .CO(n_667), .S(n_666));
   FA_X1 i_334 (.A(n_2853), .B(n_617), .CI(n_615), .CO(n_669), .S(n_668));
   FA_X1 i_335 (.A(n_613), .B(n_611), .CI(n_609), .CO(n_671), .S(n_670));
   FA_X1 i_336 (.A(n_607), .B(n_605), .CI(n_603), .CO(n_673), .S(n_672));
   FA_X1 i_337 (.A(n_601), .B(n_621), .CI(n_619), .CO(n_675), .S(n_674));
   FA_X1 i_338 (.A(n_666), .B(n_664), .CI(n_662), .CO(n_677), .S(n_676));
   FA_X1 i_339 (.A(n_660), .B(n_658), .CI(n_656), .CO(n_679), .S(n_678));
   FA_X1 i_340 (.A(n_654), .B(n_652), .CI(n_650), .CO(n_681), .S(n_680));
   FA_X1 i_341 (.A(n_623), .B(n_672), .CI(n_670), .CO(n_683), .S(n_682));
   FA_X1 i_342 (.A(n_668), .B(n_629), .CI(n_627), .CO(n_685), .S(n_684));
   FA_X1 i_343 (.A(n_625), .B(n_631), .CI(n_674), .CO(n_687), .S(n_686));
   FA_X1 i_344 (.A(n_635), .B(n_633), .CI(n_680), .CO(n_689), .S(n_688));
   FA_X1 i_345 (.A(n_678), .B(n_676), .CI(n_637), .CO(n_691), .S(n_690));
   FA_X1 i_346 (.A(n_684), .B(n_682), .CI(n_639), .CO(n_693), .S(n_692));
   FA_X1 i_347 (.A(n_686), .B(n_688), .CI(n_641), .CO(n_695), .S(n_694));
   FA_X1 i_348 (.A(n_690), .B(n_643), .CI(n_692), .CO(n_697), .S(n_696));
   FA_X1 i_349 (.A(n_694), .B(n_645), .CI(n_696), .CO(n_699), .S(n_698));
   HA_X1 i_350 (.A(n_647), .B(n_698), .CO(n_701), .S(n_700));
   FA_X1 i_351 (.A(n_1986), .B(n_2017), .CI(n_2048), .CO(n_703), .S(n_702));
   FA_X1 i_352 (.A(n_2079), .B(n_2110), .CI(n_2141), .CO(n_705), .S(n_704));
   FA_X1 i_353 (.A(n_2172), .B(n_2203), .CI(n_2234), .CO(n_707), .S(n_706));
   FA_X1 i_354 (.A(n_2265), .B(n_2296), .CI(n_2327), .CO(n_709), .S(n_708));
   FA_X1 i_355 (.A(n_2358), .B(n_2389), .CI(n_2420), .CO(n_711), .S(n_710));
   FA_X1 i_356 (.A(n_2451), .B(n_2482), .CI(n_2513), .CO(n_713), .S(n_712));
   FA_X1 i_357 (.A(n_2544), .B(n_2575), .CI(n_2606), .CO(n_715), .S(n_714));
   FA_X1 i_358 (.A(n_2637), .B(n_2668), .CI(n_2699), .CO(n_717), .S(n_716));
   FA_X1 i_359 (.A(n_2730), .B(n_2761), .CI(n_2792), .CO(n_719), .S(n_718));
   FA_X1 i_360 (.A(n_2823), .B(n_2852), .CI(n_667), .CO(n_721), .S(n_720));
   FA_X1 i_361 (.A(n_665), .B(n_663), .CI(n_661), .CO(n_723), .S(n_722));
   FA_X1 i_362 (.A(n_659), .B(n_657), .CI(n_655), .CO(n_725), .S(n_724));
   FA_X1 i_363 (.A(n_653), .B(n_651), .CI(n_673), .CO(n_727), .S(n_726));
   FA_X1 i_364 (.A(n_671), .B(n_669), .CI(n_720), .CO(n_729), .S(n_728));
   FA_X1 i_365 (.A(n_718), .B(n_716), .CI(n_714), .CO(n_731), .S(n_730));
   FA_X1 i_366 (.A(n_712), .B(n_710), .CI(n_708), .CO(n_733), .S(n_732));
   FA_X1 i_367 (.A(n_706), .B(n_704), .CI(n_702), .CO(n_735), .S(n_734));
   FA_X1 i_368 (.A(n_675), .B(n_726), .CI(n_724), .CO(n_737), .S(n_736));
   FA_X1 i_369 (.A(n_722), .B(n_681), .CI(n_679), .CO(n_739), .S(n_738));
   FA_X1 i_370 (.A(n_677), .B(n_728), .CI(n_685), .CO(n_741), .S(n_740));
   FA_X1 i_371 (.A(n_683), .B(n_734), .CI(n_732), .CO(n_743), .S(n_742));
   FA_X1 i_372 (.A(n_730), .B(n_687), .CI(n_738), .CO(n_745), .S(n_744));
   FA_X1 i_373 (.A(n_736), .B(n_689), .CI(n_691), .CO(n_747), .S(n_746));
   FA_X1 i_374 (.A(n_740), .B(n_693), .CI(n_742), .CO(n_749), .S(n_748));
   FA_X1 i_375 (.A(n_744), .B(n_695), .CI(n_746), .CO(n_751), .S(n_750));
   FA_X1 i_376 (.A(n_748), .B(n_697), .CI(n_750), .CO(n_753), .S(n_752));
   HA_X1 i_377 (.A(n_699), .B(n_752), .CO(n_755), .S(n_754));
   FA_X1 i_378 (.A(n_1954), .B(n_1985), .CI(n_2016), .CO(n_757), .S(n_756));
   FA_X1 i_379 (.A(n_2047), .B(n_2078), .CI(n_2109), .CO(n_759), .S(n_758));
   FA_X1 i_380 (.A(n_2140), .B(n_2171), .CI(n_2202), .CO(n_761), .S(n_760));
   FA_X1 i_381 (.A(n_2233), .B(n_2264), .CI(n_2295), .CO(n_763), .S(n_762));
   FA_X1 i_382 (.A(n_2326), .B(n_2357), .CI(n_2388), .CO(n_765), .S(n_764));
   FA_X1 i_383 (.A(n_2419), .B(n_2450), .CI(n_2481), .CO(n_767), .S(n_766));
   FA_X1 i_384 (.A(n_2512), .B(n_2543), .CI(n_2574), .CO(n_769), .S(n_768));
   FA_X1 i_385 (.A(n_2605), .B(n_2636), .CI(n_2667), .CO(n_771), .S(n_770));
   FA_X1 i_386 (.A(n_2698), .B(n_2729), .CI(n_2760), .CO(n_773), .S(n_772));
   FA_X1 i_387 (.A(n_2791), .B(n_2822), .CI(n_2851), .CO(n_775), .S(n_774));
   FA_X1 i_388 (.A(n_719), .B(n_717), .CI(n_715), .CO(n_777), .S(n_776));
   FA_X1 i_389 (.A(n_713), .B(n_711), .CI(n_709), .CO(n_779), .S(n_778));
   FA_X1 i_390 (.A(n_707), .B(n_705), .CI(n_703), .CO(n_781), .S(n_780));
   FA_X1 i_391 (.A(n_725), .B(n_723), .CI(n_721), .CO(n_783), .S(n_782));
   FA_X1 i_392 (.A(n_774), .B(n_772), .CI(n_770), .CO(n_785), .S(n_784));
   FA_X1 i_393 (.A(n_768), .B(n_766), .CI(n_764), .CO(n_787), .S(n_786));
   FA_X1 i_394 (.A(n_762), .B(n_760), .CI(n_758), .CO(n_789), .S(n_788));
   FA_X1 i_395 (.A(n_756), .B(n_727), .CI(n_780), .CO(n_791), .S(n_790));
   FA_X1 i_396 (.A(n_778), .B(n_776), .CI(n_735), .CO(n_793), .S(n_792));
   FA_X1 i_397 (.A(n_733), .B(n_731), .CI(n_729), .CO(n_795), .S(n_794));
   FA_X1 i_398 (.A(n_782), .B(n_739), .CI(n_737), .CO(n_797), .S(n_796));
   FA_X1 i_399 (.A(n_788), .B(n_786), .CI(n_784), .CO(n_799), .S(n_798));
   FA_X1 i_400 (.A(n_790), .B(n_741), .CI(n_794), .CO(n_801), .S(n_800));
   FA_X1 i_401 (.A(n_792), .B(n_743), .CI(n_796), .CO(n_803), .S(n_802));
   FA_X1 i_402 (.A(n_745), .B(n_747), .CI(n_798), .CO(n_805), .S(n_804));
   FA_X1 i_403 (.A(n_800), .B(n_802), .CI(n_749), .CO(n_807), .S(n_806));
   FA_X1 i_404 (.A(n_751), .B(n_804), .CI(n_806), .CO(n_809), .S(n_808));
   HA_X1 i_405 (.A(n_753), .B(n_808), .CO(n_811), .S(n_810));
   FA_X1 i_406 (.A(n_1922), .B(n_1953), .CI(n_1984), .CO(n_813), .S(n_812));
   FA_X1 i_407 (.A(n_2015), .B(n_2046), .CI(n_2077), .CO(n_815), .S(n_814));
   FA_X1 i_408 (.A(n_2108), .B(n_2139), .CI(n_2170), .CO(n_817), .S(n_816));
   FA_X1 i_409 (.A(n_2201), .B(n_2232), .CI(n_2263), .CO(n_819), .S(n_818));
   FA_X1 i_410 (.A(n_2294), .B(n_2325), .CI(n_2356), .CO(n_821), .S(n_820));
   FA_X1 i_411 (.A(n_2387), .B(n_2418), .CI(n_2449), .CO(n_823), .S(n_822));
   FA_X1 i_412 (.A(n_2480), .B(n_2511), .CI(n_2542), .CO(n_825), .S(n_824));
   FA_X1 i_413 (.A(n_2573), .B(n_2604), .CI(n_2635), .CO(n_827), .S(n_826));
   FA_X1 i_414 (.A(n_2666), .B(n_2697), .CI(n_2728), .CO(n_829), .S(n_828));
   FA_X1 i_415 (.A(n_2759), .B(n_2790), .CI(n_2821), .CO(n_831), .S(n_830));
   FA_X1 i_416 (.A(n_2850), .B(n_775), .CI(n_773), .CO(n_833), .S(n_832));
   FA_X1 i_417 (.A(n_771), .B(n_769), .CI(n_767), .CO(n_835), .S(n_834));
   FA_X1 i_418 (.A(n_765), .B(n_763), .CI(n_761), .CO(n_837), .S(n_836));
   FA_X1 i_419 (.A(n_759), .B(n_757), .CI(n_781), .CO(n_839), .S(n_838));
   FA_X1 i_420 (.A(n_779), .B(n_777), .CI(n_830), .CO(n_841), .S(n_840));
   FA_X1 i_421 (.A(n_828), .B(n_826), .CI(n_824), .CO(n_843), .S(n_842));
   FA_X1 i_422 (.A(n_822), .B(n_820), .CI(n_818), .CO(n_845), .S(n_844));
   FA_X1 i_423 (.A(n_816), .B(n_814), .CI(n_812), .CO(n_847), .S(n_846));
   FA_X1 i_424 (.A(n_783), .B(n_838), .CI(n_836), .CO(n_849), .S(n_848));
   FA_X1 i_425 (.A(n_834), .B(n_832), .CI(n_789), .CO(n_851), .S(n_850));
   FA_X1 i_426 (.A(n_787), .B(n_785), .CI(n_840), .CO(n_853), .S(n_852));
   FA_X1 i_427 (.A(n_795), .B(n_793), .CI(n_791), .CO(n_855), .S(n_854));
   FA_X1 i_428 (.A(n_846), .B(n_844), .CI(n_842), .CO(n_857), .S(n_856));
   FA_X1 i_429 (.A(n_797), .B(n_852), .CI(n_850), .CO(n_859), .S(n_858));
   FA_X1 i_430 (.A(n_848), .B(n_799), .CI(n_854), .CO(n_861), .S(n_860));
   FA_X1 i_431 (.A(n_801), .B(n_856), .CI(n_803), .CO(n_863), .S(n_862));
   FA_X1 i_432 (.A(n_860), .B(n_858), .CI(n_805), .CO(n_865), .S(n_864));
   FA_X1 i_433 (.A(n_807), .B(n_862), .CI(n_864), .CO(n_867), .S(n_866));
   HA_X1 i_434 (.A(n_809), .B(n_866), .CO(n_869), .S(n_868));
   FA_X1 i_435 (.A(n_1890), .B(n_1921), .CI(n_1952), .CO(n_871), .S(n_870));
   FA_X1 i_436 (.A(n_1983), .B(n_2014), .CI(n_2045), .CO(n_873), .S(n_872));
   FA_X1 i_437 (.A(n_2076), .B(n_2107), .CI(n_2138), .CO(n_875), .S(n_874));
   FA_X1 i_438 (.A(n_2169), .B(n_2200), .CI(n_2231), .CO(n_877), .S(n_876));
   FA_X1 i_439 (.A(n_2262), .B(n_2293), .CI(n_2324), .CO(n_879), .S(n_878));
   FA_X1 i_440 (.A(n_2355), .B(n_2386), .CI(n_2417), .CO(n_881), .S(n_880));
   FA_X1 i_441 (.A(n_2448), .B(n_2479), .CI(n_2510), .CO(n_883), .S(n_882));
   FA_X1 i_442 (.A(n_2541), .B(n_2572), .CI(n_2603), .CO(n_885), .S(n_884));
   FA_X1 i_443 (.A(n_2634), .B(n_2665), .CI(n_2696), .CO(n_887), .S(n_886));
   FA_X1 i_444 (.A(n_2727), .B(n_2758), .CI(n_2789), .CO(n_889), .S(n_888));
   FA_X1 i_445 (.A(n_2820), .B(n_2849), .CI(n_831), .CO(n_891), .S(n_890));
   FA_X1 i_446 (.A(n_829), .B(n_827), .CI(n_825), .CO(n_893), .S(n_892));
   FA_X1 i_447 (.A(n_823), .B(n_821), .CI(n_819), .CO(n_895), .S(n_894));
   FA_X1 i_448 (.A(n_817), .B(n_815), .CI(n_813), .CO(n_897), .S(n_896));
   FA_X1 i_449 (.A(n_837), .B(n_835), .CI(n_833), .CO(n_899), .S(n_898));
   FA_X1 i_450 (.A(n_890), .B(n_888), .CI(n_886), .CO(n_901), .S(n_900));
   FA_X1 i_451 (.A(n_884), .B(n_882), .CI(n_880), .CO(n_903), .S(n_902));
   FA_X1 i_452 (.A(n_878), .B(n_876), .CI(n_874), .CO(n_905), .S(n_904));
   FA_X1 i_453 (.A(n_872), .B(n_870), .CI(n_839), .CO(n_907), .S(n_906));
   FA_X1 i_454 (.A(n_896), .B(n_894), .CI(n_892), .CO(n_909), .S(n_908));
   FA_X1 i_455 (.A(n_847), .B(n_845), .CI(n_843), .CO(n_911), .S(n_910));
   FA_X1 i_456 (.A(n_841), .B(n_898), .CI(n_851), .CO(n_913), .S(n_912));
   FA_X1 i_457 (.A(n_849), .B(n_906), .CI(n_904), .CO(n_915), .S(n_914));
   FA_X1 i_458 (.A(n_902), .B(n_900), .CI(n_855), .CO(n_917), .S(n_916));
   FA_X1 i_459 (.A(n_853), .B(n_910), .CI(n_908), .CO(n_919), .S(n_918));
   FA_X1 i_460 (.A(n_857), .B(n_912), .CI(n_859), .CO(n_921), .S(n_920));
   FA_X1 i_461 (.A(n_916), .B(n_914), .CI(n_861), .CO(n_923), .S(n_922));
   FA_X1 i_462 (.A(n_918), .B(n_863), .CI(n_920), .CO(n_925), .S(n_924));
   FA_X1 i_463 (.A(n_865), .B(n_922), .CI(n_924), .CO(n_927), .S(n_926));
   HA_X1 i_464 (.A(n_867), .B(n_926), .CO(n_929), .S(n_928));
   FA_X1 i_465 (.A(n_1889), .B(n_1920), .CI(n_1951), .CO(n_931), .S(n_930));
   FA_X1 i_466 (.A(n_1982), .B(n_2013), .CI(n_2044), .CO(n_933), .S(n_932));
   FA_X1 i_467 (.A(n_2075), .B(n_2106), .CI(n_2137), .CO(n_935), .S(n_934));
   FA_X1 i_468 (.A(n_2168), .B(n_2199), .CI(n_2230), .CO(n_937), .S(n_936));
   FA_X1 i_469 (.A(n_2261), .B(n_2292), .CI(n_2323), .CO(n_939), .S(n_938));
   FA_X1 i_470 (.A(n_2354), .B(n_2385), .CI(n_2416), .CO(n_941), .S(n_940));
   FA_X1 i_471 (.A(n_2447), .B(n_2478), .CI(n_2509), .CO(n_943), .S(n_942));
   FA_X1 i_472 (.A(n_2540), .B(n_2571), .CI(n_2602), .CO(n_945), .S(n_944));
   FA_X1 i_473 (.A(n_2633), .B(n_2664), .CI(n_2695), .CO(n_947), .S(n_946));
   FA_X1 i_474 (.A(n_2726), .B(n_2757), .CI(n_2788), .CO(n_949), .S(n_948));
   FA_X1 i_475 (.A(n_2819), .B(n_889), .CI(n_887), .CO(n_951), .S(n_950));
   FA_X1 i_476 (.A(n_885), .B(n_883), .CI(n_881), .CO(n_953), .S(n_952));
   FA_X1 i_477 (.A(n_879), .B(n_877), .CI(n_875), .CO(n_955), .S(n_954));
   FA_X1 i_478 (.A(n_873), .B(n_871), .CI(n_897), .CO(n_957), .S(n_956));
   FA_X1 i_479 (.A(n_895), .B(n_893), .CI(n_891), .CO(n_959), .S(n_958));
   FA_X1 i_480 (.A(n_948), .B(n_946), .CI(n_944), .CO(n_961), .S(n_960));
   FA_X1 i_481 (.A(n_942), .B(n_940), .CI(n_938), .CO(n_963), .S(n_962));
   FA_X1 i_482 (.A(n_936), .B(n_934), .CI(n_932), .CO(n_965), .S(n_964));
   FA_X1 i_483 (.A(n_930), .B(n_899), .CI(n_956), .CO(n_967), .S(n_966));
   FA_X1 i_484 (.A(n_954), .B(n_952), .CI(n_950), .CO(n_969), .S(n_968));
   FA_X1 i_485 (.A(n_905), .B(n_903), .CI(n_901), .CO(n_971), .S(n_970));
   FA_X1 i_486 (.A(n_907), .B(n_958), .CI(n_911), .CO(n_973), .S(n_972));
   FA_X1 i_487 (.A(n_909), .B(n_964), .CI(n_962), .CO(n_975), .S(n_974));
   FA_X1 i_488 (.A(n_960), .B(n_966), .CI(n_913), .CO(n_977), .S(n_976));
   FA_X1 i_489 (.A(n_970), .B(n_968), .CI(n_915), .CO(n_979), .S(n_978));
   FA_X1 i_490 (.A(n_917), .B(n_972), .CI(n_919), .CO(n_981), .S(n_980));
   FA_X1 i_491 (.A(n_974), .B(n_976), .CI(n_921), .CO(n_983), .S(n_982));
   FA_X1 i_492 (.A(n_978), .B(n_923), .CI(n_980), .CO(n_985), .S(n_984));
   FA_X1 i_493 (.A(n_982), .B(n_925), .CI(n_984), .CO(n_987), .S(n_986));
   HA_X1 i_494 (.A(n_927), .B(n_986), .CO(n_989), .S(n_988));
   FA_X1 i_495 (.A(n_1888), .B(n_1919), .CI(n_1950), .CO(n_991), .S(n_990));
   FA_X1 i_496 (.A(n_1981), .B(n_2012), .CI(n_2043), .CO(n_993), .S(n_992));
   FA_X1 i_497 (.A(n_2074), .B(n_2105), .CI(n_2136), .CO(n_995), .S(n_994));
   FA_X1 i_498 (.A(n_2167), .B(n_2198), .CI(n_2229), .CO(n_997), .S(n_996));
   FA_X1 i_499 (.A(n_2260), .B(n_2291), .CI(n_2322), .CO(n_999), .S(n_998));
   FA_X1 i_500 (.A(n_2353), .B(n_2384), .CI(n_2415), .CO(n_1001), .S(n_1000));
   FA_X1 i_501 (.A(n_2446), .B(n_2477), .CI(n_2508), .CO(n_1003), .S(n_1002));
   FA_X1 i_502 (.A(n_2539), .B(n_2570), .CI(n_2601), .CO(n_1005), .S(n_1004));
   FA_X1 i_503 (.A(n_2632), .B(n_2663), .CI(n_2694), .CO(n_1007), .S(n_1006));
   FA_X1 i_504 (.A(n_2725), .B(n_2756), .CI(n_2787), .CO(n_1009), .S(n_1008));
   FA_X1 i_505 (.A(n_949), .B(n_947), .CI(n_945), .CO(n_1011), .S(n_1010));
   FA_X1 i_506 (.A(n_943), .B(n_941), .CI(n_939), .CO(n_1013), .S(n_1012));
   FA_X1 i_507 (.A(n_937), .B(n_935), .CI(n_933), .CO(n_1015), .S(n_1014));
   FA_X1 i_508 (.A(n_931), .B(n_955), .CI(n_953), .CO(n_1017), .S(n_1016));
   FA_X1 i_509 (.A(n_951), .B(n_1008), .CI(n_1006), .CO(n_1019), .S(n_1018));
   FA_X1 i_510 (.A(n_1004), .B(n_1002), .CI(n_1000), .CO(n_1021), .S(n_1020));
   FA_X1 i_511 (.A(n_998), .B(n_996), .CI(n_994), .CO(n_1023), .S(n_1022));
   FA_X1 i_512 (.A(n_992), .B(n_990), .CI(n_959), .CO(n_1025), .S(n_1024));
   FA_X1 i_513 (.A(n_957), .B(n_1014), .CI(n_1012), .CO(n_1027), .S(n_1026));
   FA_X1 i_514 (.A(n_1010), .B(n_965), .CI(n_963), .CO(n_1029), .S(n_1028));
   FA_X1 i_515 (.A(n_961), .B(n_1016), .CI(n_971), .CO(n_1031), .S(n_1030));
   FA_X1 i_516 (.A(n_969), .B(n_967), .CI(n_1024), .CO(n_1033), .S(n_1032));
   FA_X1 i_517 (.A(n_1022), .B(n_1020), .CI(n_1018), .CO(n_1035), .S(n_1034));
   FA_X1 i_518 (.A(n_973), .B(n_1028), .CI(n_1026), .CO(n_1037), .S(n_1036));
   FA_X1 i_519 (.A(n_975), .B(n_977), .CI(n_1032), .CO(n_1039), .S(n_1038));
   FA_X1 i_520 (.A(n_1030), .B(n_979), .CI(n_1034), .CO(n_1041), .S(n_1040));
   FA_X1 i_521 (.A(n_981), .B(n_1036), .CI(n_1038), .CO(n_1043), .S(n_1042));
   FA_X1 i_522 (.A(n_983), .B(n_1040), .CI(n_985), .CO(n_1045), .S(n_1044));
   FA_X1 i_523 (.A(n_1042), .B(n_1044), .CI(n_987), .CO(n_1047), .S(n_1046));
   FA_X1 i_524 (.A(n_1887), .B(n_1918), .CI(n_1949), .CO(n_1049), .S(n_1048));
   FA_X1 i_525 (.A(n_1980), .B(n_2011), .CI(n_2042), .CO(n_1051), .S(n_1050));
   FA_X1 i_526 (.A(n_2073), .B(n_2104), .CI(n_2135), .CO(n_1053), .S(n_1052));
   FA_X1 i_527 (.A(n_2166), .B(n_2197), .CI(n_2228), .CO(n_1055), .S(n_1054));
   FA_X1 i_528 (.A(n_2259), .B(n_2290), .CI(n_2321), .CO(n_1057), .S(n_1056));
   FA_X1 i_529 (.A(n_2352), .B(n_2383), .CI(n_2414), .CO(n_1059), .S(n_1058));
   FA_X1 i_530 (.A(n_2445), .B(n_2476), .CI(n_2507), .CO(n_1061), .S(n_1060));
   FA_X1 i_531 (.A(n_2538), .B(n_2569), .CI(n_2600), .CO(n_1063), .S(n_1062));
   FA_X1 i_532 (.A(n_2631), .B(n_2662), .CI(n_2693), .CO(n_1065), .S(n_1064));
   FA_X1 i_533 (.A(n_2724), .B(n_2755), .CI(n_1009), .CO(n_1067), .S(n_1066));
   FA_X1 i_534 (.A(n_1007), .B(n_1005), .CI(n_1003), .CO(n_1069), .S(n_1068));
   FA_X1 i_535 (.A(n_1001), .B(n_999), .CI(n_997), .CO(n_1071), .S(n_1070));
   FA_X1 i_536 (.A(n_995), .B(n_993), .CI(n_991), .CO(n_1073), .S(n_1072));
   FA_X1 i_537 (.A(n_1015), .B(n_1013), .CI(n_1011), .CO(n_1075), .S(n_1074));
   FA_X1 i_538 (.A(n_1066), .B(n_1064), .CI(n_1062), .CO(n_1077), .S(n_1076));
   FA_X1 i_539 (.A(n_1060), .B(n_1058), .CI(n_1056), .CO(n_1079), .S(n_1078));
   FA_X1 i_540 (.A(n_1054), .B(n_1052), .CI(n_1050), .CO(n_1081), .S(n_1080));
   FA_X1 i_541 (.A(n_1048), .B(n_1017), .CI(n_1072), .CO(n_1083), .S(n_1082));
   FA_X1 i_542 (.A(n_1070), .B(n_1068), .CI(n_1023), .CO(n_1085), .S(n_1084));
   FA_X1 i_543 (.A(n_1021), .B(n_1019), .CI(n_1025), .CO(n_1087), .S(n_1086));
   FA_X1 i_544 (.A(n_1074), .B(n_1029), .CI(n_1027), .CO(n_1089), .S(n_1088));
   FA_X1 i_545 (.A(n_1080), .B(n_1078), .CI(n_1076), .CO(n_1091), .S(n_1090));
   FA_X1 i_546 (.A(n_1082), .B(n_1031), .CI(n_1086), .CO(n_1093), .S(n_1092));
   FA_X1 i_547 (.A(n_1084), .B(n_1035), .CI(n_1033), .CO(n_1095), .S(n_1094));
   FA_X1 i_548 (.A(n_1088), .B(n_1037), .CI(n_1090), .CO(n_1097), .S(n_1096));
   FA_X1 i_549 (.A(n_1092), .B(n_1039), .CI(n_1094), .CO(n_1099), .S(n_1098));
   FA_X1 i_550 (.A(n_1041), .B(n_1096), .CI(n_1043), .CO(n_1101), .S(n_1100));
   FA_X1 i_551 (.A(n_1098), .B(n_1045), .CI(n_1100), .CO(n_1103), .S(n_1102));
   FA_X1 i_552 (.A(n_1886), .B(n_1917), .CI(n_1948), .CO(n_1105), .S(n_1104));
   FA_X1 i_553 (.A(n_1979), .B(n_2010), .CI(n_2041), .CO(n_1107), .S(n_1106));
   FA_X1 i_554 (.A(n_2072), .B(n_2103), .CI(n_2134), .CO(n_1109), .S(n_1108));
   FA_X1 i_555 (.A(n_2165), .B(n_2196), .CI(n_2227), .CO(n_1111), .S(n_1110));
   FA_X1 i_556 (.A(n_2258), .B(n_2289), .CI(n_2320), .CO(n_1113), .S(n_1112));
   FA_X1 i_557 (.A(n_2351), .B(n_2382), .CI(n_2413), .CO(n_1115), .S(n_1114));
   FA_X1 i_558 (.A(n_2444), .B(n_2475), .CI(n_2506), .CO(n_1117), .S(n_1116));
   FA_X1 i_559 (.A(n_2537), .B(n_2568), .CI(n_2599), .CO(n_1119), .S(n_1118));
   FA_X1 i_560 (.A(n_2630), .B(n_2661), .CI(n_2692), .CO(n_1121), .S(n_1120));
   FA_X1 i_561 (.A(n_2723), .B(n_1065), .CI(n_1063), .CO(n_1123), .S(n_1122));
   FA_X1 i_562 (.A(n_1061), .B(n_1059), .CI(n_1057), .CO(n_1125), .S(n_1124));
   FA_X1 i_563 (.A(n_1055), .B(n_1053), .CI(n_1051), .CO(n_1127), .S(n_1126));
   FA_X1 i_564 (.A(n_1049), .B(n_1073), .CI(n_1071), .CO(n_1129), .S(n_1128));
   FA_X1 i_565 (.A(n_1069), .B(n_1067), .CI(n_1120), .CO(n_1131), .S(n_1130));
   FA_X1 i_566 (.A(n_1118), .B(n_1116), .CI(n_1114), .CO(n_1133), .S(n_1132));
   FA_X1 i_567 (.A(n_1112), .B(n_1110), .CI(n_1108), .CO(n_1135), .S(n_1134));
   FA_X1 i_568 (.A(n_1106), .B(n_1104), .CI(n_1075), .CO(n_1137), .S(n_1136));
   FA_X1 i_569 (.A(n_1126), .B(n_1124), .CI(n_1122), .CO(n_1139), .S(n_1138));
   FA_X1 i_570 (.A(n_1081), .B(n_1079), .CI(n_1077), .CO(n_1141), .S(n_1140));
   FA_X1 i_571 (.A(n_1130), .B(n_1128), .CI(n_1085), .CO(n_1143), .S(n_1142));
   FA_X1 i_572 (.A(n_1083), .B(n_1087), .CI(n_1136), .CO(n_1145), .S(n_1144));
   FA_X1 i_573 (.A(n_1134), .B(n_1132), .CI(n_1089), .CO(n_1147), .S(n_1146));
   FA_X1 i_574 (.A(n_1140), .B(n_1138), .CI(n_1091), .CO(n_1149), .S(n_1148));
   FA_X1 i_575 (.A(n_1142), .B(n_1095), .CI(n_1093), .CO(n_1151), .S(n_1150));
   FA_X1 i_576 (.A(n_1144), .B(n_1146), .CI(n_1148), .CO(n_1153), .S(n_1152));
   FA_X1 i_577 (.A(n_1097), .B(n_1150), .CI(n_1099), .CO(n_1155), .S(n_1154));
   FA_X1 i_578 (.A(n_1152), .B(n_1101), .CI(n_1154), .CO(n_1157), .S(n_1156));
   FA_X1 i_579 (.A(n_1885), .B(n_1916), .CI(n_1947), .CO(n_1159), .S(n_1158));
   FA_X1 i_580 (.A(n_1978), .B(n_2009), .CI(n_2040), .CO(n_1161), .S(n_1160));
   FA_X1 i_581 (.A(n_2071), .B(n_2102), .CI(n_2133), .CO(n_1163), .S(n_1162));
   FA_X1 i_582 (.A(n_2164), .B(n_2195), .CI(n_2226), .CO(n_1165), .S(n_1164));
   FA_X1 i_583 (.A(n_2257), .B(n_2288), .CI(n_2319), .CO(n_1167), .S(n_1166));
   FA_X1 i_584 (.A(n_2350), .B(n_2381), .CI(n_2412), .CO(n_1169), .S(n_1168));
   FA_X1 i_585 (.A(n_2443), .B(n_2474), .CI(n_2505), .CO(n_1171), .S(n_1170));
   FA_X1 i_586 (.A(n_2536), .B(n_2567), .CI(n_2598), .CO(n_1173), .S(n_1172));
   FA_X1 i_587 (.A(n_2629), .B(n_2660), .CI(n_2691), .CO(n_1175), .S(n_1174));
   FA_X1 i_588 (.A(n_1121), .B(n_1119), .CI(n_1117), .CO(n_1177), .S(n_1176));
   FA_X1 i_589 (.A(n_1115), .B(n_1113), .CI(n_1111), .CO(n_1179), .S(n_1178));
   FA_X1 i_590 (.A(n_1109), .B(n_1107), .CI(n_1105), .CO(n_1181), .S(n_1180));
   FA_X1 i_591 (.A(n_1127), .B(n_1125), .CI(n_1123), .CO(n_1183), .S(n_1182));
   FA_X1 i_592 (.A(n_1174), .B(n_1172), .CI(n_1170), .CO(n_1185), .S(n_1184));
   FA_X1 i_593 (.A(n_1168), .B(n_1166), .CI(n_1164), .CO(n_1187), .S(n_1186));
   FA_X1 i_594 (.A(n_1162), .B(n_1160), .CI(n_1158), .CO(n_1189), .S(n_1188));
   FA_X1 i_595 (.A(n_1129), .B(n_1180), .CI(n_1178), .CO(n_1191), .S(n_1190));
   FA_X1 i_596 (.A(n_1176), .B(n_1135), .CI(n_1133), .CO(n_1193), .S(n_1192));
   FA_X1 i_597 (.A(n_1131), .B(n_1137), .CI(n_1182), .CO(n_1195), .S(n_1194));
   FA_X1 i_598 (.A(n_1141), .B(n_1139), .CI(n_1188), .CO(n_1197), .S(n_1196));
   FA_X1 i_599 (.A(n_1186), .B(n_1184), .CI(n_1143), .CO(n_1199), .S(n_1198));
   FA_X1 i_600 (.A(n_1192), .B(n_1190), .CI(n_1145), .CO(n_1201), .S(n_1200));
   FA_X1 i_601 (.A(n_1194), .B(n_1147), .CI(n_1196), .CO(n_1203), .S(n_1202));
   FA_X1 i_602 (.A(n_1149), .B(n_1198), .CI(n_1151), .CO(n_1205), .S(n_1204));
   FA_X1 i_603 (.A(n_1200), .B(n_1202), .CI(n_1153), .CO(n_1207), .S(n_1206));
   FA_X1 i_604 (.A(n_1204), .B(n_1155), .CI(n_1206), .CO(n_1209), .S(n_1208));
   FA_X1 i_605 (.A(n_1884), .B(n_1915), .CI(n_1946), .CO(n_1211), .S(n_1210));
   FA_X1 i_606 (.A(n_1977), .B(n_2008), .CI(n_2039), .CO(n_1213), .S(n_1212));
   FA_X1 i_607 (.A(n_2070), .B(n_2101), .CI(n_2132), .CO(n_1215), .S(n_1214));
   FA_X1 i_608 (.A(n_2163), .B(n_2194), .CI(n_2225), .CO(n_1217), .S(n_1216));
   FA_X1 i_609 (.A(n_2256), .B(n_2287), .CI(n_2318), .CO(n_1219), .S(n_1218));
   FA_X1 i_610 (.A(n_2349), .B(n_2380), .CI(n_2411), .CO(n_1221), .S(n_1220));
   FA_X1 i_611 (.A(n_2442), .B(n_2473), .CI(n_2504), .CO(n_1223), .S(n_1222));
   FA_X1 i_612 (.A(n_2535), .B(n_2566), .CI(n_2597), .CO(n_1225), .S(n_1224));
   FA_X1 i_613 (.A(n_2628), .B(n_2659), .CI(n_1175), .CO(n_1227), .S(n_1226));
   FA_X1 i_614 (.A(n_1173), .B(n_1171), .CI(n_1169), .CO(n_1229), .S(n_1228));
   FA_X1 i_615 (.A(n_1167), .B(n_1165), .CI(n_1163), .CO(n_1231), .S(n_1230));
   FA_X1 i_616 (.A(n_1161), .B(n_1159), .CI(n_1181), .CO(n_1233), .S(n_1232));
   FA_X1 i_617 (.A(n_1179), .B(n_1177), .CI(n_1226), .CO(n_1235), .S(n_1234));
   FA_X1 i_618 (.A(n_1224), .B(n_1222), .CI(n_1220), .CO(n_1237), .S(n_1236));
   FA_X1 i_619 (.A(n_1218), .B(n_1216), .CI(n_1214), .CO(n_1239), .S(n_1238));
   FA_X1 i_620 (.A(n_1212), .B(n_1210), .CI(n_1183), .CO(n_1241), .S(n_1240));
   FA_X1 i_621 (.A(n_1232), .B(n_1230), .CI(n_1228), .CO(n_1243), .S(n_1242));
   FA_X1 i_622 (.A(n_1189), .B(n_1187), .CI(n_1185), .CO(n_1245), .S(n_1244));
   FA_X1 i_623 (.A(n_1234), .B(n_1193), .CI(n_1191), .CO(n_1247), .S(n_1246));
   FA_X1 i_624 (.A(n_1240), .B(n_1238), .CI(n_1236), .CO(n_1249), .S(n_1248));
   FA_X1 i_625 (.A(n_1195), .B(n_1244), .CI(n_1242), .CO(n_1251), .S(n_1250));
   FA_X1 i_626 (.A(n_1197), .B(n_1199), .CI(n_1246), .CO(n_1253), .S(n_1252));
   FA_X1 i_627 (.A(n_1201), .B(n_1248), .CI(n_1203), .CO(n_1255), .S(n_1254));
   FA_X1 i_628 (.A(n_1250), .B(n_1252), .CI(n_1205), .CO(n_1257), .S(n_1256));
   FA_X1 i_629 (.A(n_1254), .B(n_1207), .CI(n_1256), .CO(n_1259), .S(n_1258));
   FA_X1 i_630 (.A(n_1883), .B(n_1914), .CI(n_1945), .CO(n_1261), .S(n_1260));
   FA_X1 i_631 (.A(n_1976), .B(n_2007), .CI(n_2038), .CO(n_1263), .S(n_1262));
   FA_X1 i_632 (.A(n_2069), .B(n_2100), .CI(n_2131), .CO(n_1265), .S(n_1264));
   FA_X1 i_633 (.A(n_2162), .B(n_2193), .CI(n_2224), .CO(n_1267), .S(n_1266));
   FA_X1 i_634 (.A(n_2255), .B(n_2286), .CI(n_2317), .CO(n_1269), .S(n_1268));
   FA_X1 i_635 (.A(n_2348), .B(n_2379), .CI(n_2410), .CO(n_1271), .S(n_1270));
   FA_X1 i_636 (.A(n_2441), .B(n_2472), .CI(n_2503), .CO(n_1273), .S(n_1272));
   FA_X1 i_637 (.A(n_2534), .B(n_2565), .CI(n_2596), .CO(n_1275), .S(n_1274));
   FA_X1 i_638 (.A(n_2627), .B(n_1225), .CI(n_1223), .CO(n_1277), .S(n_1276));
   FA_X1 i_639 (.A(n_1221), .B(n_1219), .CI(n_1217), .CO(n_1279), .S(n_1278));
   FA_X1 i_640 (.A(n_1215), .B(n_1213), .CI(n_1211), .CO(n_1281), .S(n_1280));
   FA_X1 i_641 (.A(n_1231), .B(n_1229), .CI(n_1227), .CO(n_1283), .S(n_1282));
   FA_X1 i_642 (.A(n_1274), .B(n_1272), .CI(n_1270), .CO(n_1285), .S(n_1284));
   FA_X1 i_643 (.A(n_1268), .B(n_1266), .CI(n_1264), .CO(n_1287), .S(n_1286));
   FA_X1 i_644 (.A(n_1262), .B(n_1260), .CI(n_1233), .CO(n_1289), .S(n_1288));
   FA_X1 i_645 (.A(n_1280), .B(n_1278), .CI(n_1276), .CO(n_1291), .S(n_1290));
   FA_X1 i_646 (.A(n_1239), .B(n_1237), .CI(n_1235), .CO(n_1293), .S(n_1292));
   FA_X1 i_647 (.A(n_1241), .B(n_1282), .CI(n_1245), .CO(n_1295), .S(n_1294));
   FA_X1 i_648 (.A(n_1243), .B(n_1288), .CI(n_1286), .CO(n_1297), .S(n_1296));
   FA_X1 i_649 (.A(n_1284), .B(n_1247), .CI(n_1292), .CO(n_1299), .S(n_1298));
   FA_X1 i_650 (.A(n_1290), .B(n_1249), .CI(n_1294), .CO(n_1301), .S(n_1300));
   FA_X1 i_651 (.A(n_1251), .B(n_1296), .CI(n_1298), .CO(n_1303), .S(n_1302));
   FA_X1 i_652 (.A(n_1253), .B(n_1300), .CI(n_1255), .CO(n_1305), .S(n_1304));
   FA_X1 i_653 (.A(n_1257), .B(n_1302), .CI(n_1304), .CO(n_1307), .S(n_1306));
   FA_X1 i_654 (.A(n_1882), .B(n_1913), .CI(n_1944), .CO(n_1309), .S(n_1308));
   FA_X1 i_655 (.A(n_1975), .B(n_2006), .CI(n_2037), .CO(n_1311), .S(n_1310));
   FA_X1 i_656 (.A(n_2068), .B(n_2099), .CI(n_2130), .CO(n_1313), .S(n_1312));
   FA_X1 i_657 (.A(n_2161), .B(n_2192), .CI(n_2223), .CO(n_1315), .S(n_1314));
   FA_X1 i_658 (.A(n_2254), .B(n_2285), .CI(n_2316), .CO(n_1317), .S(n_1316));
   FA_X1 i_659 (.A(n_2347), .B(n_2378), .CI(n_2409), .CO(n_1319), .S(n_1318));
   FA_X1 i_660 (.A(n_2440), .B(n_2471), .CI(n_2502), .CO(n_1321), .S(n_1320));
   FA_X1 i_661 (.A(n_2533), .B(n_2564), .CI(n_2595), .CO(n_1323), .S(n_1322));
   FA_X1 i_662 (.A(n_1275), .B(n_1273), .CI(n_1271), .CO(n_1325), .S(n_1324));
   FA_X1 i_663 (.A(n_1269), .B(n_1267), .CI(n_1265), .CO(n_1327), .S(n_1326));
   FA_X1 i_664 (.A(n_1263), .B(n_1261), .CI(n_1281), .CO(n_1329), .S(n_1328));
   FA_X1 i_665 (.A(n_1279), .B(n_1277), .CI(n_1322), .CO(n_1331), .S(n_1330));
   FA_X1 i_666 (.A(n_1320), .B(n_1318), .CI(n_1316), .CO(n_1333), .S(n_1332));
   FA_X1 i_667 (.A(n_1314), .B(n_1312), .CI(n_1310), .CO(n_1335), .S(n_1334));
   FA_X1 i_668 (.A(n_1308), .B(n_1283), .CI(n_1328), .CO(n_1337), .S(n_1336));
   FA_X1 i_669 (.A(n_1326), .B(n_1324), .CI(n_1287), .CO(n_1339), .S(n_1338));
   FA_X1 i_670 (.A(n_1285), .B(n_1289), .CI(n_1330), .CO(n_1341), .S(n_1340));
   FA_X1 i_671 (.A(n_1293), .B(n_1291), .CI(n_1334), .CO(n_1343), .S(n_1342));
   FA_X1 i_672 (.A(n_1332), .B(n_1336), .CI(n_1295), .CO(n_1345), .S(n_1344));
   FA_X1 i_673 (.A(n_1338), .B(n_1297), .CI(n_1340), .CO(n_1347), .S(n_1346));
   FA_X1 i_674 (.A(n_1342), .B(n_1299), .CI(n_1344), .CO(n_1349), .S(n_1348));
   FA_X1 i_675 (.A(n_1301), .B(n_1346), .CI(n_1303), .CO(n_1351), .S(n_1350));
   FA_X1 i_676 (.A(n_1348), .B(n_1305), .CI(n_1350), .CO(n_1353), .S(n_1352));
   FA_X1 i_677 (.A(n_1881), .B(n_1912), .CI(n_1943), .CO(n_1355), .S(n_1354));
   FA_X1 i_678 (.A(n_1974), .B(n_2005), .CI(n_2036), .CO(n_1357), .S(n_1356));
   FA_X1 i_679 (.A(n_2067), .B(n_2098), .CI(n_2129), .CO(n_1359), .S(n_1358));
   FA_X1 i_680 (.A(n_2160), .B(n_2191), .CI(n_2222), .CO(n_1361), .S(n_1360));
   FA_X1 i_681 (.A(n_2253), .B(n_2284), .CI(n_2315), .CO(n_1363), .S(n_1362));
   FA_X1 i_682 (.A(n_2346), .B(n_2377), .CI(n_2408), .CO(n_1365), .S(n_1364));
   FA_X1 i_683 (.A(n_2439), .B(n_2470), .CI(n_2501), .CO(n_1367), .S(n_1366));
   FA_X1 i_684 (.A(n_2532), .B(n_2563), .CI(n_1323), .CO(n_1369), .S(n_1368));
   FA_X1 i_685 (.A(n_1321), .B(n_1319), .CI(n_1317), .CO(n_1371), .S(n_1370));
   FA_X1 i_686 (.A(n_1315), .B(n_1313), .CI(n_1311), .CO(n_1373), .S(n_1372));
   FA_X1 i_687 (.A(n_1309), .B(n_1327), .CI(n_1325), .CO(n_1375), .S(n_1374));
   FA_X1 i_688 (.A(n_1368), .B(n_1366), .CI(n_1364), .CO(n_1377), .S(n_1376));
   FA_X1 i_689 (.A(n_1362), .B(n_1360), .CI(n_1358), .CO(n_1379), .S(n_1378));
   FA_X1 i_690 (.A(n_1356), .B(n_1354), .CI(n_1329), .CO(n_1381), .S(n_1380));
   FA_X1 i_691 (.A(n_1372), .B(n_1370), .CI(n_1335), .CO(n_1383), .S(n_1382));
   FA_X1 i_692 (.A(n_1333), .B(n_1331), .CI(n_1374), .CO(n_1385), .S(n_1384));
   FA_X1 i_693 (.A(n_1339), .B(n_1337), .CI(n_1380), .CO(n_1387), .S(n_1386));
   FA_X1 i_694 (.A(n_1378), .B(n_1376), .CI(n_1341), .CO(n_1389), .S(n_1388));
   FA_X1 i_695 (.A(n_1384), .B(n_1382), .CI(n_1343), .CO(n_1391), .S(n_1390));
   FA_X1 i_696 (.A(n_1345), .B(n_1386), .CI(n_1347), .CO(n_1393), .S(n_1392));
   FA_X1 i_697 (.A(n_1388), .B(n_1390), .CI(n_1349), .CO(n_1395), .S(n_1394));
   FA_X1 i_698 (.A(n_1392), .B(n_1351), .CI(n_1394), .CO(n_1397), .S(n_1396));
   FA_X1 i_699 (.A(n_1880), .B(n_1911), .CI(n_1942), .CO(n_1399), .S(n_1398));
   FA_X1 i_700 (.A(n_1973), .B(n_2004), .CI(n_2035), .CO(n_1401), .S(n_1400));
   FA_X1 i_701 (.A(n_2066), .B(n_2097), .CI(n_2128), .CO(n_1403), .S(n_1402));
   FA_X1 i_702 (.A(n_2159), .B(n_2190), .CI(n_2221), .CO(n_1405), .S(n_1404));
   FA_X1 i_703 (.A(n_2252), .B(n_2283), .CI(n_2314), .CO(n_1407), .S(n_1406));
   FA_X1 i_704 (.A(n_2345), .B(n_2376), .CI(n_2407), .CO(n_1409), .S(n_1408));
   FA_X1 i_705 (.A(n_2438), .B(n_2469), .CI(n_2500), .CO(n_1411), .S(n_1410));
   FA_X1 i_706 (.A(n_2531), .B(n_1367), .CI(n_1365), .CO(n_1413), .S(n_1412));
   FA_X1 i_707 (.A(n_1363), .B(n_1361), .CI(n_1359), .CO(n_1415), .S(n_1414));
   FA_X1 i_708 (.A(n_1357), .B(n_1355), .CI(n_1373), .CO(n_1417), .S(n_1416));
   FA_X1 i_709 (.A(n_1371), .B(n_1369), .CI(n_1410), .CO(n_1419), .S(n_1418));
   FA_X1 i_710 (.A(n_1408), .B(n_1406), .CI(n_1404), .CO(n_1421), .S(n_1420));
   FA_X1 i_711 (.A(n_1402), .B(n_1400), .CI(n_1398), .CO(n_1423), .S(n_1422));
   FA_X1 i_712 (.A(n_1375), .B(n_1416), .CI(n_1414), .CO(n_1425), .S(n_1424));
   FA_X1 i_713 (.A(n_1412), .B(n_1379), .CI(n_1377), .CO(n_1427), .S(n_1426));
   FA_X1 i_714 (.A(n_1381), .B(n_1418), .CI(n_1383), .CO(n_1429), .S(n_1428));
   FA_X1 i_715 (.A(n_1422), .B(n_1420), .CI(n_1385), .CO(n_1431), .S(n_1430));
   FA_X1 i_716 (.A(n_1426), .B(n_1424), .CI(n_1387), .CO(n_1433), .S(n_1432));
   FA_X1 i_717 (.A(n_1389), .B(n_1428), .CI(n_1391), .CO(n_1435), .S(n_1434));
   FA_X1 i_718 (.A(n_1430), .B(n_1393), .CI(n_1432), .CO(n_1437), .S(n_1436));
   FA_X1 i_719 (.A(n_1434), .B(n_1395), .CI(n_1436), .CO(n_1439), .S(n_1438));
   FA_X1 i_720 (.A(n_1879), .B(n_1910), .CI(n_1941), .CO(n_1441), .S(n_1440));
   FA_X1 i_721 (.A(n_1972), .B(n_2003), .CI(n_2034), .CO(n_1443), .S(n_1442));
   FA_X1 i_722 (.A(n_2065), .B(n_2096), .CI(n_2127), .CO(n_1445), .S(n_1444));
   FA_X1 i_723 (.A(n_2158), .B(n_2189), .CI(n_2220), .CO(n_1447), .S(n_1446));
   FA_X1 i_724 (.A(n_2251), .B(n_2282), .CI(n_2313), .CO(n_1449), .S(n_1448));
   FA_X1 i_725 (.A(n_2344), .B(n_2375), .CI(n_2406), .CO(n_1451), .S(n_1450));
   FA_X1 i_726 (.A(n_2437), .B(n_2468), .CI(n_2499), .CO(n_1453), .S(n_1452));
   FA_X1 i_727 (.A(n_1411), .B(n_1409), .CI(n_1407), .CO(n_1455), .S(n_1454));
   FA_X1 i_728 (.A(n_1405), .B(n_1403), .CI(n_1401), .CO(n_1457), .S(n_1456));
   FA_X1 i_729 (.A(n_1399), .B(n_1415), .CI(n_1413), .CO(n_1459), .S(n_1458));
   FA_X1 i_730 (.A(n_1452), .B(n_1450), .CI(n_1448), .CO(n_1461), .S(n_1460));
   FA_X1 i_731 (.A(n_1446), .B(n_1444), .CI(n_1442), .CO(n_1463), .S(n_1462));
   FA_X1 i_732 (.A(n_1440), .B(n_1417), .CI(n_1456), .CO(n_1465), .S(n_1464));
   FA_X1 i_733 (.A(n_1454), .B(n_1423), .CI(n_1421), .CO(n_1467), .S(n_1466));
   FA_X1 i_734 (.A(n_1419), .B(n_1458), .CI(n_1427), .CO(n_1469), .S(n_1468));
   FA_X1 i_735 (.A(n_1425), .B(n_1462), .CI(n_1460), .CO(n_1471), .S(n_1470));
   FA_X1 i_736 (.A(n_1464), .B(n_1429), .CI(n_1466), .CO(n_1473), .S(n_1472));
   FA_X1 i_737 (.A(n_1431), .B(n_1468), .CI(n_1433), .CO(n_1475), .S(n_1474));
   FA_X1 i_738 (.A(n_1470), .B(n_1472), .CI(n_1435), .CO(n_1477), .S(n_1476));
   FA_X1 i_739 (.A(n_1474), .B(n_1437), .CI(n_1476), .CO(n_1479), .S(n_1478));
   FA_X1 i_740 (.A(n_1878), .B(n_1909), .CI(n_1940), .CO(n_1481), .S(n_1480));
   FA_X1 i_741 (.A(n_1971), .B(n_2002), .CI(n_2033), .CO(n_1483), .S(n_1482));
   FA_X1 i_742 (.A(n_2064), .B(n_2095), .CI(n_2126), .CO(n_1485), .S(n_1484));
   FA_X1 i_743 (.A(n_2157), .B(n_2188), .CI(n_2219), .CO(n_1487), .S(n_1486));
   FA_X1 i_744 (.A(n_2250), .B(n_2281), .CI(n_2312), .CO(n_1489), .S(n_1488));
   FA_X1 i_745 (.A(n_2343), .B(n_2374), .CI(n_2405), .CO(n_1491), .S(n_1490));
   FA_X1 i_746 (.A(n_2436), .B(n_2467), .CI(n_1453), .CO(n_1493), .S(n_1492));
   FA_X1 i_747 (.A(n_1451), .B(n_1449), .CI(n_1447), .CO(n_1495), .S(n_1494));
   FA_X1 i_748 (.A(n_1445), .B(n_1443), .CI(n_1441), .CO(n_1497), .S(n_1496));
   FA_X1 i_749 (.A(n_1457), .B(n_1455), .CI(n_1492), .CO(n_1499), .S(n_1498));
   FA_X1 i_750 (.A(n_1490), .B(n_1488), .CI(n_1486), .CO(n_1501), .S(n_1500));
   FA_X1 i_751 (.A(n_1484), .B(n_1482), .CI(n_1480), .CO(n_1503), .S(n_1502));
   FA_X1 i_752 (.A(n_1459), .B(n_1496), .CI(n_1494), .CO(n_1505), .S(n_1504));
   FA_X1 i_753 (.A(n_1463), .B(n_1461), .CI(n_1498), .CO(n_1507), .S(n_1506));
   FA_X1 i_754 (.A(n_1467), .B(n_1465), .CI(n_1502), .CO(n_1509), .S(n_1508));
   FA_X1 i_755 (.A(n_1500), .B(n_1469), .CI(n_1506), .CO(n_1511), .S(n_1510));
   FA_X1 i_756 (.A(n_1504), .B(n_1471), .CI(n_1508), .CO(n_1513), .S(n_1512));
   FA_X1 i_757 (.A(n_1473), .B(n_1510), .CI(n_1475), .CO(n_1515), .S(n_1514));
   FA_X1 i_758 (.A(n_1512), .B(n_1477), .CI(n_1514), .CO(n_1517), .S(n_1516));
   FA_X1 i_759 (.A(n_1877), .B(n_1908), .CI(n_1939), .CO(n_1519), .S(n_1518));
   FA_X1 i_760 (.A(n_1970), .B(n_2001), .CI(n_2032), .CO(n_1521), .S(n_1520));
   FA_X1 i_761 (.A(n_2063), .B(n_2094), .CI(n_2125), .CO(n_1523), .S(n_1522));
   FA_X1 i_762 (.A(n_2156), .B(n_2187), .CI(n_2218), .CO(n_1525), .S(n_1524));
   FA_X1 i_763 (.A(n_2249), .B(n_2280), .CI(n_2311), .CO(n_1527), .S(n_1526));
   FA_X1 i_764 (.A(n_2342), .B(n_2373), .CI(n_2404), .CO(n_1529), .S(n_1528));
   FA_X1 i_765 (.A(n_2435), .B(n_1491), .CI(n_1489), .CO(n_1531), .S(n_1530));
   FA_X1 i_766 (.A(n_1487), .B(n_1485), .CI(n_1483), .CO(n_1533), .S(n_1532));
   FA_X1 i_767 (.A(n_1481), .B(n_1497), .CI(n_1495), .CO(n_1535), .S(n_1534));
   FA_X1 i_768 (.A(n_1493), .B(n_1528), .CI(n_1526), .CO(n_1537), .S(n_1536));
   FA_X1 i_769 (.A(n_1524), .B(n_1522), .CI(n_1520), .CO(n_1539), .S(n_1538));
   FA_X1 i_770 (.A(n_1518), .B(n_1532), .CI(n_1530), .CO(n_1541), .S(n_1540));
   FA_X1 i_771 (.A(n_1503), .B(n_1501), .CI(n_1499), .CO(n_1543), .S(n_1542));
   FA_X1 i_772 (.A(n_1534), .B(n_1505), .CI(n_1538), .CO(n_1545), .S(n_1544));
   FA_X1 i_773 (.A(n_1536), .B(n_1507), .CI(n_1542), .CO(n_1547), .S(n_1546));
   FA_X1 i_774 (.A(n_1540), .B(n_1509), .CI(n_1544), .CO(n_1549), .S(n_1548));
   FA_X1 i_775 (.A(n_1511), .B(n_1546), .CI(n_1513), .CO(n_1551), .S(n_1550));
   FA_X1 i_776 (.A(n_1548), .B(n_1515), .CI(n_1550), .CO(n_1553), .S(n_1552));
   FA_X1 i_777 (.A(n_1876), .B(n_1907), .CI(n_1938), .CO(n_1555), .S(n_1554));
   FA_X1 i_778 (.A(n_1969), .B(n_2000), .CI(n_2031), .CO(n_1557), .S(n_1556));
   FA_X1 i_779 (.A(n_2062), .B(n_2093), .CI(n_2124), .CO(n_1559), .S(n_1558));
   FA_X1 i_780 (.A(n_2155), .B(n_2186), .CI(n_2217), .CO(n_1561), .S(n_1560));
   FA_X1 i_781 (.A(n_2248), .B(n_2279), .CI(n_2310), .CO(n_1563), .S(n_1562));
   FA_X1 i_782 (.A(n_2341), .B(n_2372), .CI(n_2403), .CO(n_1565), .S(n_1564));
   FA_X1 i_783 (.A(n_1529), .B(n_1527), .CI(n_1525), .CO(n_1567), .S(n_1566));
   FA_X1 i_784 (.A(n_1523), .B(n_1521), .CI(n_1519), .CO(n_1569), .S(n_1568));
   FA_X1 i_785 (.A(n_1533), .B(n_1531), .CI(n_1564), .CO(n_1571), .S(n_1570));
   FA_X1 i_786 (.A(n_1562), .B(n_1560), .CI(n_1558), .CO(n_1573), .S(n_1572));
   FA_X1 i_787 (.A(n_1556), .B(n_1554), .CI(n_1535), .CO(n_1575), .S(n_1574));
   FA_X1 i_788 (.A(n_1568), .B(n_1566), .CI(n_1539), .CO(n_1577), .S(n_1576));
   FA_X1 i_789 (.A(n_1537), .B(n_1570), .CI(n_1543), .CO(n_1579), .S(n_1578));
   FA_X1 i_790 (.A(n_1541), .B(n_1574), .CI(n_1572), .CO(n_1581), .S(n_1580));
   FA_X1 i_791 (.A(n_1576), .B(n_1545), .CI(n_1578), .CO(n_1583), .S(n_1582));
   FA_X1 i_792 (.A(n_1547), .B(n_1580), .CI(n_1549), .CO(n_1585), .S(n_1584));
   FA_X1 i_793 (.A(n_1582), .B(n_1551), .CI(n_1584), .CO(n_1587), .S(n_1586));
   FA_X1 i_794 (.A(n_1875), .B(n_1906), .CI(n_1937), .CO(n_1589), .S(n_1588));
   FA_X1 i_795 (.A(n_1968), .B(n_1999), .CI(n_2030), .CO(n_1591), .S(n_1590));
   FA_X1 i_796 (.A(n_2061), .B(n_2092), .CI(n_2123), .CO(n_1593), .S(n_1592));
   FA_X1 i_797 (.A(n_2154), .B(n_2185), .CI(n_2216), .CO(n_1595), .S(n_1594));
   FA_X1 i_798 (.A(n_2247), .B(n_2278), .CI(n_2309), .CO(n_1597), .S(n_1596));
   FA_X1 i_799 (.A(n_2340), .B(n_2371), .CI(n_1565), .CO(n_1599), .S(n_1598));
   FA_X1 i_800 (.A(n_1563), .B(n_1561), .CI(n_1559), .CO(n_1601), .S(n_1600));
   FA_X1 i_801 (.A(n_1557), .B(n_1555), .CI(n_1569), .CO(n_1603), .S(n_1602));
   FA_X1 i_802 (.A(n_1567), .B(n_1598), .CI(n_1596), .CO(n_1605), .S(n_1604));
   FA_X1 i_803 (.A(n_1594), .B(n_1592), .CI(n_1590), .CO(n_1607), .S(n_1606));
   FA_X1 i_804 (.A(n_1588), .B(n_1602), .CI(n_1600), .CO(n_1609), .S(n_1608));
   FA_X1 i_805 (.A(n_1573), .B(n_1571), .CI(n_1575), .CO(n_1611), .S(n_1610));
   FA_X1 i_806 (.A(n_1577), .B(n_1606), .CI(n_1604), .CO(n_1613), .S(n_1612));
   FA_X1 i_807 (.A(n_1579), .B(n_1610), .CI(n_1608), .CO(n_1615), .S(n_1614));
   FA_X1 i_808 (.A(n_1581), .B(n_1612), .CI(n_1583), .CO(n_1617), .S(n_1616));
   FA_X1 i_809 (.A(n_1614), .B(n_1585), .CI(n_1616), .CO(n_1619), .S(n_1618));
   FA_X1 i_810 (.A(n_1874), .B(n_1905), .CI(n_1936), .CO(n_1621), .S(n_1620));
   FA_X1 i_811 (.A(n_1967), .B(n_1998), .CI(n_2029), .CO(n_1623), .S(n_1622));
   FA_X1 i_812 (.A(n_2060), .B(n_2091), .CI(n_2122), .CO(n_1625), .S(n_1624));
   FA_X1 i_813 (.A(n_2153), .B(n_2184), .CI(n_2215), .CO(n_1627), .S(n_1626));
   FA_X1 i_814 (.A(n_2246), .B(n_2277), .CI(n_2308), .CO(n_1629), .S(n_1628));
   FA_X1 i_815 (.A(n_2339), .B(n_1597), .CI(n_1595), .CO(n_1631), .S(n_1630));
   FA_X1 i_816 (.A(n_1593), .B(n_1591), .CI(n_1589), .CO(n_1633), .S(n_1632));
   FA_X1 i_817 (.A(n_1601), .B(n_1599), .CI(n_1628), .CO(n_1635), .S(n_1634));
   FA_X1 i_818 (.A(n_1626), .B(n_1624), .CI(n_1622), .CO(n_1637), .S(n_1636));
   FA_X1 i_819 (.A(n_1620), .B(n_1603), .CI(n_1632), .CO(n_1639), .S(n_1638));
   FA_X1 i_820 (.A(n_1630), .B(n_1607), .CI(n_1605), .CO(n_1641), .S(n_1640));
   FA_X1 i_821 (.A(n_1634), .B(n_1609), .CI(n_1611), .CO(n_1643), .S(n_1642));
   FA_X1 i_822 (.A(n_1636), .B(n_1638), .CI(n_1640), .CO(n_1645), .S(n_1644));
   FA_X1 i_823 (.A(n_1613), .B(n_1642), .CI(n_1615), .CO(n_1647), .S(n_1646));
   FA_X1 i_824 (.A(n_1644), .B(n_1617), .CI(n_1646), .CO(n_1649), .S(n_1648));
   FA_X1 i_825 (.A(n_1873), .B(n_1904), .CI(n_1935), .CO(n_1651), .S(n_1650));
   FA_X1 i_826 (.A(n_1966), .B(n_1997), .CI(n_2028), .CO(n_1653), .S(n_1652));
   FA_X1 i_827 (.A(n_2059), .B(n_2090), .CI(n_2121), .CO(n_1655), .S(n_1654));
   FA_X1 i_828 (.A(n_2152), .B(n_2183), .CI(n_2214), .CO(n_1657), .S(n_1656));
   FA_X1 i_829 (.A(n_2245), .B(n_2276), .CI(n_2307), .CO(n_1659), .S(n_1658));
   FA_X1 i_830 (.A(n_1629), .B(n_1627), .CI(n_1625), .CO(n_1661), .S(n_1660));
   FA_X1 i_831 (.A(n_1623), .B(n_1621), .CI(n_1633), .CO(n_1663), .S(n_1662));
   FA_X1 i_832 (.A(n_1631), .B(n_1658), .CI(n_1656), .CO(n_1665), .S(n_1664));
   FA_X1 i_833 (.A(n_1654), .B(n_1652), .CI(n_1650), .CO(n_1667), .S(n_1666));
   FA_X1 i_834 (.A(n_1662), .B(n_1660), .CI(n_1637), .CO(n_1669), .S(n_1668));
   FA_X1 i_835 (.A(n_1635), .B(n_1641), .CI(n_1639), .CO(n_1671), .S(n_1670));
   FA_X1 i_836 (.A(n_1666), .B(n_1664), .CI(n_1643), .CO(n_1673), .S(n_1672));
   FA_X1 i_837 (.A(n_1668), .B(n_1670), .CI(n_1645), .CO(n_1675), .S(n_1674));
   FA_X1 i_838 (.A(n_1672), .B(n_1647), .CI(n_1674), .CO(n_1677), .S(n_1676));
   FA_X1 i_839 (.A(n_1872), .B(n_1903), .CI(n_1934), .CO(n_1679), .S(n_1678));
   FA_X1 i_840 (.A(n_1965), .B(n_1996), .CI(n_2027), .CO(n_1681), .S(n_1680));
   FA_X1 i_841 (.A(n_2058), .B(n_2089), .CI(n_2120), .CO(n_1683), .S(n_1682));
   FA_X1 i_842 (.A(n_2151), .B(n_2182), .CI(n_2213), .CO(n_1685), .S(n_1684));
   FA_X1 i_843 (.A(n_2244), .B(n_2275), .CI(n_1659), .CO(n_1687), .S(n_1686));
   FA_X1 i_844 (.A(n_1657), .B(n_1655), .CI(n_1653), .CO(n_1689), .S(n_1688));
   FA_X1 i_845 (.A(n_1651), .B(n_1661), .CI(n_1686), .CO(n_1691), .S(n_1690));
   FA_X1 i_846 (.A(n_1684), .B(n_1682), .CI(n_1680), .CO(n_1693), .S(n_1692));
   FA_X1 i_847 (.A(n_1678), .B(n_1663), .CI(n_1688), .CO(n_1695), .S(n_1694));
   FA_X1 i_848 (.A(n_1667), .B(n_1665), .CI(n_1690), .CO(n_1697), .S(n_1696));
   FA_X1 i_849 (.A(n_1669), .B(n_1692), .CI(n_1694), .CO(n_1699), .S(n_1698));
   FA_X1 i_850 (.A(n_1671), .B(n_1696), .CI(n_1673), .CO(n_1701), .S(n_1700));
   FA_X1 i_851 (.A(n_1698), .B(n_1675), .CI(n_1700), .CO(n_1703), .S(n_1702));
   FA_X1 i_852 (.A(n_1871), .B(n_1902), .CI(n_1933), .CO(n_1705), .S(n_1704));
   FA_X1 i_853 (.A(n_1964), .B(n_1995), .CI(n_2026), .CO(n_1707), .S(n_1706));
   FA_X1 i_854 (.A(n_2057), .B(n_2088), .CI(n_2119), .CO(n_1709), .S(n_1708));
   FA_X1 i_855 (.A(n_2150), .B(n_2181), .CI(n_2212), .CO(n_1711), .S(n_1710));
   FA_X1 i_856 (.A(n_2243), .B(n_1685), .CI(n_1683), .CO(n_1713), .S(n_1712));
   FA_X1 i_857 (.A(n_1681), .B(n_1679), .CI(n_1689), .CO(n_1715), .S(n_1714));
   FA_X1 i_858 (.A(n_1687), .B(n_1710), .CI(n_1708), .CO(n_1717), .S(n_1716));
   FA_X1 i_859 (.A(n_1706), .B(n_1704), .CI(n_1714), .CO(n_1719), .S(n_1718));
   FA_X1 i_860 (.A(n_1712), .B(n_1693), .CI(n_1691), .CO(n_1721), .S(n_1720));
   FA_X1 i_861 (.A(n_1695), .B(n_1718), .CI(n_1716), .CO(n_1723), .S(n_1722));
   FA_X1 i_862 (.A(n_1697), .B(n_1720), .CI(n_1699), .CO(n_1725), .S(n_1724));
   FA_X1 i_863 (.A(n_1701), .B(n_1722), .CI(n_1724), .CO(n_1727), .S(n_1726));
   FA_X1 i_864 (.A(n_1870), .B(n_1901), .CI(n_1932), .CO(n_1729), .S(n_1728));
   FA_X1 i_865 (.A(n_1963), .B(n_1994), .CI(n_2025), .CO(n_1731), .S(n_1730));
   FA_X1 i_866 (.A(n_2056), .B(n_2087), .CI(n_2118), .CO(n_1733), .S(n_1732));
   FA_X1 i_867 (.A(n_2149), .B(n_2180), .CI(n_2211), .CO(n_1735), .S(n_1734));
   FA_X1 i_868 (.A(n_1711), .B(n_1709), .CI(n_1707), .CO(n_1737), .S(n_1736));
   FA_X1 i_869 (.A(n_1705), .B(n_1713), .CI(n_1734), .CO(n_1739), .S(n_1738));
   FA_X1 i_870 (.A(n_1732), .B(n_1730), .CI(n_1728), .CO(n_1741), .S(n_1740));
   FA_X1 i_871 (.A(n_1715), .B(n_1736), .CI(n_1717), .CO(n_1743), .S(n_1742));
   FA_X1 i_872 (.A(n_1738), .B(n_1721), .CI(n_1719), .CO(n_1745), .S(n_1744));
   FA_X1 i_873 (.A(n_1740), .B(n_1742), .CI(n_1723), .CO(n_1747), .S(n_1746));
   FA_X1 i_874 (.A(n_1744), .B(n_1725), .CI(n_1746), .CO(n_1749), .S(n_1748));
   FA_X1 i_875 (.A(n_1869), .B(n_1900), .CI(n_1931), .CO(n_1751), .S(n_1750));
   FA_X1 i_876 (.A(n_1962), .B(n_1993), .CI(n_2024), .CO(n_1753), .S(n_1752));
   FA_X1 i_877 (.A(n_2055), .B(n_2086), .CI(n_2117), .CO(n_1755), .S(n_1754));
   FA_X1 i_878 (.A(n_2148), .B(n_2179), .CI(n_1735), .CO(n_1757), .S(n_1756));
   FA_X1 i_879 (.A(n_1733), .B(n_1731), .CI(n_1729), .CO(n_1759), .S(n_1758));
   FA_X1 i_880 (.A(n_1737), .B(n_1756), .CI(n_1754), .CO(n_1761), .S(n_1760));
   FA_X1 i_881 (.A(n_1752), .B(n_1750), .CI(n_1758), .CO(n_1763), .S(n_1762));
   FA_X1 i_882 (.A(n_1741), .B(n_1739), .CI(n_1743), .CO(n_1765), .S(n_1764));
   FA_X1 i_883 (.A(n_1762), .B(n_1760), .CI(n_1745), .CO(n_1767), .S(n_1766));
   FA_X1 i_884 (.A(n_1764), .B(n_1747), .CI(n_1766), .CO(n_1769), .S(n_1768));
   FA_X1 i_885 (.A(n_1868), .B(n_1899), .CI(n_1930), .CO(n_1771), .S(n_1770));
   FA_X1 i_886 (.A(n_1961), .B(n_1992), .CI(n_2023), .CO(n_1773), .S(n_1772));
   FA_X1 i_887 (.A(n_2054), .B(n_2085), .CI(n_2116), .CO(n_1775), .S(n_1774));
   FA_X1 i_888 (.A(n_2147), .B(n_1755), .CI(n_1753), .CO(n_1777), .S(n_1776));
   FA_X1 i_889 (.A(n_1751), .B(n_1759), .CI(n_1757), .CO(n_1779), .S(n_1778));
   FA_X1 i_890 (.A(n_1774), .B(n_1772), .CI(n_1770), .CO(n_1781), .S(n_1780));
   FA_X1 i_891 (.A(n_1776), .B(n_1761), .CI(n_1778), .CO(n_1783), .S(n_1782));
   FA_X1 i_892 (.A(n_1763), .B(n_1780), .CI(n_1765), .CO(n_1785), .S(n_1784));
   FA_X1 i_893 (.A(n_1782), .B(n_1767), .CI(n_1784), .CO(n_1787), .S(n_1786));
   FA_X1 i_894 (.A(n_1867), .B(n_1898), .CI(n_1929), .CO(n_1789), .S(n_1788));
   FA_X1 i_895 (.A(n_1960), .B(n_1991), .CI(n_2022), .CO(n_1791), .S(n_1790));
   FA_X1 i_896 (.A(n_2053), .B(n_2084), .CI(n_2115), .CO(n_1793), .S(n_1792));
   FA_X1 i_897 (.A(n_1775), .B(n_1773), .CI(n_1771), .CO(n_1795), .S(n_1794));
   FA_X1 i_898 (.A(n_1777), .B(n_1792), .CI(n_1790), .CO(n_1797), .S(n_1796));
   FA_X1 i_899 (.A(n_1788), .B(n_1779), .CI(n_1794), .CO(n_1799), .S(n_1798));
   FA_X1 i_900 (.A(n_1781), .B(n_1796), .CI(n_1798), .CO(n_1801), .S(n_1800));
   FA_X1 i_901 (.A(n_1783), .B(n_1785), .CI(n_1800), .CO(n_1803), .S(n_1802));
   FA_X1 i_902 (.A(n_1866), .B(n_1897), .CI(n_1928), .CO(n_1805), .S(n_1804));
   FA_X1 i_903 (.A(n_1959), .B(n_1990), .CI(n_2021), .CO(n_1807), .S(n_1806));
   FA_X1 i_904 (.A(n_2052), .B(n_2083), .CI(n_1793), .CO(n_1809), .S(n_1808));
   FA_X1 i_905 (.A(n_1791), .B(n_1789), .CI(n_1795), .CO(n_1811), .S(n_1810));
   FA_X1 i_906 (.A(n_1808), .B(n_1806), .CI(n_1804), .CO(n_1813), .S(n_1812));
   FA_X1 i_907 (.A(n_1810), .B(n_1797), .CI(n_1799), .CO(n_1815), .S(n_1814));
   FA_X1 i_908 (.A(n_1812), .B(n_1814), .CI(n_1801), .CO(n_1817), .S(n_1816));
   FA_X1 i_909 (.A(n_1865), .B(n_1896), .CI(n_1927), .CO(n_1819), .S(n_1818));
   FA_X1 i_910 (.A(n_1958), .B(n_1989), .CI(n_2020), .CO(n_1821), .S(n_1820));
   FA_X1 i_911 (.A(n_2051), .B(n_1807), .CI(n_1805), .CO(n_1823), .S(n_1822));
   FA_X1 i_912 (.A(n_1809), .B(n_1820), .CI(n_1818), .CO(n_1825), .S(n_1824));
   FA_X1 i_913 (.A(n_1811), .B(n_1822), .CI(n_1813), .CO(n_1827), .S(n_1826));
   FA_X1 i_914 (.A(n_1824), .B(n_1815), .CI(n_1826), .CO(n_1829), .S(n_1828));
   FA_X1 i_915 (.A(n_1864), .B(n_1895), .CI(n_1926), .CO(n_1831), .S(n_1830));
   FA_X1 i_916 (.A(n_1957), .B(n_1988), .CI(n_2019), .CO(n_1833), .S(n_1832));
   FA_X1 i_917 (.A(n_1821), .B(n_1819), .CI(n_1823), .CO(n_1835), .S(n_1834));
   FA_X1 i_918 (.A(n_1832), .B(n_1830), .CI(n_1834), .CO(n_1837), .S(n_1836));
   FA_X1 i_919 (.A(n_1825), .B(n_1827), .CI(n_1836), .CO(n_1839), .S(n_1838));
   FA_X1 i_920 (.A(n_1863), .B(n_1894), .CI(n_1925), .CO(n_1841), .S(n_1840));
   FA_X1 i_921 (.A(n_1956), .B(n_1987), .CI(n_1833), .CO(n_1843), .S(n_1842));
   FA_X1 i_922 (.A(n_1831), .B(n_1842), .CI(n_1840), .CO(n_1845), .S(n_1844));
   FA_X1 i_923 (.A(n_1835), .B(n_1837), .CI(n_1844), .CO(n_1847), .S(n_1846));
   FA_X1 i_924 (.A(n_1862), .B(n_1893), .CI(n_1924), .CO(n_1849), .S(n_1848));
   FA_X1 i_925 (.A(n_1955), .B(n_1841), .CI(n_1843), .CO(n_1851), .S(n_1850));
   FA_X1 i_926 (.A(n_1848), .B(n_1850), .CI(n_1845), .CO(n_1853), .S(n_1852));
   FA_X1 i_927 (.A(n_1861), .B(n_1892), .CI(n_1923), .CO(n_1855), .S(n_1854));
   FA_X1 i_928 (.A(n_1849), .B(n_1854), .CI(n_1851), .CO(n_1857), .S(n_1856));
   FA_X1 i_929 (.A(n_1860), .B(n_1891), .CI(n_1855), .CO(n_1859), .S(n_1858));
   NOR2_X1 i_930 (.A1(n_3309), .A2(n_3276), .ZN(n_1860));
   NOR2_X1 i_931 (.A1(n_3309), .A2(n_3275), .ZN(n_1861));
   NOR2_X1 i_932 (.A1(n_3309), .A2(n_3274), .ZN(n_1862));
   NOR2_X1 i_933 (.A1(n_3309), .A2(n_3273), .ZN(n_1863));
   NOR2_X1 i_934 (.A1(n_3309), .A2(n_3272), .ZN(n_1864));
   NOR2_X1 i_935 (.A1(n_3309), .A2(n_3271), .ZN(n_1865));
   NOR2_X1 i_936 (.A1(n_3309), .A2(n_3270), .ZN(n_1866));
   NOR2_X1 i_937 (.A1(n_3309), .A2(n_3269), .ZN(n_1867));
   NOR2_X1 i_938 (.A1(n_3309), .A2(n_3268), .ZN(n_1868));
   NOR2_X1 i_939 (.A1(n_3309), .A2(n_3267), .ZN(n_1869));
   NOR2_X1 i_940 (.A1(n_3309), .A2(n_3266), .ZN(n_1870));
   NOR2_X1 i_941 (.A1(n_3309), .A2(n_3265), .ZN(n_1871));
   NOR2_X1 i_942 (.A1(n_3309), .A2(n_3264), .ZN(n_1872));
   NOR2_X1 i_943 (.A1(n_3309), .A2(n_3263), .ZN(n_1873));
   NOR2_X1 i_944 (.A1(n_3309), .A2(n_3262), .ZN(n_1874));
   NOR2_X1 i_945 (.A1(n_3309), .A2(n_3261), .ZN(n_1875));
   NOR2_X1 i_946 (.A1(n_3309), .A2(n_3260), .ZN(n_1876));
   NOR2_X1 i_947 (.A1(n_3309), .A2(n_3259), .ZN(n_1877));
   NOR2_X1 i_948 (.A1(n_3309), .A2(n_3258), .ZN(n_1878));
   NOR2_X1 i_949 (.A1(n_3309), .A2(n_3257), .ZN(n_1879));
   NOR2_X1 i_950 (.A1(n_3309), .A2(n_3256), .ZN(n_1880));
   NOR2_X1 i_951 (.A1(n_3309), .A2(n_3255), .ZN(n_1881));
   NOR2_X1 i_952 (.A1(n_3309), .A2(n_3254), .ZN(n_1882));
   NOR2_X1 i_953 (.A1(n_3309), .A2(n_3253), .ZN(n_1883));
   NOR2_X1 i_954 (.A1(n_3309), .A2(n_3252), .ZN(n_1884));
   NOR2_X1 i_955 (.A1(n_3309), .A2(n_3251), .ZN(n_1885));
   NOR2_X1 i_956 (.A1(n_3309), .A2(n_3250), .ZN(n_1886));
   NOR2_X1 i_957 (.A1(n_3309), .A2(n_3249), .ZN(n_1887));
   NOR2_X1 i_958 (.A1(n_3309), .A2(n_3248), .ZN(n_1888));
   NOR2_X1 i_959 (.A1(n_3309), .A2(n_3247), .ZN(n_1889));
   NOR2_X1 i_960 (.A1(n_3309), .A2(n_3246), .ZN(n_1890));
   NOR2_X1 i_961 (.A1(n_3308), .A2(n_3277), .ZN(n_1891));
   NOR2_X1 i_962 (.A1(n_3308), .A2(n_3276), .ZN(n_1892));
   NOR2_X1 i_963 (.A1(n_3308), .A2(n_3275), .ZN(n_1893));
   NOR2_X1 i_964 (.A1(n_3308), .A2(n_3274), .ZN(n_1894));
   NOR2_X1 i_965 (.A1(n_3308), .A2(n_3273), .ZN(n_1895));
   NOR2_X1 i_966 (.A1(n_3308), .A2(n_3272), .ZN(n_1896));
   NOR2_X1 i_967 (.A1(n_3308), .A2(n_3271), .ZN(n_1897));
   NOR2_X1 i_968 (.A1(n_3308), .A2(n_3270), .ZN(n_1898));
   NOR2_X1 i_969 (.A1(n_3308), .A2(n_3269), .ZN(n_1899));
   NOR2_X1 i_970 (.A1(n_3308), .A2(n_3268), .ZN(n_1900));
   NOR2_X1 i_971 (.A1(n_3308), .A2(n_3267), .ZN(n_1901));
   NOR2_X1 i_972 (.A1(n_3308), .A2(n_3266), .ZN(n_1902));
   NOR2_X1 i_973 (.A1(n_3308), .A2(n_3265), .ZN(n_1903));
   NOR2_X1 i_974 (.A1(n_3308), .A2(n_3264), .ZN(n_1904));
   NOR2_X1 i_975 (.A1(n_3308), .A2(n_3263), .ZN(n_1905));
   NOR2_X1 i_976 (.A1(n_3308), .A2(n_3262), .ZN(n_1906));
   NOR2_X1 i_977 (.A1(n_3308), .A2(n_3261), .ZN(n_1907));
   NOR2_X1 i_978 (.A1(n_3308), .A2(n_3260), .ZN(n_1908));
   NOR2_X1 i_979 (.A1(n_3308), .A2(n_3259), .ZN(n_1909));
   NOR2_X1 i_980 (.A1(n_3308), .A2(n_3258), .ZN(n_1910));
   NOR2_X1 i_981 (.A1(n_3308), .A2(n_3257), .ZN(n_1911));
   NOR2_X1 i_982 (.A1(n_3308), .A2(n_3256), .ZN(n_1912));
   NOR2_X1 i_983 (.A1(n_3308), .A2(n_3255), .ZN(n_1913));
   NOR2_X1 i_984 (.A1(n_3308), .A2(n_3254), .ZN(n_1914));
   NOR2_X1 i_985 (.A1(n_3308), .A2(n_3253), .ZN(n_1915));
   NOR2_X1 i_986 (.A1(n_3308), .A2(n_3252), .ZN(n_1916));
   NOR2_X1 i_987 (.A1(n_3308), .A2(n_3251), .ZN(n_1917));
   NOR2_X1 i_988 (.A1(n_3308), .A2(n_3250), .ZN(n_1918));
   NOR2_X1 i_989 (.A1(n_3308), .A2(n_3249), .ZN(n_1919));
   NOR2_X1 i_990 (.A1(n_3308), .A2(n_3248), .ZN(n_1920));
   NOR2_X1 i_991 (.A1(n_3308), .A2(n_3247), .ZN(n_1921));
   NOR2_X1 i_992 (.A1(n_3308), .A2(n_3246), .ZN(n_1922));
   NOR2_X1 i_993 (.A1(n_3307), .A2(n_3277), .ZN(n_1923));
   NOR2_X1 i_994 (.A1(n_3307), .A2(n_3276), .ZN(n_1924));
   NOR2_X1 i_995 (.A1(n_3307), .A2(n_3275), .ZN(n_1925));
   NOR2_X1 i_996 (.A1(n_3307), .A2(n_3274), .ZN(n_1926));
   NOR2_X1 i_997 (.A1(n_3307), .A2(n_3273), .ZN(n_1927));
   NOR2_X1 i_998 (.A1(n_3307), .A2(n_3272), .ZN(n_1928));
   NOR2_X1 i_999 (.A1(n_3307), .A2(n_3271), .ZN(n_1929));
   NOR2_X1 i_1000 (.A1(n_3307), .A2(n_3270), .ZN(n_1930));
   NOR2_X1 i_1001 (.A1(n_3307), .A2(n_3269), .ZN(n_1931));
   NOR2_X1 i_1002 (.A1(n_3307), .A2(n_3268), .ZN(n_1932));
   NOR2_X1 i_1003 (.A1(n_3307), .A2(n_3267), .ZN(n_1933));
   NOR2_X1 i_1004 (.A1(n_3307), .A2(n_3266), .ZN(n_1934));
   NOR2_X1 i_1005 (.A1(n_3307), .A2(n_3265), .ZN(n_1935));
   NOR2_X1 i_1006 (.A1(n_3307), .A2(n_3264), .ZN(n_1936));
   NOR2_X1 i_1007 (.A1(n_3307), .A2(n_3263), .ZN(n_1937));
   NOR2_X1 i_1008 (.A1(n_3307), .A2(n_3262), .ZN(n_1938));
   NOR2_X1 i_1009 (.A1(n_3307), .A2(n_3261), .ZN(n_1939));
   NOR2_X1 i_1010 (.A1(n_3307), .A2(n_3260), .ZN(n_1940));
   NOR2_X1 i_1011 (.A1(n_3307), .A2(n_3259), .ZN(n_1941));
   NOR2_X1 i_1012 (.A1(n_3307), .A2(n_3258), .ZN(n_1942));
   NOR2_X1 i_1013 (.A1(n_3307), .A2(n_3257), .ZN(n_1943));
   NOR2_X1 i_1014 (.A1(n_3307), .A2(n_3256), .ZN(n_1944));
   NOR2_X1 i_1015 (.A1(n_3307), .A2(n_3255), .ZN(n_1945));
   NOR2_X1 i_1016 (.A1(n_3307), .A2(n_3254), .ZN(n_1946));
   NOR2_X1 i_1017 (.A1(n_3307), .A2(n_3253), .ZN(n_1947));
   NOR2_X1 i_1018 (.A1(n_3307), .A2(n_3252), .ZN(n_1948));
   NOR2_X1 i_1019 (.A1(n_3307), .A2(n_3251), .ZN(n_1949));
   NOR2_X1 i_1020 (.A1(n_3307), .A2(n_3250), .ZN(n_1950));
   NOR2_X1 i_1021 (.A1(n_3307), .A2(n_3249), .ZN(n_1951));
   NOR2_X1 i_1022 (.A1(n_3307), .A2(n_3248), .ZN(n_1952));
   NOR2_X1 i_1023 (.A1(n_3307), .A2(n_3247), .ZN(n_1953));
   NOR2_X1 i_1024 (.A1(n_3307), .A2(n_3246), .ZN(n_1954));
   NOR2_X1 i_1025 (.A1(n_3306), .A2(n_3277), .ZN(n_1955));
   NOR2_X1 i_1026 (.A1(n_3306), .A2(n_3276), .ZN(n_1956));
   NOR2_X1 i_1027 (.A1(n_3306), .A2(n_3275), .ZN(n_1957));
   NOR2_X1 i_1028 (.A1(n_3306), .A2(n_3274), .ZN(n_1958));
   NOR2_X1 i_1029 (.A1(n_3306), .A2(n_3273), .ZN(n_1959));
   NOR2_X1 i_1030 (.A1(n_3306), .A2(n_3272), .ZN(n_1960));
   NOR2_X1 i_1031 (.A1(n_3306), .A2(n_3271), .ZN(n_1961));
   NOR2_X1 i_1032 (.A1(n_3306), .A2(n_3270), .ZN(n_1962));
   NOR2_X1 i_1033 (.A1(n_3306), .A2(n_3269), .ZN(n_1963));
   NOR2_X1 i_1034 (.A1(n_3306), .A2(n_3268), .ZN(n_1964));
   NOR2_X1 i_1035 (.A1(n_3306), .A2(n_3267), .ZN(n_1965));
   NOR2_X1 i_1036 (.A1(n_3306), .A2(n_3266), .ZN(n_1966));
   NOR2_X1 i_1037 (.A1(n_3306), .A2(n_3265), .ZN(n_1967));
   NOR2_X1 i_1038 (.A1(n_3306), .A2(n_3264), .ZN(n_1968));
   NOR2_X1 i_1039 (.A1(n_3306), .A2(n_3263), .ZN(n_1969));
   NOR2_X1 i_1040 (.A1(n_3306), .A2(n_3262), .ZN(n_1970));
   NOR2_X1 i_1041 (.A1(n_3306), .A2(n_3261), .ZN(n_1971));
   NOR2_X1 i_1042 (.A1(n_3306), .A2(n_3260), .ZN(n_1972));
   NOR2_X1 i_1043 (.A1(n_3306), .A2(n_3259), .ZN(n_1973));
   NOR2_X1 i_1044 (.A1(n_3306), .A2(n_3258), .ZN(n_1974));
   NOR2_X1 i_1045 (.A1(n_3306), .A2(n_3257), .ZN(n_1975));
   NOR2_X1 i_1046 (.A1(n_3306), .A2(n_3256), .ZN(n_1976));
   NOR2_X1 i_1047 (.A1(n_3306), .A2(n_3255), .ZN(n_1977));
   NOR2_X1 i_1048 (.A1(n_3306), .A2(n_3254), .ZN(n_1978));
   NOR2_X1 i_1049 (.A1(n_3306), .A2(n_3253), .ZN(n_1979));
   NOR2_X1 i_1050 (.A1(n_3306), .A2(n_3252), .ZN(n_1980));
   NOR2_X1 i_1051 (.A1(n_3306), .A2(n_3251), .ZN(n_1981));
   NOR2_X1 i_1052 (.A1(n_3306), .A2(n_3250), .ZN(n_1982));
   NOR2_X1 i_1053 (.A1(n_3306), .A2(n_3249), .ZN(n_1983));
   NOR2_X1 i_1054 (.A1(n_3306), .A2(n_3248), .ZN(n_1984));
   NOR2_X1 i_1055 (.A1(n_3306), .A2(n_3247), .ZN(n_1985));
   NOR2_X1 i_1056 (.A1(n_3306), .A2(n_3246), .ZN(n_1986));
   NOR2_X1 i_1057 (.A1(n_3305), .A2(n_3277), .ZN(n_1987));
   NOR2_X1 i_1058 (.A1(n_3305), .A2(n_3276), .ZN(n_1988));
   NOR2_X1 i_1059 (.A1(n_3305), .A2(n_3275), .ZN(n_1989));
   NOR2_X1 i_1060 (.A1(n_3305), .A2(n_3274), .ZN(n_1990));
   NOR2_X1 i_1061 (.A1(n_3305), .A2(n_3273), .ZN(n_1991));
   NOR2_X1 i_1062 (.A1(n_3305), .A2(n_3272), .ZN(n_1992));
   NOR2_X1 i_1063 (.A1(n_3305), .A2(n_3271), .ZN(n_1993));
   NOR2_X1 i_1064 (.A1(n_3305), .A2(n_3270), .ZN(n_1994));
   NOR2_X1 i_1065 (.A1(n_3305), .A2(n_3269), .ZN(n_1995));
   NOR2_X1 i_1066 (.A1(n_3305), .A2(n_3268), .ZN(n_1996));
   NOR2_X1 i_1067 (.A1(n_3305), .A2(n_3267), .ZN(n_1997));
   NOR2_X1 i_1068 (.A1(n_3305), .A2(n_3266), .ZN(n_1998));
   NOR2_X1 i_1069 (.A1(n_3305), .A2(n_3265), .ZN(n_1999));
   NOR2_X1 i_1070 (.A1(n_3305), .A2(n_3264), .ZN(n_2000));
   NOR2_X1 i_1071 (.A1(n_3305), .A2(n_3263), .ZN(n_2001));
   NOR2_X1 i_1072 (.A1(n_3305), .A2(n_3262), .ZN(n_2002));
   NOR2_X1 i_1073 (.A1(n_3305), .A2(n_3261), .ZN(n_2003));
   NOR2_X1 i_1074 (.A1(n_3305), .A2(n_3260), .ZN(n_2004));
   NOR2_X1 i_1075 (.A1(n_3305), .A2(n_3259), .ZN(n_2005));
   NOR2_X1 i_1076 (.A1(n_3305), .A2(n_3258), .ZN(n_2006));
   NOR2_X1 i_1077 (.A1(n_3305), .A2(n_3257), .ZN(n_2007));
   NOR2_X1 i_1078 (.A1(n_3305), .A2(n_3256), .ZN(n_2008));
   NOR2_X1 i_1079 (.A1(n_3305), .A2(n_3255), .ZN(n_2009));
   NOR2_X1 i_1080 (.A1(n_3305), .A2(n_3254), .ZN(n_2010));
   NOR2_X1 i_1081 (.A1(n_3305), .A2(n_3253), .ZN(n_2011));
   NOR2_X1 i_1082 (.A1(n_3305), .A2(n_3252), .ZN(n_2012));
   NOR2_X1 i_1083 (.A1(n_3305), .A2(n_3251), .ZN(n_2013));
   NOR2_X1 i_1084 (.A1(n_3305), .A2(n_3250), .ZN(n_2014));
   NOR2_X1 i_1085 (.A1(n_3305), .A2(n_3249), .ZN(n_2015));
   NOR2_X1 i_1086 (.A1(n_3305), .A2(n_3248), .ZN(n_2016));
   NOR2_X1 i_1087 (.A1(n_3305), .A2(n_3247), .ZN(n_2017));
   NOR2_X1 i_1088 (.A1(n_3305), .A2(n_3246), .ZN(n_2018));
   NOR2_X1 i_1089 (.A1(n_3304), .A2(n_3277), .ZN(n_2019));
   NOR2_X1 i_1090 (.A1(n_3304), .A2(n_3276), .ZN(n_2020));
   NOR2_X1 i_1091 (.A1(n_3304), .A2(n_3275), .ZN(n_2021));
   NOR2_X1 i_1092 (.A1(n_3304), .A2(n_3274), .ZN(n_2022));
   NOR2_X1 i_1093 (.A1(n_3304), .A2(n_3273), .ZN(n_2023));
   NOR2_X1 i_1094 (.A1(n_3304), .A2(n_3272), .ZN(n_2024));
   NOR2_X1 i_1095 (.A1(n_3304), .A2(n_3271), .ZN(n_2025));
   NOR2_X1 i_1096 (.A1(n_3304), .A2(n_3270), .ZN(n_2026));
   NOR2_X1 i_1097 (.A1(n_3304), .A2(n_3269), .ZN(n_2027));
   NOR2_X1 i_1098 (.A1(n_3304), .A2(n_3268), .ZN(n_2028));
   NOR2_X1 i_1099 (.A1(n_3304), .A2(n_3267), .ZN(n_2029));
   NOR2_X1 i_1100 (.A1(n_3304), .A2(n_3266), .ZN(n_2030));
   NOR2_X1 i_1101 (.A1(n_3304), .A2(n_3265), .ZN(n_2031));
   NOR2_X1 i_1102 (.A1(n_3304), .A2(n_3264), .ZN(n_2032));
   NOR2_X1 i_1103 (.A1(n_3304), .A2(n_3263), .ZN(n_2033));
   NOR2_X1 i_1104 (.A1(n_3304), .A2(n_3262), .ZN(n_2034));
   NOR2_X1 i_1105 (.A1(n_3304), .A2(n_3261), .ZN(n_2035));
   NOR2_X1 i_1106 (.A1(n_3304), .A2(n_3260), .ZN(n_2036));
   NOR2_X1 i_1107 (.A1(n_3304), .A2(n_3259), .ZN(n_2037));
   NOR2_X1 i_1108 (.A1(n_3304), .A2(n_3258), .ZN(n_2038));
   NOR2_X1 i_1109 (.A1(n_3304), .A2(n_3257), .ZN(n_2039));
   NOR2_X1 i_1110 (.A1(n_3304), .A2(n_3256), .ZN(n_2040));
   NOR2_X1 i_1111 (.A1(n_3304), .A2(n_3255), .ZN(n_2041));
   NOR2_X1 i_1112 (.A1(n_3304), .A2(n_3254), .ZN(n_2042));
   NOR2_X1 i_1113 (.A1(n_3304), .A2(n_3253), .ZN(n_2043));
   NOR2_X1 i_1114 (.A1(n_3304), .A2(n_3252), .ZN(n_2044));
   NOR2_X1 i_1115 (.A1(n_3304), .A2(n_3251), .ZN(n_2045));
   NOR2_X1 i_1116 (.A1(n_3304), .A2(n_3250), .ZN(n_2046));
   NOR2_X1 i_1117 (.A1(n_3304), .A2(n_3249), .ZN(n_2047));
   NOR2_X1 i_1118 (.A1(n_3304), .A2(n_3248), .ZN(n_2048));
   NOR2_X1 i_1119 (.A1(n_3304), .A2(n_3247), .ZN(n_2049));
   NOR2_X1 i_1120 (.A1(n_3304), .A2(n_3246), .ZN(n_2050));
   NOR2_X1 i_1121 (.A1(n_3303), .A2(n_3277), .ZN(n_2051));
   NOR2_X1 i_1122 (.A1(n_3303), .A2(n_3276), .ZN(n_2052));
   NOR2_X1 i_1123 (.A1(n_3303), .A2(n_3275), .ZN(n_2053));
   NOR2_X1 i_1124 (.A1(n_3303), .A2(n_3274), .ZN(n_2054));
   NOR2_X1 i_1125 (.A1(n_3303), .A2(n_3273), .ZN(n_2055));
   NOR2_X1 i_1126 (.A1(n_3303), .A2(n_3272), .ZN(n_2056));
   NOR2_X1 i_1127 (.A1(n_3303), .A2(n_3271), .ZN(n_2057));
   NOR2_X1 i_1128 (.A1(n_3303), .A2(n_3270), .ZN(n_2058));
   NOR2_X1 i_1129 (.A1(n_3303), .A2(n_3269), .ZN(n_2059));
   NOR2_X1 i_1130 (.A1(n_3303), .A2(n_3268), .ZN(n_2060));
   NOR2_X1 i_1131 (.A1(n_3303), .A2(n_3267), .ZN(n_2061));
   NOR2_X1 i_1132 (.A1(n_3303), .A2(n_3266), .ZN(n_2062));
   NOR2_X1 i_1133 (.A1(n_3303), .A2(n_3265), .ZN(n_2063));
   NOR2_X1 i_1134 (.A1(n_3303), .A2(n_3264), .ZN(n_2064));
   NOR2_X1 i_1135 (.A1(n_3303), .A2(n_3263), .ZN(n_2065));
   NOR2_X1 i_1136 (.A1(n_3303), .A2(n_3262), .ZN(n_2066));
   NOR2_X1 i_1137 (.A1(n_3303), .A2(n_3261), .ZN(n_2067));
   NOR2_X1 i_1138 (.A1(n_3303), .A2(n_3260), .ZN(n_2068));
   NOR2_X1 i_1139 (.A1(n_3303), .A2(n_3259), .ZN(n_2069));
   NOR2_X1 i_1140 (.A1(n_3303), .A2(n_3258), .ZN(n_2070));
   NOR2_X1 i_1141 (.A1(n_3303), .A2(n_3257), .ZN(n_2071));
   NOR2_X1 i_1142 (.A1(n_3303), .A2(n_3256), .ZN(n_2072));
   NOR2_X1 i_1143 (.A1(n_3303), .A2(n_3255), .ZN(n_2073));
   NOR2_X1 i_1144 (.A1(n_3303), .A2(n_3254), .ZN(n_2074));
   NOR2_X1 i_1145 (.A1(n_3303), .A2(n_3253), .ZN(n_2075));
   NOR2_X1 i_1146 (.A1(n_3303), .A2(n_3252), .ZN(n_2076));
   NOR2_X1 i_1147 (.A1(n_3303), .A2(n_3251), .ZN(n_2077));
   NOR2_X1 i_1148 (.A1(n_3303), .A2(n_3250), .ZN(n_2078));
   NOR2_X1 i_1149 (.A1(n_3303), .A2(n_3249), .ZN(n_2079));
   NOR2_X1 i_1150 (.A1(n_3303), .A2(n_3248), .ZN(n_2080));
   NOR2_X1 i_1151 (.A1(n_3303), .A2(n_3247), .ZN(n_2081));
   NOR2_X1 i_1152 (.A1(n_3303), .A2(n_3246), .ZN(n_2082));
   NOR2_X1 i_1153 (.A1(n_3302), .A2(n_3277), .ZN(n_2083));
   NOR2_X1 i_1154 (.A1(n_3302), .A2(n_3276), .ZN(n_2084));
   NOR2_X1 i_1155 (.A1(n_3302), .A2(n_3275), .ZN(n_2085));
   NOR2_X1 i_1156 (.A1(n_3302), .A2(n_3274), .ZN(n_2086));
   NOR2_X1 i_1157 (.A1(n_3302), .A2(n_3273), .ZN(n_2087));
   NOR2_X1 i_1158 (.A1(n_3302), .A2(n_3272), .ZN(n_2088));
   NOR2_X1 i_1159 (.A1(n_3302), .A2(n_3271), .ZN(n_2089));
   NOR2_X1 i_1160 (.A1(n_3302), .A2(n_3270), .ZN(n_2090));
   NOR2_X1 i_1161 (.A1(n_3302), .A2(n_3269), .ZN(n_2091));
   NOR2_X1 i_1162 (.A1(n_3302), .A2(n_3268), .ZN(n_2092));
   NOR2_X1 i_1163 (.A1(n_3302), .A2(n_3267), .ZN(n_2093));
   NOR2_X1 i_1164 (.A1(n_3302), .A2(n_3266), .ZN(n_2094));
   NOR2_X1 i_1165 (.A1(n_3302), .A2(n_3265), .ZN(n_2095));
   NOR2_X1 i_1166 (.A1(n_3302), .A2(n_3264), .ZN(n_2096));
   NOR2_X1 i_1167 (.A1(n_3302), .A2(n_3263), .ZN(n_2097));
   NOR2_X1 i_1168 (.A1(n_3302), .A2(n_3262), .ZN(n_2098));
   NOR2_X1 i_1169 (.A1(n_3302), .A2(n_3261), .ZN(n_2099));
   NOR2_X1 i_1170 (.A1(n_3302), .A2(n_3260), .ZN(n_2100));
   NOR2_X1 i_1171 (.A1(n_3302), .A2(n_3259), .ZN(n_2101));
   NOR2_X1 i_1172 (.A1(n_3302), .A2(n_3258), .ZN(n_2102));
   NOR2_X1 i_1173 (.A1(n_3302), .A2(n_3257), .ZN(n_2103));
   NOR2_X1 i_1174 (.A1(n_3302), .A2(n_3256), .ZN(n_2104));
   NOR2_X1 i_1175 (.A1(n_3302), .A2(n_3255), .ZN(n_2105));
   NOR2_X1 i_1176 (.A1(n_3302), .A2(n_3254), .ZN(n_2106));
   NOR2_X1 i_1177 (.A1(n_3302), .A2(n_3253), .ZN(n_2107));
   NOR2_X1 i_1178 (.A1(n_3302), .A2(n_3252), .ZN(n_2108));
   NOR2_X1 i_1179 (.A1(n_3302), .A2(n_3251), .ZN(n_2109));
   NOR2_X1 i_1180 (.A1(n_3302), .A2(n_3250), .ZN(n_2110));
   NOR2_X1 i_1181 (.A1(n_3302), .A2(n_3249), .ZN(n_2111));
   NOR2_X1 i_1182 (.A1(n_3302), .A2(n_3248), .ZN(n_2112));
   NOR2_X1 i_1183 (.A1(n_3302), .A2(n_3247), .ZN(n_2113));
   NOR2_X1 i_1184 (.A1(n_3302), .A2(n_3246), .ZN(n_2114));
   NOR2_X1 i_1185 (.A1(n_3301), .A2(n_3277), .ZN(n_2115));
   NOR2_X1 i_1186 (.A1(n_3301), .A2(n_3276), .ZN(n_2116));
   NOR2_X1 i_1187 (.A1(n_3301), .A2(n_3275), .ZN(n_2117));
   NOR2_X1 i_1188 (.A1(n_3301), .A2(n_3274), .ZN(n_2118));
   NOR2_X1 i_1189 (.A1(n_3301), .A2(n_3273), .ZN(n_2119));
   NOR2_X1 i_1190 (.A1(n_3301), .A2(n_3272), .ZN(n_2120));
   NOR2_X1 i_1191 (.A1(n_3301), .A2(n_3271), .ZN(n_2121));
   NOR2_X1 i_1192 (.A1(n_3301), .A2(n_3270), .ZN(n_2122));
   NOR2_X1 i_1193 (.A1(n_3301), .A2(n_3269), .ZN(n_2123));
   NOR2_X1 i_1194 (.A1(n_3301), .A2(n_3268), .ZN(n_2124));
   NOR2_X1 i_1195 (.A1(n_3301), .A2(n_3267), .ZN(n_2125));
   NOR2_X1 i_1196 (.A1(n_3301), .A2(n_3266), .ZN(n_2126));
   NOR2_X1 i_1197 (.A1(n_3301), .A2(n_3265), .ZN(n_2127));
   NOR2_X1 i_1198 (.A1(n_3301), .A2(n_3264), .ZN(n_2128));
   NOR2_X1 i_1199 (.A1(n_3301), .A2(n_3263), .ZN(n_2129));
   NOR2_X1 i_1200 (.A1(n_3301), .A2(n_3262), .ZN(n_2130));
   NOR2_X1 i_1201 (.A1(n_3301), .A2(n_3261), .ZN(n_2131));
   NOR2_X1 i_1202 (.A1(n_3301), .A2(n_3260), .ZN(n_2132));
   NOR2_X1 i_1203 (.A1(n_3301), .A2(n_3259), .ZN(n_2133));
   NOR2_X1 i_1204 (.A1(n_3301), .A2(n_3258), .ZN(n_2134));
   NOR2_X1 i_1205 (.A1(n_3301), .A2(n_3257), .ZN(n_2135));
   NOR2_X1 i_1206 (.A1(n_3301), .A2(n_3256), .ZN(n_2136));
   NOR2_X1 i_1207 (.A1(n_3301), .A2(n_3255), .ZN(n_2137));
   NOR2_X1 i_1208 (.A1(n_3301), .A2(n_3254), .ZN(n_2138));
   NOR2_X1 i_1209 (.A1(n_3301), .A2(n_3253), .ZN(n_2139));
   NOR2_X1 i_1210 (.A1(n_3301), .A2(n_3252), .ZN(n_2140));
   NOR2_X1 i_1211 (.A1(n_3301), .A2(n_3251), .ZN(n_2141));
   NOR2_X1 i_1212 (.A1(n_3301), .A2(n_3250), .ZN(n_2142));
   NOR2_X1 i_1213 (.A1(n_3301), .A2(n_3249), .ZN(n_2143));
   NOR2_X1 i_1214 (.A1(n_3301), .A2(n_3248), .ZN(n_2144));
   NOR2_X1 i_1215 (.A1(n_3301), .A2(n_3247), .ZN(n_2145));
   NOR2_X1 i_1216 (.A1(n_3301), .A2(n_3246), .ZN(n_2146));
   NOR2_X1 i_1217 (.A1(n_3300), .A2(n_3277), .ZN(n_2147));
   NOR2_X1 i_1218 (.A1(n_3300), .A2(n_3276), .ZN(n_2148));
   NOR2_X1 i_1219 (.A1(n_3300), .A2(n_3275), .ZN(n_2149));
   NOR2_X1 i_1220 (.A1(n_3300), .A2(n_3274), .ZN(n_2150));
   NOR2_X1 i_1221 (.A1(n_3300), .A2(n_3273), .ZN(n_2151));
   NOR2_X1 i_1222 (.A1(n_3300), .A2(n_3272), .ZN(n_2152));
   NOR2_X1 i_1223 (.A1(n_3300), .A2(n_3271), .ZN(n_2153));
   NOR2_X1 i_1224 (.A1(n_3300), .A2(n_3270), .ZN(n_2154));
   NOR2_X1 i_1225 (.A1(n_3300), .A2(n_3269), .ZN(n_2155));
   NOR2_X1 i_1226 (.A1(n_3300), .A2(n_3268), .ZN(n_2156));
   NOR2_X1 i_1227 (.A1(n_3300), .A2(n_3267), .ZN(n_2157));
   NOR2_X1 i_1228 (.A1(n_3300), .A2(n_3266), .ZN(n_2158));
   NOR2_X1 i_1229 (.A1(n_3300), .A2(n_3265), .ZN(n_2159));
   NOR2_X1 i_1230 (.A1(n_3300), .A2(n_3264), .ZN(n_2160));
   NOR2_X1 i_1231 (.A1(n_3300), .A2(n_3263), .ZN(n_2161));
   NOR2_X1 i_1232 (.A1(n_3300), .A2(n_3262), .ZN(n_2162));
   NOR2_X1 i_1233 (.A1(n_3300), .A2(n_3261), .ZN(n_2163));
   NOR2_X1 i_1234 (.A1(n_3300), .A2(n_3260), .ZN(n_2164));
   NOR2_X1 i_1235 (.A1(n_3300), .A2(n_3259), .ZN(n_2165));
   NOR2_X1 i_1236 (.A1(n_3300), .A2(n_3258), .ZN(n_2166));
   NOR2_X1 i_1237 (.A1(n_3300), .A2(n_3257), .ZN(n_2167));
   NOR2_X1 i_1238 (.A1(n_3300), .A2(n_3256), .ZN(n_2168));
   NOR2_X1 i_1239 (.A1(n_3300), .A2(n_3255), .ZN(n_2169));
   NOR2_X1 i_1240 (.A1(n_3300), .A2(n_3254), .ZN(n_2170));
   NOR2_X1 i_1241 (.A1(n_3300), .A2(n_3253), .ZN(n_2171));
   NOR2_X1 i_1242 (.A1(n_3300), .A2(n_3252), .ZN(n_2172));
   NOR2_X1 i_1243 (.A1(n_3300), .A2(n_3251), .ZN(n_2173));
   NOR2_X1 i_1244 (.A1(n_3300), .A2(n_3250), .ZN(n_2174));
   NOR2_X1 i_1245 (.A1(n_3300), .A2(n_3249), .ZN(n_2175));
   NOR2_X1 i_1246 (.A1(n_3300), .A2(n_3248), .ZN(n_2176));
   NOR2_X1 i_1247 (.A1(n_3300), .A2(n_3247), .ZN(n_2177));
   NOR2_X1 i_1248 (.A1(n_3300), .A2(n_3246), .ZN(n_2178));
   NOR2_X1 i_1249 (.A1(n_3299), .A2(n_3277), .ZN(n_2179));
   NOR2_X1 i_1250 (.A1(n_3299), .A2(n_3276), .ZN(n_2180));
   NOR2_X1 i_1251 (.A1(n_3299), .A2(n_3275), .ZN(n_2181));
   NOR2_X1 i_1252 (.A1(n_3299), .A2(n_3274), .ZN(n_2182));
   NOR2_X1 i_1253 (.A1(n_3299), .A2(n_3273), .ZN(n_2183));
   NOR2_X1 i_1254 (.A1(n_3299), .A2(n_3272), .ZN(n_2184));
   NOR2_X1 i_1255 (.A1(n_3299), .A2(n_3271), .ZN(n_2185));
   NOR2_X1 i_1256 (.A1(n_3299), .A2(n_3270), .ZN(n_2186));
   NOR2_X1 i_1257 (.A1(n_3299), .A2(n_3269), .ZN(n_2187));
   NOR2_X1 i_1258 (.A1(n_3299), .A2(n_3268), .ZN(n_2188));
   NOR2_X1 i_1259 (.A1(n_3299), .A2(n_3267), .ZN(n_2189));
   NOR2_X1 i_1260 (.A1(n_3299), .A2(n_3266), .ZN(n_2190));
   NOR2_X1 i_1261 (.A1(n_3299), .A2(n_3265), .ZN(n_2191));
   NOR2_X1 i_1262 (.A1(n_3299), .A2(n_3264), .ZN(n_2192));
   NOR2_X1 i_1263 (.A1(n_3299), .A2(n_3263), .ZN(n_2193));
   NOR2_X1 i_1264 (.A1(n_3299), .A2(n_3262), .ZN(n_2194));
   NOR2_X1 i_1265 (.A1(n_3299), .A2(n_3261), .ZN(n_2195));
   NOR2_X1 i_1266 (.A1(n_3299), .A2(n_3260), .ZN(n_2196));
   NOR2_X1 i_1267 (.A1(n_3299), .A2(n_3259), .ZN(n_2197));
   NOR2_X1 i_1268 (.A1(n_3299), .A2(n_3258), .ZN(n_2198));
   NOR2_X1 i_1269 (.A1(n_3299), .A2(n_3257), .ZN(n_2199));
   NOR2_X1 i_1270 (.A1(n_3299), .A2(n_3256), .ZN(n_2200));
   NOR2_X1 i_1271 (.A1(n_3299), .A2(n_3255), .ZN(n_2201));
   NOR2_X1 i_1272 (.A1(n_3299), .A2(n_3254), .ZN(n_2202));
   NOR2_X1 i_1273 (.A1(n_3299), .A2(n_3253), .ZN(n_2203));
   NOR2_X1 i_1274 (.A1(n_3299), .A2(n_3252), .ZN(n_2204));
   NOR2_X1 i_1275 (.A1(n_3299), .A2(n_3251), .ZN(n_2205));
   NOR2_X1 i_1276 (.A1(n_3299), .A2(n_3250), .ZN(n_2206));
   NOR2_X1 i_1277 (.A1(n_3299), .A2(n_3249), .ZN(n_2207));
   NOR2_X1 i_1278 (.A1(n_3299), .A2(n_3248), .ZN(n_2208));
   NOR2_X1 i_1279 (.A1(n_3299), .A2(n_3247), .ZN(n_2209));
   NOR2_X1 i_1280 (.A1(n_3299), .A2(n_3246), .ZN(n_2210));
   NOR2_X1 i_1281 (.A1(n_3298), .A2(n_3277), .ZN(n_2211));
   NOR2_X1 i_1282 (.A1(n_3298), .A2(n_3276), .ZN(n_2212));
   NOR2_X1 i_1283 (.A1(n_3298), .A2(n_3275), .ZN(n_2213));
   NOR2_X1 i_1284 (.A1(n_3298), .A2(n_3274), .ZN(n_2214));
   NOR2_X1 i_1285 (.A1(n_3298), .A2(n_3273), .ZN(n_2215));
   NOR2_X1 i_1286 (.A1(n_3298), .A2(n_3272), .ZN(n_2216));
   NOR2_X1 i_1287 (.A1(n_3298), .A2(n_3271), .ZN(n_2217));
   NOR2_X1 i_1288 (.A1(n_3298), .A2(n_3270), .ZN(n_2218));
   NOR2_X1 i_1289 (.A1(n_3298), .A2(n_3269), .ZN(n_2219));
   NOR2_X1 i_1290 (.A1(n_3298), .A2(n_3268), .ZN(n_2220));
   NOR2_X1 i_1291 (.A1(n_3298), .A2(n_3267), .ZN(n_2221));
   NOR2_X1 i_1292 (.A1(n_3298), .A2(n_3266), .ZN(n_2222));
   NOR2_X1 i_1293 (.A1(n_3298), .A2(n_3265), .ZN(n_2223));
   NOR2_X1 i_1294 (.A1(n_3298), .A2(n_3264), .ZN(n_2224));
   NOR2_X1 i_1295 (.A1(n_3298), .A2(n_3263), .ZN(n_2225));
   NOR2_X1 i_1296 (.A1(n_3298), .A2(n_3262), .ZN(n_2226));
   NOR2_X1 i_1297 (.A1(n_3298), .A2(n_3261), .ZN(n_2227));
   NOR2_X1 i_1298 (.A1(n_3298), .A2(n_3260), .ZN(n_2228));
   NOR2_X1 i_1299 (.A1(n_3298), .A2(n_3259), .ZN(n_2229));
   NOR2_X1 i_1300 (.A1(n_3298), .A2(n_3258), .ZN(n_2230));
   NOR2_X1 i_1301 (.A1(n_3298), .A2(n_3257), .ZN(n_2231));
   NOR2_X1 i_1302 (.A1(n_3298), .A2(n_3256), .ZN(n_2232));
   NOR2_X1 i_1303 (.A1(n_3298), .A2(n_3255), .ZN(n_2233));
   NOR2_X1 i_1304 (.A1(n_3298), .A2(n_3254), .ZN(n_2234));
   NOR2_X1 i_1305 (.A1(n_3298), .A2(n_3253), .ZN(n_2235));
   NOR2_X1 i_1306 (.A1(n_3298), .A2(n_3252), .ZN(n_2236));
   NOR2_X1 i_1307 (.A1(n_3298), .A2(n_3251), .ZN(n_2237));
   NOR2_X1 i_1308 (.A1(n_3298), .A2(n_3250), .ZN(n_2238));
   NOR2_X1 i_1309 (.A1(n_3298), .A2(n_3249), .ZN(n_2239));
   NOR2_X1 i_1310 (.A1(n_3298), .A2(n_3248), .ZN(n_2240));
   NOR2_X1 i_1311 (.A1(n_3298), .A2(n_3247), .ZN(n_2241));
   NOR2_X1 i_1312 (.A1(n_3298), .A2(n_3246), .ZN(n_2242));
   NOR2_X1 i_1313 (.A1(n_3297), .A2(n_3277), .ZN(n_2243));
   NOR2_X1 i_1314 (.A1(n_3297), .A2(n_3276), .ZN(n_2244));
   NOR2_X1 i_1315 (.A1(n_3297), .A2(n_3275), .ZN(n_2245));
   NOR2_X1 i_1316 (.A1(n_3297), .A2(n_3274), .ZN(n_2246));
   NOR2_X1 i_1317 (.A1(n_3297), .A2(n_3273), .ZN(n_2247));
   NOR2_X1 i_1318 (.A1(n_3297), .A2(n_3272), .ZN(n_2248));
   NOR2_X1 i_1319 (.A1(n_3297), .A2(n_3271), .ZN(n_2249));
   NOR2_X1 i_1320 (.A1(n_3297), .A2(n_3270), .ZN(n_2250));
   NOR2_X1 i_1321 (.A1(n_3297), .A2(n_3269), .ZN(n_2251));
   NOR2_X1 i_1322 (.A1(n_3297), .A2(n_3268), .ZN(n_2252));
   NOR2_X1 i_1323 (.A1(n_3297), .A2(n_3267), .ZN(n_2253));
   NOR2_X1 i_1324 (.A1(n_3297), .A2(n_3266), .ZN(n_2254));
   NOR2_X1 i_1325 (.A1(n_3297), .A2(n_3265), .ZN(n_2255));
   NOR2_X1 i_1326 (.A1(n_3297), .A2(n_3264), .ZN(n_2256));
   NOR2_X1 i_1327 (.A1(n_3297), .A2(n_3263), .ZN(n_2257));
   NOR2_X1 i_1328 (.A1(n_3297), .A2(n_3262), .ZN(n_2258));
   NOR2_X1 i_1329 (.A1(n_3297), .A2(n_3261), .ZN(n_2259));
   NOR2_X1 i_1330 (.A1(n_3297), .A2(n_3260), .ZN(n_2260));
   NOR2_X1 i_1331 (.A1(n_3297), .A2(n_3259), .ZN(n_2261));
   NOR2_X1 i_1332 (.A1(n_3297), .A2(n_3258), .ZN(n_2262));
   NOR2_X1 i_1333 (.A1(n_3297), .A2(n_3257), .ZN(n_2263));
   NOR2_X1 i_1334 (.A1(n_3297), .A2(n_3256), .ZN(n_2264));
   NOR2_X1 i_1335 (.A1(n_3297), .A2(n_3255), .ZN(n_2265));
   NOR2_X1 i_1336 (.A1(n_3297), .A2(n_3254), .ZN(n_2266));
   NOR2_X1 i_1337 (.A1(n_3297), .A2(n_3253), .ZN(n_2267));
   NOR2_X1 i_1338 (.A1(n_3297), .A2(n_3252), .ZN(n_2268));
   NOR2_X1 i_1339 (.A1(n_3297), .A2(n_3251), .ZN(n_2269));
   NOR2_X1 i_1340 (.A1(n_3297), .A2(n_3250), .ZN(n_2270));
   NOR2_X1 i_1341 (.A1(n_3297), .A2(n_3249), .ZN(n_2271));
   NOR2_X1 i_1342 (.A1(n_3297), .A2(n_3248), .ZN(n_2272));
   NOR2_X1 i_1343 (.A1(n_3297), .A2(n_3247), .ZN(n_2273));
   NOR2_X1 i_1344 (.A1(n_3297), .A2(n_3246), .ZN(n_2274));
   NOR2_X1 i_1345 (.A1(n_3296), .A2(n_3277), .ZN(n_2275));
   NOR2_X1 i_1346 (.A1(n_3296), .A2(n_3276), .ZN(n_2276));
   NOR2_X1 i_1347 (.A1(n_3296), .A2(n_3275), .ZN(n_2277));
   NOR2_X1 i_1348 (.A1(n_3296), .A2(n_3274), .ZN(n_2278));
   NOR2_X1 i_1349 (.A1(n_3296), .A2(n_3273), .ZN(n_2279));
   NOR2_X1 i_1350 (.A1(n_3296), .A2(n_3272), .ZN(n_2280));
   NOR2_X1 i_1351 (.A1(n_3296), .A2(n_3271), .ZN(n_2281));
   NOR2_X1 i_1352 (.A1(n_3296), .A2(n_3270), .ZN(n_2282));
   NOR2_X1 i_1353 (.A1(n_3296), .A2(n_3269), .ZN(n_2283));
   NOR2_X1 i_1354 (.A1(n_3296), .A2(n_3268), .ZN(n_2284));
   NOR2_X1 i_1355 (.A1(n_3296), .A2(n_3267), .ZN(n_2285));
   NOR2_X1 i_1356 (.A1(n_3296), .A2(n_3266), .ZN(n_2286));
   NOR2_X1 i_1357 (.A1(n_3296), .A2(n_3265), .ZN(n_2287));
   NOR2_X1 i_1358 (.A1(n_3296), .A2(n_3264), .ZN(n_2288));
   NOR2_X1 i_1359 (.A1(n_3296), .A2(n_3263), .ZN(n_2289));
   NOR2_X1 i_1360 (.A1(n_3296), .A2(n_3262), .ZN(n_2290));
   NOR2_X1 i_1361 (.A1(n_3296), .A2(n_3261), .ZN(n_2291));
   NOR2_X1 i_1362 (.A1(n_3296), .A2(n_3260), .ZN(n_2292));
   NOR2_X1 i_1363 (.A1(n_3296), .A2(n_3259), .ZN(n_2293));
   NOR2_X1 i_1364 (.A1(n_3296), .A2(n_3258), .ZN(n_2294));
   NOR2_X1 i_1365 (.A1(n_3296), .A2(n_3257), .ZN(n_2295));
   NOR2_X1 i_1366 (.A1(n_3296), .A2(n_3256), .ZN(n_2296));
   NOR2_X1 i_1367 (.A1(n_3296), .A2(n_3255), .ZN(n_2297));
   NOR2_X1 i_1368 (.A1(n_3296), .A2(n_3254), .ZN(n_2298));
   NOR2_X1 i_1369 (.A1(n_3296), .A2(n_3253), .ZN(n_2299));
   NOR2_X1 i_1370 (.A1(n_3296), .A2(n_3252), .ZN(n_2300));
   NOR2_X1 i_1371 (.A1(n_3296), .A2(n_3251), .ZN(n_2301));
   NOR2_X1 i_1372 (.A1(n_3296), .A2(n_3250), .ZN(n_2302));
   NOR2_X1 i_1373 (.A1(n_3296), .A2(n_3249), .ZN(n_2303));
   NOR2_X1 i_1374 (.A1(n_3296), .A2(n_3248), .ZN(n_2304));
   NOR2_X1 i_1375 (.A1(n_3296), .A2(n_3247), .ZN(n_2305));
   NOR2_X1 i_1376 (.A1(n_3296), .A2(n_3246), .ZN(n_2306));
   NOR2_X1 i_1377 (.A1(n_3295), .A2(n_3277), .ZN(n_2307));
   NOR2_X1 i_1378 (.A1(n_3295), .A2(n_3276), .ZN(n_2308));
   NOR2_X1 i_1379 (.A1(n_3295), .A2(n_3275), .ZN(n_2309));
   NOR2_X1 i_1380 (.A1(n_3295), .A2(n_3274), .ZN(n_2310));
   NOR2_X1 i_1381 (.A1(n_3295), .A2(n_3273), .ZN(n_2311));
   NOR2_X1 i_1382 (.A1(n_3295), .A2(n_3272), .ZN(n_2312));
   NOR2_X1 i_1383 (.A1(n_3295), .A2(n_3271), .ZN(n_2313));
   NOR2_X1 i_1384 (.A1(n_3295), .A2(n_3270), .ZN(n_2314));
   NOR2_X1 i_1385 (.A1(n_3295), .A2(n_3269), .ZN(n_2315));
   NOR2_X1 i_1386 (.A1(n_3295), .A2(n_3268), .ZN(n_2316));
   NOR2_X1 i_1387 (.A1(n_3295), .A2(n_3267), .ZN(n_2317));
   NOR2_X1 i_1388 (.A1(n_3295), .A2(n_3266), .ZN(n_2318));
   NOR2_X1 i_1389 (.A1(n_3295), .A2(n_3265), .ZN(n_2319));
   NOR2_X1 i_1390 (.A1(n_3295), .A2(n_3264), .ZN(n_2320));
   NOR2_X1 i_1391 (.A1(n_3295), .A2(n_3263), .ZN(n_2321));
   NOR2_X1 i_1392 (.A1(n_3295), .A2(n_3262), .ZN(n_2322));
   NOR2_X1 i_1393 (.A1(n_3295), .A2(n_3261), .ZN(n_2323));
   NOR2_X1 i_1394 (.A1(n_3295), .A2(n_3260), .ZN(n_2324));
   NOR2_X1 i_1395 (.A1(n_3295), .A2(n_3259), .ZN(n_2325));
   NOR2_X1 i_1396 (.A1(n_3295), .A2(n_3258), .ZN(n_2326));
   NOR2_X1 i_1397 (.A1(n_3295), .A2(n_3257), .ZN(n_2327));
   NOR2_X1 i_1398 (.A1(n_3295), .A2(n_3256), .ZN(n_2328));
   NOR2_X1 i_1399 (.A1(n_3295), .A2(n_3255), .ZN(n_2329));
   NOR2_X1 i_1400 (.A1(n_3295), .A2(n_3254), .ZN(n_2330));
   NOR2_X1 i_1401 (.A1(n_3295), .A2(n_3253), .ZN(n_2331));
   NOR2_X1 i_1402 (.A1(n_3295), .A2(n_3252), .ZN(n_2332));
   NOR2_X1 i_1403 (.A1(n_3295), .A2(n_3251), .ZN(n_2333));
   NOR2_X1 i_1404 (.A1(n_3295), .A2(n_3250), .ZN(n_2334));
   NOR2_X1 i_1405 (.A1(n_3295), .A2(n_3249), .ZN(n_2335));
   NOR2_X1 i_1406 (.A1(n_3295), .A2(n_3248), .ZN(n_2336));
   NOR2_X1 i_1407 (.A1(n_3295), .A2(n_3247), .ZN(n_2337));
   NOR2_X1 i_1408 (.A1(n_3295), .A2(n_3246), .ZN(n_2338));
   NOR2_X1 i_1409 (.A1(n_3294), .A2(n_3277), .ZN(n_2339));
   NOR2_X1 i_1410 (.A1(n_3294), .A2(n_3276), .ZN(n_2340));
   NOR2_X1 i_1411 (.A1(n_3294), .A2(n_3275), .ZN(n_2341));
   NOR2_X1 i_1412 (.A1(n_3294), .A2(n_3274), .ZN(n_2342));
   NOR2_X1 i_1413 (.A1(n_3294), .A2(n_3273), .ZN(n_2343));
   NOR2_X1 i_1414 (.A1(n_3294), .A2(n_3272), .ZN(n_2344));
   NOR2_X1 i_1415 (.A1(n_3294), .A2(n_3271), .ZN(n_2345));
   NOR2_X1 i_1416 (.A1(n_3294), .A2(n_3270), .ZN(n_2346));
   NOR2_X1 i_1417 (.A1(n_3294), .A2(n_3269), .ZN(n_2347));
   NOR2_X1 i_1418 (.A1(n_3294), .A2(n_3268), .ZN(n_2348));
   NOR2_X1 i_1419 (.A1(n_3294), .A2(n_3267), .ZN(n_2349));
   NOR2_X1 i_1420 (.A1(n_3294), .A2(n_3266), .ZN(n_2350));
   NOR2_X1 i_1421 (.A1(n_3294), .A2(n_3265), .ZN(n_2351));
   NOR2_X1 i_1422 (.A1(n_3294), .A2(n_3264), .ZN(n_2352));
   NOR2_X1 i_1423 (.A1(n_3294), .A2(n_3263), .ZN(n_2353));
   NOR2_X1 i_1424 (.A1(n_3294), .A2(n_3262), .ZN(n_2354));
   NOR2_X1 i_1425 (.A1(n_3294), .A2(n_3261), .ZN(n_2355));
   NOR2_X1 i_1426 (.A1(n_3294), .A2(n_3260), .ZN(n_2356));
   NOR2_X1 i_1427 (.A1(n_3294), .A2(n_3259), .ZN(n_2357));
   NOR2_X1 i_1428 (.A1(n_3294), .A2(n_3258), .ZN(n_2358));
   NOR2_X1 i_1429 (.A1(n_3294), .A2(n_3257), .ZN(n_2359));
   NOR2_X1 i_1430 (.A1(n_3294), .A2(n_3256), .ZN(n_2360));
   NOR2_X1 i_1431 (.A1(n_3294), .A2(n_3255), .ZN(n_2361));
   NOR2_X1 i_1432 (.A1(n_3294), .A2(n_3254), .ZN(n_2362));
   NOR2_X1 i_1433 (.A1(n_3294), .A2(n_3253), .ZN(n_2363));
   NOR2_X1 i_1434 (.A1(n_3294), .A2(n_3252), .ZN(n_2364));
   NOR2_X1 i_1435 (.A1(n_3294), .A2(n_3251), .ZN(n_2365));
   NOR2_X1 i_1436 (.A1(n_3294), .A2(n_3250), .ZN(n_2366));
   NOR2_X1 i_1437 (.A1(n_3294), .A2(n_3249), .ZN(n_2367));
   NOR2_X1 i_1438 (.A1(n_3294), .A2(n_3248), .ZN(n_2368));
   NOR2_X1 i_1439 (.A1(n_3294), .A2(n_3247), .ZN(n_2369));
   NOR2_X1 i_1440 (.A1(n_3294), .A2(n_3246), .ZN(n_2370));
   NOR2_X1 i_1441 (.A1(n_3293), .A2(n_3277), .ZN(n_2371));
   NOR2_X1 i_1442 (.A1(n_3293), .A2(n_3276), .ZN(n_2372));
   NOR2_X1 i_1443 (.A1(n_3293), .A2(n_3275), .ZN(n_2373));
   NOR2_X1 i_1444 (.A1(n_3293), .A2(n_3274), .ZN(n_2374));
   NOR2_X1 i_1445 (.A1(n_3293), .A2(n_3273), .ZN(n_2375));
   NOR2_X1 i_1446 (.A1(n_3293), .A2(n_3272), .ZN(n_2376));
   NOR2_X1 i_1447 (.A1(n_3293), .A2(n_3271), .ZN(n_2377));
   NOR2_X1 i_1448 (.A1(n_3293), .A2(n_3270), .ZN(n_2378));
   NOR2_X1 i_1449 (.A1(n_3293), .A2(n_3269), .ZN(n_2379));
   NOR2_X1 i_1450 (.A1(n_3293), .A2(n_3268), .ZN(n_2380));
   NOR2_X1 i_1451 (.A1(n_3293), .A2(n_3267), .ZN(n_2381));
   NOR2_X1 i_1452 (.A1(n_3293), .A2(n_3266), .ZN(n_2382));
   NOR2_X1 i_1453 (.A1(n_3293), .A2(n_3265), .ZN(n_2383));
   NOR2_X1 i_1454 (.A1(n_3293), .A2(n_3264), .ZN(n_2384));
   NOR2_X1 i_1455 (.A1(n_3293), .A2(n_3263), .ZN(n_2385));
   NOR2_X1 i_1456 (.A1(n_3293), .A2(n_3262), .ZN(n_2386));
   NOR2_X1 i_1457 (.A1(n_3293), .A2(n_3261), .ZN(n_2387));
   NOR2_X1 i_1458 (.A1(n_3293), .A2(n_3260), .ZN(n_2388));
   NOR2_X1 i_1459 (.A1(n_3293), .A2(n_3259), .ZN(n_2389));
   NOR2_X1 i_1460 (.A1(n_3293), .A2(n_3258), .ZN(n_2390));
   NOR2_X1 i_1461 (.A1(n_3293), .A2(n_3257), .ZN(n_2391));
   NOR2_X1 i_1462 (.A1(n_3293), .A2(n_3256), .ZN(n_2392));
   NOR2_X1 i_1463 (.A1(n_3293), .A2(n_3255), .ZN(n_2393));
   NOR2_X1 i_1464 (.A1(n_3293), .A2(n_3254), .ZN(n_2394));
   NOR2_X1 i_1465 (.A1(n_3293), .A2(n_3253), .ZN(n_2395));
   NOR2_X1 i_1466 (.A1(n_3293), .A2(n_3252), .ZN(n_2396));
   NOR2_X1 i_1467 (.A1(n_3293), .A2(n_3251), .ZN(n_2397));
   NOR2_X1 i_1468 (.A1(n_3293), .A2(n_3250), .ZN(n_2398));
   NOR2_X1 i_1469 (.A1(n_3293), .A2(n_3249), .ZN(n_2399));
   NOR2_X1 i_1470 (.A1(n_3293), .A2(n_3248), .ZN(n_2400));
   NOR2_X1 i_1471 (.A1(n_3293), .A2(n_3247), .ZN(n_2401));
   NOR2_X1 i_1472 (.A1(n_3293), .A2(n_3246), .ZN(n_2402));
   NOR2_X1 i_1473 (.A1(n_3292), .A2(n_3277), .ZN(n_2403));
   NOR2_X1 i_1474 (.A1(n_3292), .A2(n_3276), .ZN(n_2404));
   NOR2_X1 i_1475 (.A1(n_3292), .A2(n_3275), .ZN(n_2405));
   NOR2_X1 i_1476 (.A1(n_3292), .A2(n_3274), .ZN(n_2406));
   NOR2_X1 i_1477 (.A1(n_3292), .A2(n_3273), .ZN(n_2407));
   NOR2_X1 i_1478 (.A1(n_3292), .A2(n_3272), .ZN(n_2408));
   NOR2_X1 i_1479 (.A1(n_3292), .A2(n_3271), .ZN(n_2409));
   NOR2_X1 i_1480 (.A1(n_3292), .A2(n_3270), .ZN(n_2410));
   NOR2_X1 i_1481 (.A1(n_3292), .A2(n_3269), .ZN(n_2411));
   NOR2_X1 i_1482 (.A1(n_3292), .A2(n_3268), .ZN(n_2412));
   NOR2_X1 i_1483 (.A1(n_3292), .A2(n_3267), .ZN(n_2413));
   NOR2_X1 i_1484 (.A1(n_3292), .A2(n_3266), .ZN(n_2414));
   NOR2_X1 i_1485 (.A1(n_3292), .A2(n_3265), .ZN(n_2415));
   NOR2_X1 i_1486 (.A1(n_3292), .A2(n_3264), .ZN(n_2416));
   NOR2_X1 i_1487 (.A1(n_3292), .A2(n_3263), .ZN(n_2417));
   NOR2_X1 i_1488 (.A1(n_3292), .A2(n_3262), .ZN(n_2418));
   NOR2_X1 i_1489 (.A1(n_3292), .A2(n_3261), .ZN(n_2419));
   NOR2_X1 i_1490 (.A1(n_3292), .A2(n_3260), .ZN(n_2420));
   NOR2_X1 i_1491 (.A1(n_3292), .A2(n_3259), .ZN(n_2421));
   NOR2_X1 i_1492 (.A1(n_3292), .A2(n_3258), .ZN(n_2422));
   NOR2_X1 i_1493 (.A1(n_3292), .A2(n_3257), .ZN(n_2423));
   NOR2_X1 i_1494 (.A1(n_3292), .A2(n_3256), .ZN(n_2424));
   NOR2_X1 i_1495 (.A1(n_3292), .A2(n_3255), .ZN(n_2425));
   NOR2_X1 i_1496 (.A1(n_3292), .A2(n_3254), .ZN(n_2426));
   NOR2_X1 i_1497 (.A1(n_3292), .A2(n_3253), .ZN(n_2427));
   NOR2_X1 i_1498 (.A1(n_3292), .A2(n_3252), .ZN(n_2428));
   NOR2_X1 i_1499 (.A1(n_3292), .A2(n_3251), .ZN(n_2429));
   NOR2_X1 i_1500 (.A1(n_3292), .A2(n_3250), .ZN(n_2430));
   NOR2_X1 i_1501 (.A1(n_3292), .A2(n_3249), .ZN(n_2431));
   NOR2_X1 i_1502 (.A1(n_3292), .A2(n_3248), .ZN(n_2432));
   NOR2_X1 i_1503 (.A1(n_3292), .A2(n_3247), .ZN(n_2433));
   NOR2_X1 i_1504 (.A1(n_3292), .A2(n_3246), .ZN(n_2434));
   NOR2_X1 i_1505 (.A1(n_3291), .A2(n_3277), .ZN(n_2435));
   NOR2_X1 i_1506 (.A1(n_3291), .A2(n_3276), .ZN(n_2436));
   NOR2_X1 i_1507 (.A1(n_3291), .A2(n_3275), .ZN(n_2437));
   NOR2_X1 i_1508 (.A1(n_3291), .A2(n_3274), .ZN(n_2438));
   NOR2_X1 i_1509 (.A1(n_3291), .A2(n_3273), .ZN(n_2439));
   NOR2_X1 i_1510 (.A1(n_3291), .A2(n_3272), .ZN(n_2440));
   NOR2_X1 i_1511 (.A1(n_3291), .A2(n_3271), .ZN(n_2441));
   NOR2_X1 i_1512 (.A1(n_3291), .A2(n_3270), .ZN(n_2442));
   NOR2_X1 i_1513 (.A1(n_3291), .A2(n_3269), .ZN(n_2443));
   NOR2_X1 i_1514 (.A1(n_3291), .A2(n_3268), .ZN(n_2444));
   NOR2_X1 i_1515 (.A1(n_3291), .A2(n_3267), .ZN(n_2445));
   NOR2_X1 i_1516 (.A1(n_3291), .A2(n_3266), .ZN(n_2446));
   NOR2_X1 i_1517 (.A1(n_3291), .A2(n_3265), .ZN(n_2447));
   NOR2_X1 i_1518 (.A1(n_3291), .A2(n_3264), .ZN(n_2448));
   NOR2_X1 i_1519 (.A1(n_3291), .A2(n_3263), .ZN(n_2449));
   NOR2_X1 i_1520 (.A1(n_3291), .A2(n_3262), .ZN(n_2450));
   NOR2_X1 i_1521 (.A1(n_3291), .A2(n_3261), .ZN(n_2451));
   NOR2_X1 i_1522 (.A1(n_3291), .A2(n_3260), .ZN(n_2452));
   NOR2_X1 i_1523 (.A1(n_3291), .A2(n_3259), .ZN(n_2453));
   NOR2_X1 i_1524 (.A1(n_3291), .A2(n_3258), .ZN(n_2454));
   NOR2_X1 i_1525 (.A1(n_3291), .A2(n_3257), .ZN(n_2455));
   NOR2_X1 i_1526 (.A1(n_3291), .A2(n_3256), .ZN(n_2456));
   NOR2_X1 i_1527 (.A1(n_3291), .A2(n_3255), .ZN(n_2457));
   NOR2_X1 i_1528 (.A1(n_3291), .A2(n_3254), .ZN(n_2458));
   NOR2_X1 i_1529 (.A1(n_3291), .A2(n_3253), .ZN(n_2459));
   NOR2_X1 i_1530 (.A1(n_3291), .A2(n_3252), .ZN(n_2460));
   NOR2_X1 i_1531 (.A1(n_3291), .A2(n_3251), .ZN(n_2461));
   NOR2_X1 i_1532 (.A1(n_3291), .A2(n_3250), .ZN(n_2462));
   NOR2_X1 i_1533 (.A1(n_3291), .A2(n_3249), .ZN(n_2463));
   NOR2_X1 i_1534 (.A1(n_3291), .A2(n_3248), .ZN(n_2464));
   NOR2_X1 i_1535 (.A1(n_3291), .A2(n_3247), .ZN(n_2465));
   NOR2_X1 i_1536 (.A1(n_3291), .A2(n_3246), .ZN(n_2466));
   NOR2_X1 i_1537 (.A1(n_3290), .A2(n_3277), .ZN(n_2467));
   NOR2_X1 i_1538 (.A1(n_3290), .A2(n_3276), .ZN(n_2468));
   NOR2_X1 i_1539 (.A1(n_3290), .A2(n_3275), .ZN(n_2469));
   NOR2_X1 i_1540 (.A1(n_3290), .A2(n_3274), .ZN(n_2470));
   NOR2_X1 i_1541 (.A1(n_3290), .A2(n_3273), .ZN(n_2471));
   NOR2_X1 i_1542 (.A1(n_3290), .A2(n_3272), .ZN(n_2472));
   NOR2_X1 i_1543 (.A1(n_3290), .A2(n_3271), .ZN(n_2473));
   NOR2_X1 i_1544 (.A1(n_3290), .A2(n_3270), .ZN(n_2474));
   NOR2_X1 i_1545 (.A1(n_3290), .A2(n_3269), .ZN(n_2475));
   NOR2_X1 i_1546 (.A1(n_3290), .A2(n_3268), .ZN(n_2476));
   NOR2_X1 i_1547 (.A1(n_3290), .A2(n_3267), .ZN(n_2477));
   NOR2_X1 i_1548 (.A1(n_3290), .A2(n_3266), .ZN(n_2478));
   NOR2_X1 i_1549 (.A1(n_3290), .A2(n_3265), .ZN(n_2479));
   NOR2_X1 i_1550 (.A1(n_3290), .A2(n_3264), .ZN(n_2480));
   NOR2_X1 i_1551 (.A1(n_3290), .A2(n_3263), .ZN(n_2481));
   NOR2_X1 i_1552 (.A1(n_3290), .A2(n_3262), .ZN(n_2482));
   NOR2_X1 i_1553 (.A1(n_3290), .A2(n_3261), .ZN(n_2483));
   NOR2_X1 i_1554 (.A1(n_3290), .A2(n_3260), .ZN(n_2484));
   NOR2_X1 i_1555 (.A1(n_3290), .A2(n_3259), .ZN(n_2485));
   NOR2_X1 i_1556 (.A1(n_3290), .A2(n_3258), .ZN(n_2486));
   NOR2_X1 i_1557 (.A1(n_3290), .A2(n_3257), .ZN(n_2487));
   NOR2_X1 i_1558 (.A1(n_3290), .A2(n_3256), .ZN(n_2488));
   NOR2_X1 i_1559 (.A1(n_3290), .A2(n_3255), .ZN(n_2489));
   NOR2_X1 i_1560 (.A1(n_3290), .A2(n_3254), .ZN(n_2490));
   NOR2_X1 i_1561 (.A1(n_3290), .A2(n_3253), .ZN(n_2491));
   NOR2_X1 i_1562 (.A1(n_3290), .A2(n_3252), .ZN(n_2492));
   NOR2_X1 i_1563 (.A1(n_3290), .A2(n_3251), .ZN(n_2493));
   NOR2_X1 i_1564 (.A1(n_3290), .A2(n_3250), .ZN(n_2494));
   NOR2_X1 i_1565 (.A1(n_3290), .A2(n_3249), .ZN(n_2495));
   NOR2_X1 i_1566 (.A1(n_3290), .A2(n_3248), .ZN(n_2496));
   NOR2_X1 i_1567 (.A1(n_3290), .A2(n_3247), .ZN(n_2497));
   NOR2_X1 i_1568 (.A1(n_3290), .A2(n_3246), .ZN(n_2498));
   NOR2_X1 i_1569 (.A1(n_3289), .A2(n_3277), .ZN(n_2499));
   NOR2_X1 i_1570 (.A1(n_3289), .A2(n_3276), .ZN(n_2500));
   NOR2_X1 i_1571 (.A1(n_3289), .A2(n_3275), .ZN(n_2501));
   NOR2_X1 i_1572 (.A1(n_3289), .A2(n_3274), .ZN(n_2502));
   NOR2_X1 i_1573 (.A1(n_3289), .A2(n_3273), .ZN(n_2503));
   NOR2_X1 i_1574 (.A1(n_3289), .A2(n_3272), .ZN(n_2504));
   NOR2_X1 i_1575 (.A1(n_3289), .A2(n_3271), .ZN(n_2505));
   NOR2_X1 i_1576 (.A1(n_3289), .A2(n_3270), .ZN(n_2506));
   NOR2_X1 i_1577 (.A1(n_3289), .A2(n_3269), .ZN(n_2507));
   NOR2_X1 i_1578 (.A1(n_3289), .A2(n_3268), .ZN(n_2508));
   NOR2_X1 i_1579 (.A1(n_3289), .A2(n_3267), .ZN(n_2509));
   NOR2_X1 i_1580 (.A1(n_3289), .A2(n_3266), .ZN(n_2510));
   NOR2_X1 i_1581 (.A1(n_3289), .A2(n_3265), .ZN(n_2511));
   NOR2_X1 i_1582 (.A1(n_3289), .A2(n_3264), .ZN(n_2512));
   NOR2_X1 i_1583 (.A1(n_3289), .A2(n_3263), .ZN(n_2513));
   NOR2_X1 i_1584 (.A1(n_3289), .A2(n_3262), .ZN(n_2514));
   NOR2_X1 i_1585 (.A1(n_3289), .A2(n_3261), .ZN(n_2515));
   NOR2_X1 i_1586 (.A1(n_3289), .A2(n_3260), .ZN(n_2516));
   NOR2_X1 i_1587 (.A1(n_3289), .A2(n_3259), .ZN(n_2517));
   NOR2_X1 i_1588 (.A1(n_3289), .A2(n_3258), .ZN(n_2518));
   NOR2_X1 i_1589 (.A1(n_3289), .A2(n_3257), .ZN(n_2519));
   NOR2_X1 i_1590 (.A1(n_3289), .A2(n_3256), .ZN(n_2520));
   NOR2_X1 i_1591 (.A1(n_3289), .A2(n_3255), .ZN(n_2521));
   NOR2_X1 i_1592 (.A1(n_3289), .A2(n_3254), .ZN(n_2522));
   NOR2_X1 i_1593 (.A1(n_3289), .A2(n_3253), .ZN(n_2523));
   NOR2_X1 i_1594 (.A1(n_3289), .A2(n_3252), .ZN(n_2524));
   NOR2_X1 i_1595 (.A1(n_3289), .A2(n_3251), .ZN(n_2525));
   NOR2_X1 i_1596 (.A1(n_3289), .A2(n_3250), .ZN(n_2526));
   NOR2_X1 i_1597 (.A1(n_3289), .A2(n_3249), .ZN(n_2527));
   NOR2_X1 i_1598 (.A1(n_3289), .A2(n_3248), .ZN(n_2528));
   NOR2_X1 i_1599 (.A1(n_3289), .A2(n_3247), .ZN(n_2529));
   NOR2_X1 i_1600 (.A1(n_3289), .A2(n_3246), .ZN(n_2530));
   NOR2_X1 i_1601 (.A1(n_3288), .A2(n_3277), .ZN(n_2531));
   NOR2_X1 i_1602 (.A1(n_3288), .A2(n_3276), .ZN(n_2532));
   NOR2_X1 i_1603 (.A1(n_3288), .A2(n_3275), .ZN(n_2533));
   NOR2_X1 i_1604 (.A1(n_3288), .A2(n_3274), .ZN(n_2534));
   NOR2_X1 i_1605 (.A1(n_3288), .A2(n_3273), .ZN(n_2535));
   NOR2_X1 i_1606 (.A1(n_3288), .A2(n_3272), .ZN(n_2536));
   NOR2_X1 i_1607 (.A1(n_3288), .A2(n_3271), .ZN(n_2537));
   NOR2_X1 i_1608 (.A1(n_3288), .A2(n_3270), .ZN(n_2538));
   NOR2_X1 i_1609 (.A1(n_3288), .A2(n_3269), .ZN(n_2539));
   NOR2_X1 i_1610 (.A1(n_3288), .A2(n_3268), .ZN(n_2540));
   NOR2_X1 i_1611 (.A1(n_3288), .A2(n_3267), .ZN(n_2541));
   NOR2_X1 i_1612 (.A1(n_3288), .A2(n_3266), .ZN(n_2542));
   NOR2_X1 i_1613 (.A1(n_3288), .A2(n_3265), .ZN(n_2543));
   NOR2_X1 i_1614 (.A1(n_3288), .A2(n_3264), .ZN(n_2544));
   NOR2_X1 i_1615 (.A1(n_3288), .A2(n_3263), .ZN(n_2545));
   NOR2_X1 i_1616 (.A1(n_3288), .A2(n_3262), .ZN(n_2546));
   NOR2_X1 i_1617 (.A1(n_3288), .A2(n_3261), .ZN(n_2547));
   NOR2_X1 i_1618 (.A1(n_3288), .A2(n_3260), .ZN(n_2548));
   NOR2_X1 i_1619 (.A1(n_3288), .A2(n_3259), .ZN(n_2549));
   NOR2_X1 i_1620 (.A1(n_3288), .A2(n_3258), .ZN(n_2550));
   NOR2_X1 i_1621 (.A1(n_3288), .A2(n_3257), .ZN(n_2551));
   NOR2_X1 i_1622 (.A1(n_3288), .A2(n_3256), .ZN(n_2552));
   NOR2_X1 i_1623 (.A1(n_3288), .A2(n_3255), .ZN(n_2553));
   NOR2_X1 i_1624 (.A1(n_3288), .A2(n_3254), .ZN(n_2554));
   NOR2_X1 i_1625 (.A1(n_3288), .A2(n_3253), .ZN(n_2555));
   NOR2_X1 i_1626 (.A1(n_3288), .A2(n_3252), .ZN(n_2556));
   NOR2_X1 i_1627 (.A1(n_3288), .A2(n_3251), .ZN(n_2557));
   NOR2_X1 i_1628 (.A1(n_3288), .A2(n_3250), .ZN(n_2558));
   NOR2_X1 i_1629 (.A1(n_3288), .A2(n_3249), .ZN(n_2559));
   NOR2_X1 i_1630 (.A1(n_3288), .A2(n_3248), .ZN(n_2560));
   NOR2_X1 i_1631 (.A1(n_3288), .A2(n_3247), .ZN(n_2561));
   NOR2_X1 i_1632 (.A1(n_3288), .A2(n_3246), .ZN(n_2562));
   NOR2_X1 i_1633 (.A1(n_3287), .A2(n_3277), .ZN(n_2563));
   NOR2_X1 i_1634 (.A1(n_3287), .A2(n_3276), .ZN(n_2564));
   NOR2_X1 i_1635 (.A1(n_3287), .A2(n_3275), .ZN(n_2565));
   NOR2_X1 i_1636 (.A1(n_3287), .A2(n_3274), .ZN(n_2566));
   NOR2_X1 i_1637 (.A1(n_3287), .A2(n_3273), .ZN(n_2567));
   NOR2_X1 i_1638 (.A1(n_3287), .A2(n_3272), .ZN(n_2568));
   NOR2_X1 i_1639 (.A1(n_3287), .A2(n_3271), .ZN(n_2569));
   NOR2_X1 i_1640 (.A1(n_3287), .A2(n_3270), .ZN(n_2570));
   NOR2_X1 i_1641 (.A1(n_3287), .A2(n_3269), .ZN(n_2571));
   NOR2_X1 i_1642 (.A1(n_3287), .A2(n_3268), .ZN(n_2572));
   NOR2_X1 i_1643 (.A1(n_3287), .A2(n_3267), .ZN(n_2573));
   NOR2_X1 i_1644 (.A1(n_3287), .A2(n_3266), .ZN(n_2574));
   NOR2_X1 i_1645 (.A1(n_3287), .A2(n_3265), .ZN(n_2575));
   NOR2_X1 i_1646 (.A1(n_3287), .A2(n_3264), .ZN(n_2576));
   NOR2_X1 i_1647 (.A1(n_3287), .A2(n_3263), .ZN(n_2577));
   NOR2_X1 i_1648 (.A1(n_3287), .A2(n_3262), .ZN(n_2578));
   NOR2_X1 i_1649 (.A1(n_3287), .A2(n_3261), .ZN(n_2579));
   NOR2_X1 i_1650 (.A1(n_3287), .A2(n_3260), .ZN(n_2580));
   NOR2_X1 i_1651 (.A1(n_3287), .A2(n_3259), .ZN(n_2581));
   NOR2_X1 i_1652 (.A1(n_3287), .A2(n_3258), .ZN(n_2582));
   NOR2_X1 i_1653 (.A1(n_3287), .A2(n_3257), .ZN(n_2583));
   NOR2_X1 i_1654 (.A1(n_3287), .A2(n_3256), .ZN(n_2584));
   NOR2_X1 i_1655 (.A1(n_3287), .A2(n_3255), .ZN(n_2585));
   NOR2_X1 i_1656 (.A1(n_3287), .A2(n_3254), .ZN(n_2586));
   NOR2_X1 i_1657 (.A1(n_3287), .A2(n_3253), .ZN(n_2587));
   NOR2_X1 i_1658 (.A1(n_3287), .A2(n_3252), .ZN(n_2588));
   NOR2_X1 i_1659 (.A1(n_3287), .A2(n_3251), .ZN(n_2589));
   NOR2_X1 i_1660 (.A1(n_3287), .A2(n_3250), .ZN(n_2590));
   NOR2_X1 i_1661 (.A1(n_3287), .A2(n_3249), .ZN(n_2591));
   NOR2_X1 i_1662 (.A1(n_3287), .A2(n_3248), .ZN(n_2592));
   NOR2_X1 i_1663 (.A1(n_3287), .A2(n_3247), .ZN(n_2593));
   NOR2_X1 i_1664 (.A1(n_3287), .A2(n_3246), .ZN(n_2594));
   NOR2_X1 i_1665 (.A1(n_3286), .A2(n_3277), .ZN(n_2595));
   NOR2_X1 i_1666 (.A1(n_3286), .A2(n_3276), .ZN(n_2596));
   NOR2_X1 i_1667 (.A1(n_3286), .A2(n_3275), .ZN(n_2597));
   NOR2_X1 i_1668 (.A1(n_3286), .A2(n_3274), .ZN(n_2598));
   NOR2_X1 i_1669 (.A1(n_3286), .A2(n_3273), .ZN(n_2599));
   NOR2_X1 i_1670 (.A1(n_3286), .A2(n_3272), .ZN(n_2600));
   NOR2_X1 i_1671 (.A1(n_3286), .A2(n_3271), .ZN(n_2601));
   NOR2_X1 i_1672 (.A1(n_3286), .A2(n_3270), .ZN(n_2602));
   NOR2_X1 i_1673 (.A1(n_3286), .A2(n_3269), .ZN(n_2603));
   NOR2_X1 i_1674 (.A1(n_3286), .A2(n_3268), .ZN(n_2604));
   NOR2_X1 i_1675 (.A1(n_3286), .A2(n_3267), .ZN(n_2605));
   NOR2_X1 i_1676 (.A1(n_3286), .A2(n_3266), .ZN(n_2606));
   NOR2_X1 i_1677 (.A1(n_3286), .A2(n_3265), .ZN(n_2607));
   NOR2_X1 i_1678 (.A1(n_3286), .A2(n_3264), .ZN(n_2608));
   NOR2_X1 i_1679 (.A1(n_3286), .A2(n_3263), .ZN(n_2609));
   NOR2_X1 i_1680 (.A1(n_3286), .A2(n_3262), .ZN(n_2610));
   NOR2_X1 i_1681 (.A1(n_3286), .A2(n_3261), .ZN(n_2611));
   NOR2_X1 i_1682 (.A1(n_3286), .A2(n_3260), .ZN(n_2612));
   NOR2_X1 i_1683 (.A1(n_3286), .A2(n_3259), .ZN(n_2613));
   NOR2_X1 i_1684 (.A1(n_3286), .A2(n_3258), .ZN(n_2614));
   NOR2_X1 i_1685 (.A1(n_3286), .A2(n_3257), .ZN(n_2615));
   NOR2_X1 i_1686 (.A1(n_3286), .A2(n_3256), .ZN(n_2616));
   NOR2_X1 i_1687 (.A1(n_3286), .A2(n_3255), .ZN(n_2617));
   NOR2_X1 i_1688 (.A1(n_3286), .A2(n_3254), .ZN(n_2618));
   NOR2_X1 i_1689 (.A1(n_3286), .A2(n_3253), .ZN(n_2619));
   NOR2_X1 i_1690 (.A1(n_3286), .A2(n_3252), .ZN(n_2620));
   NOR2_X1 i_1691 (.A1(n_3286), .A2(n_3251), .ZN(n_2621));
   NOR2_X1 i_1692 (.A1(n_3286), .A2(n_3250), .ZN(n_2622));
   NOR2_X1 i_1693 (.A1(n_3286), .A2(n_3249), .ZN(n_2623));
   NOR2_X1 i_1694 (.A1(n_3286), .A2(n_3248), .ZN(n_2624));
   NOR2_X1 i_1695 (.A1(n_3286), .A2(n_3247), .ZN(n_2625));
   NOR2_X1 i_1696 (.A1(n_3286), .A2(n_3246), .ZN(n_2626));
   NOR2_X1 i_1697 (.A1(n_3285), .A2(n_3277), .ZN(n_2627));
   NOR2_X1 i_1698 (.A1(n_3285), .A2(n_3276), .ZN(n_2628));
   NOR2_X1 i_1699 (.A1(n_3285), .A2(n_3275), .ZN(n_2629));
   NOR2_X1 i_1700 (.A1(n_3285), .A2(n_3274), .ZN(n_2630));
   NOR2_X1 i_1701 (.A1(n_3285), .A2(n_3273), .ZN(n_2631));
   NOR2_X1 i_1702 (.A1(n_3285), .A2(n_3272), .ZN(n_2632));
   NOR2_X1 i_1703 (.A1(n_3285), .A2(n_3271), .ZN(n_2633));
   NOR2_X1 i_1704 (.A1(n_3285), .A2(n_3270), .ZN(n_2634));
   NOR2_X1 i_1705 (.A1(n_3285), .A2(n_3269), .ZN(n_2635));
   NOR2_X1 i_1706 (.A1(n_3285), .A2(n_3268), .ZN(n_2636));
   NOR2_X1 i_1707 (.A1(n_3285), .A2(n_3267), .ZN(n_2637));
   NOR2_X1 i_1708 (.A1(n_3285), .A2(n_3266), .ZN(n_2638));
   NOR2_X1 i_1709 (.A1(n_3285), .A2(n_3265), .ZN(n_2639));
   NOR2_X1 i_1710 (.A1(n_3285), .A2(n_3264), .ZN(n_2640));
   NOR2_X1 i_1711 (.A1(n_3285), .A2(n_3263), .ZN(n_2641));
   NOR2_X1 i_1712 (.A1(n_3285), .A2(n_3262), .ZN(n_2642));
   NOR2_X1 i_1713 (.A1(n_3285), .A2(n_3261), .ZN(n_2643));
   NOR2_X1 i_1714 (.A1(n_3285), .A2(n_3260), .ZN(n_2644));
   NOR2_X1 i_1715 (.A1(n_3285), .A2(n_3259), .ZN(n_2645));
   NOR2_X1 i_1716 (.A1(n_3285), .A2(n_3258), .ZN(n_2646));
   NOR2_X1 i_1717 (.A1(n_3285), .A2(n_3257), .ZN(n_2647));
   NOR2_X1 i_1718 (.A1(n_3285), .A2(n_3256), .ZN(n_2648));
   NOR2_X1 i_1719 (.A1(n_3285), .A2(n_3255), .ZN(n_2649));
   NOR2_X1 i_1720 (.A1(n_3285), .A2(n_3254), .ZN(n_2650));
   NOR2_X1 i_1721 (.A1(n_3285), .A2(n_3253), .ZN(n_2651));
   NOR2_X1 i_1722 (.A1(n_3285), .A2(n_3252), .ZN(n_2652));
   NOR2_X1 i_1723 (.A1(n_3285), .A2(n_3251), .ZN(n_2653));
   NOR2_X1 i_1724 (.A1(n_3285), .A2(n_3250), .ZN(n_2654));
   NOR2_X1 i_1725 (.A1(n_3285), .A2(n_3249), .ZN(n_2655));
   NOR2_X1 i_1726 (.A1(n_3285), .A2(n_3248), .ZN(n_2656));
   NOR2_X1 i_1727 (.A1(n_3285), .A2(n_3247), .ZN(n_2657));
   NOR2_X1 i_1728 (.A1(n_3285), .A2(n_3246), .ZN(n_2658));
   NOR2_X1 i_1729 (.A1(n_3284), .A2(n_3277), .ZN(n_2659));
   NOR2_X1 i_1730 (.A1(n_3284), .A2(n_3276), .ZN(n_2660));
   NOR2_X1 i_1731 (.A1(n_3284), .A2(n_3275), .ZN(n_2661));
   NOR2_X1 i_1732 (.A1(n_3284), .A2(n_3274), .ZN(n_2662));
   NOR2_X1 i_1733 (.A1(n_3284), .A2(n_3273), .ZN(n_2663));
   NOR2_X1 i_1734 (.A1(n_3284), .A2(n_3272), .ZN(n_2664));
   NOR2_X1 i_1735 (.A1(n_3284), .A2(n_3271), .ZN(n_2665));
   NOR2_X1 i_1736 (.A1(n_3284), .A2(n_3270), .ZN(n_2666));
   NOR2_X1 i_1737 (.A1(n_3284), .A2(n_3269), .ZN(n_2667));
   NOR2_X1 i_1738 (.A1(n_3284), .A2(n_3268), .ZN(n_2668));
   NOR2_X1 i_1739 (.A1(n_3284), .A2(n_3267), .ZN(n_2669));
   NOR2_X1 i_1740 (.A1(n_3284), .A2(n_3266), .ZN(n_2670));
   NOR2_X1 i_1741 (.A1(n_3284), .A2(n_3265), .ZN(n_2671));
   NOR2_X1 i_1742 (.A1(n_3284), .A2(n_3264), .ZN(n_2672));
   NOR2_X1 i_1743 (.A1(n_3284), .A2(n_3263), .ZN(n_2673));
   NOR2_X1 i_1744 (.A1(n_3284), .A2(n_3262), .ZN(n_2674));
   NOR2_X1 i_1745 (.A1(n_3284), .A2(n_3261), .ZN(n_2675));
   NOR2_X1 i_1746 (.A1(n_3284), .A2(n_3260), .ZN(n_2676));
   NOR2_X1 i_1747 (.A1(n_3284), .A2(n_3259), .ZN(n_2677));
   NOR2_X1 i_1748 (.A1(n_3284), .A2(n_3258), .ZN(n_2678));
   NOR2_X1 i_1749 (.A1(n_3284), .A2(n_3257), .ZN(n_2679));
   NOR2_X1 i_1750 (.A1(n_3284), .A2(n_3256), .ZN(n_2680));
   NOR2_X1 i_1751 (.A1(n_3284), .A2(n_3255), .ZN(n_2681));
   NOR2_X1 i_1752 (.A1(n_3284), .A2(n_3254), .ZN(n_2682));
   NOR2_X1 i_1753 (.A1(n_3284), .A2(n_3253), .ZN(n_2683));
   NOR2_X1 i_1754 (.A1(n_3284), .A2(n_3252), .ZN(n_2684));
   NOR2_X1 i_1755 (.A1(n_3284), .A2(n_3251), .ZN(n_2685));
   NOR2_X1 i_1756 (.A1(n_3284), .A2(n_3250), .ZN(n_2686));
   NOR2_X1 i_1757 (.A1(n_3284), .A2(n_3249), .ZN(n_2687));
   NOR2_X1 i_1758 (.A1(n_3284), .A2(n_3248), .ZN(n_2688));
   NOR2_X1 i_1759 (.A1(n_3284), .A2(n_3247), .ZN(n_2689));
   NOR2_X1 i_1760 (.A1(n_3284), .A2(n_3246), .ZN(n_2690));
   NOR2_X1 i_1761 (.A1(n_3283), .A2(n_3277), .ZN(n_2691));
   NOR2_X1 i_1762 (.A1(n_3283), .A2(n_3276), .ZN(n_2692));
   NOR2_X1 i_1763 (.A1(n_3283), .A2(n_3275), .ZN(n_2693));
   NOR2_X1 i_1764 (.A1(n_3283), .A2(n_3274), .ZN(n_2694));
   NOR2_X1 i_1765 (.A1(n_3283), .A2(n_3273), .ZN(n_2695));
   NOR2_X1 i_1766 (.A1(n_3283), .A2(n_3272), .ZN(n_2696));
   NOR2_X1 i_1767 (.A1(n_3283), .A2(n_3271), .ZN(n_2697));
   NOR2_X1 i_1768 (.A1(n_3283), .A2(n_3270), .ZN(n_2698));
   NOR2_X1 i_1769 (.A1(n_3283), .A2(n_3269), .ZN(n_2699));
   NOR2_X1 i_1770 (.A1(n_3283), .A2(n_3268), .ZN(n_2700));
   NOR2_X1 i_1771 (.A1(n_3283), .A2(n_3267), .ZN(n_2701));
   NOR2_X1 i_1772 (.A1(n_3283), .A2(n_3266), .ZN(n_2702));
   NOR2_X1 i_1773 (.A1(n_3283), .A2(n_3265), .ZN(n_2703));
   NOR2_X1 i_1774 (.A1(n_3283), .A2(n_3264), .ZN(n_2704));
   NOR2_X1 i_1775 (.A1(n_3283), .A2(n_3263), .ZN(n_2705));
   NOR2_X1 i_1776 (.A1(n_3283), .A2(n_3262), .ZN(n_2706));
   NOR2_X1 i_1777 (.A1(n_3283), .A2(n_3261), .ZN(n_2707));
   NOR2_X1 i_1778 (.A1(n_3283), .A2(n_3260), .ZN(n_2708));
   NOR2_X1 i_1779 (.A1(n_3283), .A2(n_3259), .ZN(n_2709));
   NOR2_X1 i_1780 (.A1(n_3283), .A2(n_3258), .ZN(n_2710));
   NOR2_X1 i_1781 (.A1(n_3283), .A2(n_3257), .ZN(n_2711));
   NOR2_X1 i_1782 (.A1(n_3283), .A2(n_3256), .ZN(n_2712));
   NOR2_X1 i_1783 (.A1(n_3283), .A2(n_3255), .ZN(n_2713));
   NOR2_X1 i_1784 (.A1(n_3283), .A2(n_3254), .ZN(n_2714));
   NOR2_X1 i_1785 (.A1(n_3283), .A2(n_3253), .ZN(n_2715));
   NOR2_X1 i_1786 (.A1(n_3283), .A2(n_3252), .ZN(n_2716));
   NOR2_X1 i_1787 (.A1(n_3283), .A2(n_3251), .ZN(n_2717));
   NOR2_X1 i_1788 (.A1(n_3283), .A2(n_3250), .ZN(n_2718));
   NOR2_X1 i_1789 (.A1(n_3283), .A2(n_3249), .ZN(n_2719));
   NOR2_X1 i_1790 (.A1(n_3283), .A2(n_3248), .ZN(n_2720));
   NOR2_X1 i_1791 (.A1(n_3283), .A2(n_3247), .ZN(n_2721));
   NOR2_X1 i_1792 (.A1(n_3283), .A2(n_3246), .ZN(n_2722));
   NOR2_X1 i_1793 (.A1(n_3282), .A2(n_3277), .ZN(n_2723));
   NOR2_X1 i_1794 (.A1(n_3282), .A2(n_3276), .ZN(n_2724));
   NOR2_X1 i_1795 (.A1(n_3282), .A2(n_3275), .ZN(n_2725));
   NOR2_X1 i_1796 (.A1(n_3282), .A2(n_3274), .ZN(n_2726));
   NOR2_X1 i_1797 (.A1(n_3282), .A2(n_3273), .ZN(n_2727));
   NOR2_X1 i_1798 (.A1(n_3282), .A2(n_3272), .ZN(n_2728));
   NOR2_X1 i_1799 (.A1(n_3282), .A2(n_3271), .ZN(n_2729));
   NOR2_X1 i_1800 (.A1(n_3282), .A2(n_3270), .ZN(n_2730));
   NOR2_X1 i_1801 (.A1(n_3282), .A2(n_3269), .ZN(n_2731));
   NOR2_X1 i_1802 (.A1(n_3282), .A2(n_3268), .ZN(n_2732));
   NOR2_X1 i_1803 (.A1(n_3282), .A2(n_3267), .ZN(n_2733));
   NOR2_X1 i_1804 (.A1(n_3282), .A2(n_3266), .ZN(n_2734));
   NOR2_X1 i_1805 (.A1(n_3282), .A2(n_3265), .ZN(n_2735));
   NOR2_X1 i_1806 (.A1(n_3282), .A2(n_3264), .ZN(n_2736));
   NOR2_X1 i_1807 (.A1(n_3282), .A2(n_3263), .ZN(n_2737));
   NOR2_X1 i_1808 (.A1(n_3282), .A2(n_3262), .ZN(n_2738));
   NOR2_X1 i_1809 (.A1(n_3282), .A2(n_3261), .ZN(n_2739));
   NOR2_X1 i_1810 (.A1(n_3282), .A2(n_3260), .ZN(n_2740));
   NOR2_X1 i_1811 (.A1(n_3282), .A2(n_3259), .ZN(n_2741));
   NOR2_X1 i_1812 (.A1(n_3282), .A2(n_3258), .ZN(n_2742));
   NOR2_X1 i_1813 (.A1(n_3282), .A2(n_3257), .ZN(n_2743));
   NOR2_X1 i_1814 (.A1(n_3282), .A2(n_3256), .ZN(n_2744));
   NOR2_X1 i_1815 (.A1(n_3282), .A2(n_3255), .ZN(n_2745));
   NOR2_X1 i_1816 (.A1(n_3282), .A2(n_3254), .ZN(n_2746));
   NOR2_X1 i_1817 (.A1(n_3282), .A2(n_3253), .ZN(n_2747));
   NOR2_X1 i_1818 (.A1(n_3282), .A2(n_3252), .ZN(n_2748));
   NOR2_X1 i_1819 (.A1(n_3282), .A2(n_3251), .ZN(n_2749));
   NOR2_X1 i_1820 (.A1(n_3282), .A2(n_3250), .ZN(n_2750));
   NOR2_X1 i_1821 (.A1(n_3282), .A2(n_3249), .ZN(n_2751));
   NOR2_X1 i_1822 (.A1(n_3282), .A2(n_3248), .ZN(n_2752));
   NOR2_X1 i_1823 (.A1(n_3282), .A2(n_3247), .ZN(n_2753));
   NOR2_X1 i_1824 (.A1(n_3282), .A2(n_3246), .ZN(n_2754));
   NOR2_X1 i_1825 (.A1(n_3281), .A2(n_3277), .ZN(n_2755));
   NOR2_X1 i_1826 (.A1(n_3281), .A2(n_3276), .ZN(n_2756));
   NOR2_X1 i_1827 (.A1(n_3281), .A2(n_3275), .ZN(n_2757));
   NOR2_X1 i_1828 (.A1(n_3281), .A2(n_3274), .ZN(n_2758));
   NOR2_X1 i_1829 (.A1(n_3281), .A2(n_3273), .ZN(n_2759));
   NOR2_X1 i_1830 (.A1(n_3281), .A2(n_3272), .ZN(n_2760));
   NOR2_X1 i_1831 (.A1(n_3281), .A2(n_3271), .ZN(n_2761));
   NOR2_X1 i_1832 (.A1(n_3281), .A2(n_3270), .ZN(n_2762));
   NOR2_X1 i_1833 (.A1(n_3281), .A2(n_3269), .ZN(n_2763));
   NOR2_X1 i_1834 (.A1(n_3281), .A2(n_3268), .ZN(n_2764));
   NOR2_X1 i_1835 (.A1(n_3281), .A2(n_3267), .ZN(n_2765));
   NOR2_X1 i_1836 (.A1(n_3281), .A2(n_3266), .ZN(n_2766));
   NOR2_X1 i_1837 (.A1(n_3281), .A2(n_3265), .ZN(n_2767));
   NOR2_X1 i_1838 (.A1(n_3281), .A2(n_3264), .ZN(n_2768));
   NOR2_X1 i_1839 (.A1(n_3281), .A2(n_3263), .ZN(n_2769));
   NOR2_X1 i_1840 (.A1(n_3281), .A2(n_3262), .ZN(n_2770));
   NOR2_X1 i_1841 (.A1(n_3281), .A2(n_3261), .ZN(n_2771));
   NOR2_X1 i_1842 (.A1(n_3281), .A2(n_3260), .ZN(n_2772));
   NOR2_X1 i_1843 (.A1(n_3281), .A2(n_3259), .ZN(n_2773));
   NOR2_X1 i_1844 (.A1(n_3281), .A2(n_3258), .ZN(n_2774));
   NOR2_X1 i_1845 (.A1(n_3281), .A2(n_3257), .ZN(n_2775));
   NOR2_X1 i_1846 (.A1(n_3281), .A2(n_3256), .ZN(n_2776));
   NOR2_X1 i_1847 (.A1(n_3281), .A2(n_3255), .ZN(n_2777));
   NOR2_X1 i_1848 (.A1(n_3281), .A2(n_3254), .ZN(n_2778));
   NOR2_X1 i_1849 (.A1(n_3281), .A2(n_3253), .ZN(n_2779));
   NOR2_X1 i_1850 (.A1(n_3281), .A2(n_3252), .ZN(n_2780));
   NOR2_X1 i_1851 (.A1(n_3281), .A2(n_3251), .ZN(n_2781));
   NOR2_X1 i_1852 (.A1(n_3281), .A2(n_3250), .ZN(n_2782));
   NOR2_X1 i_1853 (.A1(n_3281), .A2(n_3249), .ZN(n_2783));
   NOR2_X1 i_1854 (.A1(n_3281), .A2(n_3248), .ZN(n_2784));
   NOR2_X1 i_1855 (.A1(n_3281), .A2(n_3247), .ZN(n_2785));
   NOR2_X1 i_1856 (.A1(n_3281), .A2(n_3246), .ZN(n_2786));
   NOR2_X1 i_1857 (.A1(n_3280), .A2(n_3277), .ZN(n_2787));
   NOR2_X1 i_1858 (.A1(n_3280), .A2(n_3276), .ZN(n_2788));
   NOR2_X1 i_1859 (.A1(n_3280), .A2(n_3275), .ZN(n_2789));
   NOR2_X1 i_1860 (.A1(n_3280), .A2(n_3274), .ZN(n_2790));
   NOR2_X1 i_1861 (.A1(n_3280), .A2(n_3273), .ZN(n_2791));
   NOR2_X1 i_1862 (.A1(n_3280), .A2(n_3272), .ZN(n_2792));
   NOR2_X1 i_1863 (.A1(n_3280), .A2(n_3271), .ZN(n_2793));
   NOR2_X1 i_1864 (.A1(n_3280), .A2(n_3270), .ZN(n_2794));
   NOR2_X1 i_1865 (.A1(n_3280), .A2(n_3269), .ZN(n_2795));
   NOR2_X1 i_1866 (.A1(n_3280), .A2(n_3268), .ZN(n_2796));
   NOR2_X1 i_1867 (.A1(n_3280), .A2(n_3267), .ZN(n_2797));
   NOR2_X1 i_1868 (.A1(n_3280), .A2(n_3266), .ZN(n_2798));
   NOR2_X1 i_1869 (.A1(n_3280), .A2(n_3265), .ZN(n_2799));
   NOR2_X1 i_1870 (.A1(n_3280), .A2(n_3264), .ZN(n_2800));
   NOR2_X1 i_1871 (.A1(n_3280), .A2(n_3263), .ZN(n_2801));
   NOR2_X1 i_1872 (.A1(n_3280), .A2(n_3262), .ZN(n_2802));
   NOR2_X1 i_1873 (.A1(n_3280), .A2(n_3261), .ZN(n_2803));
   NOR2_X1 i_1874 (.A1(n_3280), .A2(n_3260), .ZN(n_2804));
   NOR2_X1 i_1875 (.A1(n_3280), .A2(n_3259), .ZN(n_2805));
   NOR2_X1 i_1876 (.A1(n_3280), .A2(n_3258), .ZN(n_2806));
   NOR2_X1 i_1877 (.A1(n_3280), .A2(n_3257), .ZN(n_2807));
   NOR2_X1 i_1878 (.A1(n_3280), .A2(n_3256), .ZN(n_2808));
   NOR2_X1 i_1879 (.A1(n_3280), .A2(n_3255), .ZN(n_2809));
   NOR2_X1 i_1880 (.A1(n_3280), .A2(n_3254), .ZN(n_2810));
   NOR2_X1 i_1881 (.A1(n_3280), .A2(n_3253), .ZN(n_2811));
   NOR2_X1 i_1882 (.A1(n_3280), .A2(n_3252), .ZN(n_2812));
   NOR2_X1 i_1883 (.A1(n_3280), .A2(n_3251), .ZN(n_2813));
   NOR2_X1 i_1884 (.A1(n_3280), .A2(n_3250), .ZN(n_2814));
   NOR2_X1 i_1885 (.A1(n_3280), .A2(n_3249), .ZN(n_2815));
   NOR2_X1 i_1886 (.A1(n_3280), .A2(n_3248), .ZN(n_2816));
   NOR2_X1 i_1887 (.A1(n_3280), .A2(n_3247), .ZN(n_2817));
   NOR2_X1 i_1888 (.A1(n_3280), .A2(n_3246), .ZN(n_2818));
   NOR2_X1 i_1889 (.A1(n_3279), .A2(n_3277), .ZN(n_2819));
   NOR2_X1 i_1890 (.A1(n_3279), .A2(n_3276), .ZN(n_2820));
   NOR2_X1 i_1891 (.A1(n_3279), .A2(n_3275), .ZN(n_2821));
   NOR2_X1 i_1892 (.A1(n_3279), .A2(n_3274), .ZN(n_2822));
   NOR2_X1 i_1893 (.A1(n_3279), .A2(n_3273), .ZN(n_2823));
   NOR2_X1 i_1894 (.A1(n_3279), .A2(n_3272), .ZN(n_2824));
   NOR2_X1 i_1895 (.A1(n_3279), .A2(n_3271), .ZN(n_2825));
   NOR2_X1 i_1896 (.A1(n_3279), .A2(n_3270), .ZN(n_2826));
   NOR2_X1 i_1897 (.A1(n_3279), .A2(n_3269), .ZN(n_2827));
   NOR2_X1 i_1898 (.A1(n_3279), .A2(n_3268), .ZN(n_2828));
   NOR2_X1 i_1899 (.A1(n_3279), .A2(n_3267), .ZN(n_2829));
   NOR2_X1 i_1900 (.A1(n_3279), .A2(n_3266), .ZN(n_2830));
   NOR2_X1 i_1901 (.A1(n_3279), .A2(n_3265), .ZN(n_2831));
   NOR2_X1 i_1902 (.A1(n_3279), .A2(n_3264), .ZN(n_2832));
   NOR2_X1 i_1903 (.A1(n_3279), .A2(n_3263), .ZN(n_2833));
   NOR2_X1 i_1904 (.A1(n_3279), .A2(n_3262), .ZN(n_2834));
   NOR2_X1 i_1905 (.A1(n_3279), .A2(n_3261), .ZN(n_2835));
   NOR2_X1 i_1906 (.A1(n_3279), .A2(n_3260), .ZN(n_2836));
   NOR2_X1 i_1907 (.A1(n_3279), .A2(n_3259), .ZN(n_2837));
   NOR2_X1 i_1908 (.A1(n_3279), .A2(n_3258), .ZN(n_2838));
   NOR2_X1 i_1909 (.A1(n_3279), .A2(n_3257), .ZN(n_2839));
   NOR2_X1 i_1910 (.A1(n_3279), .A2(n_3256), .ZN(n_2840));
   NOR2_X1 i_1911 (.A1(n_3279), .A2(n_3255), .ZN(n_2841));
   NOR2_X1 i_1912 (.A1(n_3279), .A2(n_3254), .ZN(n_2842));
   NOR2_X1 i_1913 (.A1(n_3279), .A2(n_3253), .ZN(n_2843));
   NOR2_X1 i_1914 (.A1(n_3279), .A2(n_3252), .ZN(n_2844));
   NOR2_X1 i_1915 (.A1(n_3279), .A2(n_3251), .ZN(n_2845));
   NOR2_X1 i_1916 (.A1(n_3279), .A2(n_3250), .ZN(n_2846));
   NOR2_X1 i_1917 (.A1(n_3279), .A2(n_3249), .ZN(n_2847));
   NOR2_X1 i_1918 (.A1(n_3279), .A2(n_3248), .ZN(n_2848));
   NOR2_X1 i_1919 (.A1(n_3278), .A2(n_3277), .ZN(n_2849));
   NOR2_X1 i_1920 (.A1(n_3278), .A2(n_3276), .ZN(n_2850));
   NOR2_X1 i_1921 (.A1(n_3278), .A2(n_3275), .ZN(n_2851));
   NOR2_X1 i_1922 (.A1(n_3278), .A2(n_3274), .ZN(n_2852));
   NOR2_X1 i_1923 (.A1(n_3278), .A2(n_3273), .ZN(n_2853));
   NOR2_X1 i_1924 (.A1(n_3278), .A2(n_3272), .ZN(n_2854));
   NOR2_X1 i_1925 (.A1(n_3278), .A2(n_3271), .ZN(n_2855));
   NOR2_X1 i_1926 (.A1(n_3278), .A2(n_3270), .ZN(n_2856));
   NOR2_X1 i_1927 (.A1(n_3278), .A2(n_3269), .ZN(n_2857));
   NOR2_X1 i_1928 (.A1(n_3278), .A2(n_3268), .ZN(n_2858));
   NOR2_X1 i_1929 (.A1(n_3278), .A2(n_3267), .ZN(n_2859));
   NOR2_X1 i_1930 (.A1(n_3278), .A2(n_3266), .ZN(n_2860));
   NOR2_X1 i_1931 (.A1(n_3278), .A2(n_3265), .ZN(n_2861));
   NOR2_X1 i_1932 (.A1(n_3278), .A2(n_3264), .ZN(n_2862));
   NOR2_X1 i_1933 (.A1(n_3278), .A2(n_3263), .ZN(n_2863));
   NOR2_X1 i_1934 (.A1(n_3278), .A2(n_3262), .ZN(n_2864));
   NOR2_X1 i_1935 (.A1(n_3278), .A2(n_3261), .ZN(n_2865));
   NOR2_X1 i_1936 (.A1(n_3278), .A2(n_3260), .ZN(n_2866));
   NOR2_X1 i_1937 (.A1(n_3278), .A2(n_3259), .ZN(n_2867));
   NOR2_X1 i_1938 (.A1(n_3278), .A2(n_3258), .ZN(n_2868));
   NOR2_X1 i_1939 (.A1(n_3278), .A2(n_3257), .ZN(n_2869));
   NOR2_X1 i_1940 (.A1(n_3278), .A2(n_3256), .ZN(n_2870));
   NOR2_X1 i_1941 (.A1(n_3278), .A2(n_3255), .ZN(n_2871));
   NOR2_X1 i_1942 (.A1(n_3278), .A2(n_3254), .ZN(n_2872));
   NOR2_X1 i_1943 (.A1(n_3278), .A2(n_3253), .ZN(n_2873));
   NOR2_X1 i_1944 (.A1(n_3278), .A2(n_3252), .ZN(n_2874));
   NOR2_X1 i_1945 (.A1(n_3278), .A2(n_3251), .ZN(n_2875));
   NOR2_X1 i_1946 (.A1(n_3278), .A2(n_3250), .ZN(n_2876));
   NOR2_X1 i_1947 (.A1(n_3278), .A2(n_3249), .ZN(n_2877));
   INV_X1 i_1948 (.A(n_2878), .ZN(p_0[1]));
   OAI21_X1 i_1949 (.A(n_3230), .B1(n_3233), .B2(n_3232), .ZN(n_2878));
   XOR2_X1 i_1950 (.A(n_3230), .B(n_2879), .Z(p_0[2]));
   OAI21_X1 i_1951 (.A(n_3229), .B1(n_0), .B2(n_3235), .ZN(n_2879));
   XNOR2_X1 i_1952 (.A(n_3228), .B(n_2880), .ZN(p_0[3]));
   OAI21_X1 i_1953 (.A(n_3236), .B1(n_2), .B2(n_4), .ZN(n_2880));
   XOR2_X1 i_1954 (.A(n_3226), .B(n_2881), .Z(p_0[4]));
   XOR2_X1 i_1955 (.A(n_6), .B(n_10), .Z(n_2881));
   XOR2_X1 i_1956 (.A(n_3225), .B(n_2888), .Z(p_0[5]));
   XOR2_X1 i_1957 (.A(n_2887), .B(n_2884), .Z(p_0[6]));
   XOR2_X1 i_1958 (.A(n_2885), .B(n_2882), .Z(p_0[7]));
   NOR2_X1 i_1959 (.A1(n_3222), .A2(n_3213), .ZN(n_2882));
   XNOR2_X1 i_1960 (.A(n_2889), .B(n_2883), .ZN(p_0[8]));
   OAI22_X1 i_1961 (.A1(n_38), .A2(n_40), .B1(n_3213), .B2(n_2885), .ZN(n_2883));
   AOI21_X1 i_1962 (.A(n_3223), .B1(n_26), .B2(n_28), .ZN(n_2884));
   AOI21_X1 i_1963 (.A(n_3223), .B1(n_3217), .B2(n_2886), .ZN(n_2885));
   INV_X1 i_1964 (.A(n_2887), .ZN(n_2886));
   AOI21_X1 i_1965 (.A(n_3220), .B1(n_3225), .B2(n_3218), .ZN(n_2887));
   OAI21_X1 i_1966 (.A(n_3218), .B1(n_16), .B2(n_18), .ZN(n_2888));
   NOR2_X1 i_1967 (.A1(n_3224), .A2(n_3215), .ZN(n_2889));
   XOR2_X1 i_1968 (.A(n_3211), .B(n_2896), .Z(p_0[9]));
   XOR2_X1 i_1969 (.A(n_2895), .B(n_2892), .Z(p_0[10]));
   XOR2_X1 i_1970 (.A(n_2893), .B(n_2890), .Z(p_0[11]));
   NOR2_X1 i_1971 (.A1(n_3208), .A2(n_3199), .ZN(n_2890));
   XNOR2_X1 i_1972 (.A(n_2897), .B(n_2891), .ZN(p_0[12]));
   OAI22_X1 i_1973 (.A1(n_106), .A2(n_108), .B1(n_3199), .B2(n_2893), .ZN(n_2891));
   AOI21_X1 i_1974 (.A(n_3209), .B1(n_86), .B2(n_88), .ZN(n_2892));
   AOI21_X1 i_1975 (.A(n_3209), .B1(n_3203), .B2(n_2894), .ZN(n_2893));
   INV_X1 i_1976 (.A(n_2895), .ZN(n_2894));
   AOI21_X1 i_1977 (.A(n_3206), .B1(n_3211), .B2(n_3204), .ZN(n_2895));
   OAI21_X1 i_1978 (.A(n_3204), .B1(n_68), .B2(n_70), .ZN(n_2896));
   NOR2_X1 i_1979 (.A1(n_3210), .A2(n_3201), .ZN(n_2897));
   XOR2_X1 i_1980 (.A(n_3197), .B(n_2904), .Z(p_0[13]));
   XOR2_X1 i_1981 (.A(n_2903), .B(n_2900), .Z(p_0[14]));
   XOR2_X1 i_1982 (.A(n_2901), .B(n_2898), .Z(p_0[15]));
   NOR2_X1 i_1983 (.A1(n_3194), .A2(n_3185), .ZN(n_2898));
   XNOR2_X1 i_1984 (.A(n_2905), .B(n_2899), .ZN(p_0[16]));
   OAI22_X1 i_1985 (.A1(n_206), .A2(n_208), .B1(n_3185), .B2(n_2901), .ZN(n_2899));
   AOI21_X1 i_1986 (.A(n_3195), .B1(n_178), .B2(n_180), .ZN(n_2900));
   AOI21_X1 i_1987 (.A(n_3195), .B1(n_3189), .B2(n_2902), .ZN(n_2901));
   INV_X1 i_1988 (.A(n_2903), .ZN(n_2902));
   AOI21_X1 i_1989 (.A(n_3192), .B1(n_3197), .B2(n_3190), .ZN(n_2903));
   OAI21_X1 i_1990 (.A(n_3190), .B1(n_152), .B2(n_154), .ZN(n_2904));
   NOR2_X1 i_1991 (.A1(n_3196), .A2(n_3187), .ZN(n_2905));
   XOR2_X1 i_1992 (.A(n_3183), .B(n_2912), .Z(p_0[17]));
   XOR2_X1 i_1993 (.A(n_2911), .B(n_2908), .Z(p_0[18]));
   XOR2_X1 i_1994 (.A(n_2909), .B(n_2906), .Z(p_0[19]));
   NOR2_X1 i_1995 (.A1(n_3149), .A2(n_3139), .ZN(n_2906));
   XNOR2_X1 i_1996 (.A(n_2913), .B(n_2907), .ZN(p_0[20]));
   OAI21_X1 i_1997 (.A(n_3148), .B1(n_3139), .B2(n_2909), .ZN(n_2907));
   NOR2_X1 i_1998 (.A1(n_3151), .A2(n_3141), .ZN(n_2908));
   INV_X1 i_1999 (.A(n_2910), .ZN(n_2909));
   OAI21_X1 i_2000 (.A(n_3150), .B1(n_3141), .B2(n_2911), .ZN(n_2910));
   AOI21_X1 i_2001 (.A(n_3146), .B1(n_3183), .B2(n_3143), .ZN(n_2911));
   OAI21_X1 i_2002 (.A(n_3143), .B1(n_268), .B2(n_270), .ZN(n_2912));
   AOI21_X1 i_2003 (.A(n_3153), .B1(n_376), .B2(n_378), .ZN(n_2913));
   XOR2_X1 i_2004 (.A(n_2941), .B(n_2920), .Z(p_0[21]));
   XOR2_X1 i_2005 (.A(n_2919), .B(n_2916), .Z(p_0[22]));
   XOR2_X1 i_2006 (.A(n_2917), .B(n_2914), .Z(p_0[23]));
   NOR2_X1 i_2007 (.A1(n_3177), .A2(n_3121), .ZN(n_2914));
   XNOR2_X1 i_2008 (.A(n_2921), .B(n_2915), .ZN(p_0[24]));
   OAI21_X1 i_2009 (.A(n_3176), .B1(n_3121), .B2(n_2917), .ZN(n_2915));
   NOR2_X1 i_2010 (.A1(n_3179), .A2(n_3123), .ZN(n_2916));
   INV_X1 i_2011 (.A(n_2918), .ZN(n_2917));
   OAI21_X1 i_2012 (.A(n_3178), .B1(n_3123), .B2(n_2919), .ZN(n_2918));
   AOI21_X1 i_2013 (.A(n_3182), .B1(n_3125), .B2(n_2941), .ZN(n_2919));
   OAI21_X1 i_2014 (.A(n_3125), .B1(n_379), .B2(n_418), .ZN(n_2920));
   AOI21_X1 i_2015 (.A(n_3181), .B1(n_505), .B2(n_550), .ZN(n_2921));
   XOR2_X1 i_2016 (.A(n_2939), .B(n_2928), .Z(p_0[25]));
   XOR2_X1 i_2017 (.A(n_2927), .B(n_2924), .Z(p_0[26]));
   XOR2_X1 i_2018 (.A(n_2925), .B(n_2922), .Z(p_0[27]));
   NOR2_X1 i_2019 (.A1(n_3160), .A2(n_3133), .ZN(n_2922));
   XNOR2_X1 i_2020 (.A(n_2929), .B(n_2923), .ZN(p_0[28]));
   OAI21_X1 i_2021 (.A(n_3159), .B1(n_3133), .B2(n_2925), .ZN(n_2923));
   NOR2_X1 i_2022 (.A1(n_3162), .A2(n_3135), .ZN(n_2924));
   INV_X1 i_2023 (.A(n_2926), .ZN(n_2925));
   OAI21_X1 i_2024 (.A(n_3161), .B1(n_3135), .B2(n_2927), .ZN(n_2926));
   AOI21_X1 i_2025 (.A(n_3157), .B1(n_3137), .B2(n_2939), .ZN(n_2927));
   OAI21_X1 i_2026 (.A(n_3137), .B1(n_596), .B2(n_598), .ZN(n_2928));
   AOI21_X1 i_2027 (.A(n_3164), .B1(n_701), .B2(n_754), .ZN(n_2929));
   XOR2_X1 i_2028 (.A(n_2937), .B(n_2936), .Z(p_0[29]));
   XOR2_X1 i_2029 (.A(n_2935), .B(n_2932), .Z(p_0[30]));
   XOR2_X1 i_2030 (.A(n_2933), .B(n_2930), .Z(p_0[31]));
   NOR2_X1 i_2031 (.A1(n_3169), .A2(n_3127), .ZN(n_2930));
   XOR2_X1 i_2032 (.A(n_2943), .B(n_2931), .Z(p_0[32]));
   OAI21_X1 i_2033 (.A(n_3168), .B1(n_3127), .B2(n_2933), .ZN(n_2931));
   NOR2_X1 i_2034 (.A1(n_3171), .A2(n_3130), .ZN(n_2932));
   INV_X1 i_2035 (.A(n_2934), .ZN(n_2933));
   OAI21_X1 i_2036 (.A(n_3170), .B1(n_3130), .B2(n_2935), .ZN(n_2934));
   AOI21_X1 i_2037 (.A(n_3166), .B1(n_3131), .B2(n_2937), .ZN(n_2935));
   OAI21_X1 i_2038 (.A(n_3131), .B1(n_755), .B2(n_810), .ZN(n_2936));
   INV_X1 i_2039 (.A(n_2938), .ZN(n_2937));
   OAI21_X1 i_2040 (.A(n_3132), .B1(n_3156), .B2(n_2939), .ZN(n_2938));
   INV_X1 i_2041 (.A(n_2940), .ZN(n_2939));
   OAI21_X1 i_2042 (.A(n_3120), .B1(n_3174), .B2(n_2941), .ZN(n_2940));
   INV_X1 i_2043 (.A(n_2942), .ZN(n_2941));
   OAI21_X1 i_2044 (.A(n_3138), .B1(n_3183), .B2(n_3145), .ZN(n_2942));
   OAI21_X1 i_2045 (.A(n_3172), .B1(n_3245), .B2(n_3244), .ZN(n_2943));
   XOR2_X1 i_2046 (.A(n_3118), .B(n_2950), .Z(p_0[33]));
   XOR2_X1 i_2047 (.A(n_2949), .B(n_2946), .Z(p_0[34]));
   XOR2_X1 i_2048 (.A(n_2947), .B(n_2944), .Z(p_0[35]));
   NOR2_X1 i_2049 (.A1(n_3087), .A2(n_3077), .ZN(n_2944));
   XNOR2_X1 i_2050 (.A(n_2951), .B(n_2945), .ZN(p_0[36]));
   OAI21_X1 i_2051 (.A(n_3086), .B1(n_3077), .B2(n_2947), .ZN(n_2945));
   NOR2_X1 i_2052 (.A1(n_3089), .A2(n_3079), .ZN(n_2946));
   INV_X1 i_2053 (.A(n_2948), .ZN(n_2947));
   OAI21_X1 i_2054 (.A(n_3088), .B1(n_3079), .B2(n_2949), .ZN(n_2948));
   AOI21_X1 i_2055 (.A(n_3084), .B1(n_3118), .B2(n_3081), .ZN(n_2949));
   OAI21_X1 i_2056 (.A(n_3081), .B1(n_989), .B2(n_1046), .ZN(n_2950));
   AOI21_X1 i_2057 (.A(n_3091), .B1(n_1157), .B2(n_1208), .ZN(n_2951));
   XOR2_X1 i_2058 (.A(n_2979), .B(n_2958), .Z(p_0[37]));
   XOR2_X1 i_2059 (.A(n_2957), .B(n_2954), .Z(p_0[38]));
   XOR2_X1 i_2060 (.A(n_2955), .B(n_2952), .Z(p_0[39]));
   NOR2_X1 i_2061 (.A1(n_3112), .A2(n_3070), .ZN(n_2952));
   XNOR2_X1 i_2062 (.A(n_2959), .B(n_2953), .ZN(p_0[40]));
   OAI21_X1 i_2063 (.A(n_3111), .B1(n_3070), .B2(n_2955), .ZN(n_2953));
   NOR2_X1 i_2064 (.A1(n_3114), .A2(n_3072), .ZN(n_2954));
   INV_X1 i_2065 (.A(n_2956), .ZN(n_2955));
   OAI21_X1 i_2066 (.A(n_3113), .B1(n_3072), .B2(n_2957), .ZN(n_2956));
   AOI21_X1 i_2067 (.A(n_3117), .B1(n_3074), .B2(n_2979), .ZN(n_2957));
   OAI21_X1 i_2068 (.A(n_3074), .B1(n_1209), .B2(n_1258), .ZN(n_2958));
   AOI21_X1 i_2069 (.A(n_3116), .B1(n_1353), .B2(n_1396), .ZN(n_2959));
   XOR2_X1 i_2070 (.A(n_2977), .B(n_2966), .Z(p_0[41]));
   XOR2_X1 i_2071 (.A(n_2965), .B(n_2962), .Z(p_0[42]));
   XOR2_X1 i_2072 (.A(n_2963), .B(n_2960), .Z(p_0[43]));
   NOR2_X1 i_2073 (.A1(n_3098), .A2(n_3056), .ZN(n_2960));
   XNOR2_X1 i_2074 (.A(n_2967), .B(n_2961), .ZN(p_0[44]));
   OAI21_X1 i_2075 (.A(n_3097), .B1(n_3056), .B2(n_2963), .ZN(n_2961));
   NOR2_X1 i_2076 (.A1(n_3100), .A2(n_3058), .ZN(n_2962));
   INV_X1 i_2077 (.A(n_2964), .ZN(n_2963));
   OAI21_X1 i_2078 (.A(n_3099), .B1(n_3058), .B2(n_2965), .ZN(n_2964));
   AOI21_X1 i_2079 (.A(n_3095), .B1(n_3060), .B2(n_2977), .ZN(n_2965));
   OAI21_X1 i_2080 (.A(n_3060), .B1(n_1397), .B2(n_1438), .ZN(n_2966));
   AOI21_X1 i_2081 (.A(n_3102), .B1(n_1517), .B2(n_1552), .ZN(n_2967));
   XNOR2_X1 i_2082 (.A(n_2976), .B(n_2975), .ZN(p_0[45]));
   XOR2_X1 i_2083 (.A(n_2973), .B(n_2972), .Z(p_0[46]));
   XNOR2_X1 i_2084 (.A(n_2969), .B(n_2968), .ZN(p_0[47]));
   OAI22_X1 i_2085 (.A1(n_1587), .A2(n_1618), .B1(n_3066), .B2(n_2973), .ZN(
      n_2968));
   NOR2_X1 i_2086 (.A1(n_3106), .A2(n_3063), .ZN(n_2969));
   XNOR2_X1 i_2087 (.A(n_2981), .B(n_2970), .ZN(p_0[48]));
   OAI21_X1 i_2088 (.A(n_2971), .B1(n_3105), .B2(n_3063), .ZN(n_2970));
   NAND3_X1 i_2089 (.A1(n_3064), .A2(n_2972), .A3(n_2974), .ZN(n_2971));
   NOR2_X1 i_2090 (.A1(n_3107), .A2(n_3066), .ZN(n_2972));
   INV_X1 i_2091 (.A(n_2974), .ZN(n_2973));
   OAI22_X1 i_2092 (.A1(n_1553), .A2(n_1586), .B1(n_3067), .B2(n_2976), .ZN(
      n_2974));
   OAI21_X1 i_2093 (.A(n_3068), .B1(n_1553), .B2(n_1586), .ZN(n_2975));
   OAI21_X1 i_2094 (.A(n_3055), .B1(n_3094), .B2(n_2977), .ZN(n_2976));
   INV_X1 i_2095 (.A(n_2978), .ZN(n_2977));
   OAI21_X1 i_2096 (.A(n_3069), .B1(n_3109), .B2(n_2979), .ZN(n_2978));
   INV_X1 i_2097 (.A(n_2980), .ZN(n_2979));
   OAI21_X1 i_2098 (.A(n_3076), .B1(n_3118), .B2(n_3083), .ZN(n_2980));
   AOI21_X1 i_2099 (.A(n_3108), .B1(n_1649), .B2(n_1676), .ZN(n_2981));
   XOR2_X1 i_2100 (.A(n_3053), .B(n_2988), .Z(p_0[49]));
   XOR2_X1 i_2101 (.A(n_2987), .B(n_2984), .Z(p_0[50]));
   XOR2_X1 i_2102 (.A(n_2985), .B(n_2982), .Z(p_0[51]));
   NOR2_X1 i_2103 (.A1(n_3050), .A2(n_3041), .ZN(n_2982));
   XNOR2_X1 i_2104 (.A(n_2989), .B(n_2983), .ZN(p_0[52]));
   OAI22_X1 i_2105 (.A1(n_1727), .A2(n_1748), .B1(n_3041), .B2(n_2985), .ZN(
      n_2983));
   AOI21_X1 i_2106 (.A(n_3051), .B1(n_1703), .B2(n_1726), .ZN(n_2984));
   AOI21_X1 i_2107 (.A(n_3051), .B1(n_3045), .B2(n_2986), .ZN(n_2985));
   INV_X1 i_2108 (.A(n_2987), .ZN(n_2986));
   AOI21_X1 i_2109 (.A(n_3048), .B1(n_3053), .B2(n_3046), .ZN(n_2987));
   OAI21_X1 i_2110 (.A(n_3046), .B1(n_1677), .B2(n_1702), .ZN(n_2988));
   NOR2_X1 i_2111 (.A1(n_3052), .A2(n_3043), .ZN(n_2989));
   XOR2_X1 i_2112 (.A(n_3039), .B(n_2996), .Z(p_0[53]));
   XOR2_X1 i_2113 (.A(n_2995), .B(n_2992), .Z(p_0[54]));
   XOR2_X1 i_2114 (.A(n_2993), .B(n_2990), .Z(p_0[55]));
   NOR2_X1 i_2115 (.A1(n_3036), .A2(n_3027), .ZN(n_2990));
   XNOR2_X1 i_2116 (.A(n_2997), .B(n_2991), .ZN(p_0[56]));
   OAI22_X1 i_2117 (.A1(n_1803), .A2(n_1816), .B1(n_3027), .B2(n_2993), .ZN(
      n_2991));
   AOI21_X1 i_2118 (.A(n_3037), .B1(n_1787), .B2(n_1802), .ZN(n_2992));
   AOI21_X1 i_2119 (.A(n_3037), .B1(n_3031), .B2(n_2994), .ZN(n_2993));
   INV_X1 i_2120 (.A(n_2995), .ZN(n_2994));
   AOI21_X1 i_2121 (.A(n_3034), .B1(n_3039), .B2(n_3032), .ZN(n_2995));
   OAI21_X1 i_2122 (.A(n_3032), .B1(n_1769), .B2(n_1786), .ZN(n_2996));
   NOR2_X1 i_2123 (.A1(n_3038), .A2(n_3029), .ZN(n_2997));
   XOR2_X1 i_2124 (.A(n_3025), .B(n_3004), .Z(p_0[57]));
   XOR2_X1 i_2125 (.A(n_3003), .B(n_3002), .Z(p_0[58]));
   XNOR2_X1 i_2126 (.A(n_2999), .B(n_2998), .ZN(p_0[59]));
   OAI22_X1 i_2127 (.A1(n_1839), .A2(n_1846), .B1(n_3015), .B2(n_3003), .ZN(
      n_2998));
   NOR2_X1 i_2128 (.A1(n_3022), .A2(n_3011), .ZN(n_2999));
   XNOR2_X1 i_2129 (.A(n_3005), .B(n_3000), .ZN(p_0[60]));
   OAI22_X1 i_2130 (.A1(n_3003), .A2(n_3001), .B1(n_3021), .B2(n_3011), .ZN(
      n_3000));
   NAND2_X1 i_2131 (.A1(n_3012), .A2(n_3002), .ZN(n_3001));
   NOR2_X1 i_2132 (.A1(n_3023), .A2(n_3015), .ZN(n_3002));
   AOI21_X1 i_2133 (.A(n_3019), .B1(n_3025), .B2(n_3017), .ZN(n_3003));
   OAI21_X1 i_2134 (.A(n_3017), .B1(n_1829), .B2(n_1838), .ZN(n_3004));
   NOR2_X1 i_2135 (.A1(n_3024), .A2(n_3013), .ZN(n_3005));
   XOR2_X1 i_2136 (.A(n_3009), .B(n_3006), .Z(p_0[61]));
   AOI21_X1 i_2137 (.A(n_3238), .B1(n_3243), .B2(n_3242), .ZN(n_3006));
   XNOR2_X1 i_2138 (.A(n_3008), .B(n_3007), .ZN(p_0[62]));
   AOI21_X1 i_2139 (.A(n_3240), .B1(n_1859), .B2(n_3241), .ZN(n_3007));
   AOI21_X1 i_2140 (.A(n_3240), .B1(n_3239), .B2(n_3008), .ZN(p_0[63]));
   OAI22_X1 i_2141 (.A1(n_1857), .A2(n_1858), .B1(n_3238), .B2(n_3009), .ZN(
      n_3008));
   OR4_X1 i_2142 (.A1(n_3013), .A2(n_3010), .A3(n_3014), .A4(n_3018), .ZN(n_3009));
   NOR2_X1 i_2143 (.A1(n_3024), .A2(n_3012), .ZN(n_3010));
   INV_X1 i_2144 (.A(n_3012), .ZN(n_3011));
   NAND2_X1 i_2145 (.A1(n_1847), .A2(n_1852), .ZN(n_3012));
   AND2_X1 i_2146 (.A1(n_1853), .A2(n_1856), .ZN(n_3013));
   AOI21_X1 i_2147 (.A(n_3020), .B1(n_3017), .B2(n_3016), .ZN(n_3014));
   INV_X1 i_2148 (.A(n_3016), .ZN(n_3015));
   NAND2_X1 i_2149 (.A1(n_1839), .A2(n_1846), .ZN(n_3016));
   NAND2_X1 i_2150 (.A1(n_1829), .A2(n_1838), .ZN(n_3017));
   NOR3_X1 i_2151 (.A1(n_3020), .A2(n_3019), .A3(n_3025), .ZN(n_3018));
   NOR2_X1 i_2152 (.A1(n_1829), .A2(n_1838), .ZN(n_3019));
   OAI21_X1 i_2153 (.A(n_3021), .B1(n_1853), .B2(n_1856), .ZN(n_3020));
   NOR2_X1 i_2154 (.A1(n_3023), .A2(n_3022), .ZN(n_3021));
   NOR2_X1 i_2155 (.A1(n_1847), .A2(n_1852), .ZN(n_3022));
   NOR2_X1 i_2156 (.A1(n_1839), .A2(n_1846), .ZN(n_3023));
   NOR2_X1 i_2157 (.A1(n_1853), .A2(n_1856), .ZN(n_3024));
   NOR4_X1 i_2158 (.A1(n_3029), .A2(n_3026), .A3(n_3030), .A4(n_3033), .ZN(
      n_3025));
   NOR2_X1 i_2159 (.A1(n_3038), .A2(n_3028), .ZN(n_3026));
   INV_X1 i_2160 (.A(n_3028), .ZN(n_3027));
   NAND2_X1 i_2161 (.A1(n_1803), .A2(n_1816), .ZN(n_3028));
   AND2_X1 i_2162 (.A1(n_1817), .A2(n_1828), .ZN(n_3029));
   AOI21_X1 i_2163 (.A(n_3035), .B1(n_3032), .B2(n_3031), .ZN(n_3030));
   NAND2_X1 i_2164 (.A1(n_1787), .A2(n_1802), .ZN(n_3031));
   NAND2_X1 i_2165 (.A1(n_1769), .A2(n_1786), .ZN(n_3032));
   NOR3_X1 i_2166 (.A1(n_3035), .A2(n_3034), .A3(n_3039), .ZN(n_3033));
   NOR2_X1 i_2167 (.A1(n_1769), .A2(n_1786), .ZN(n_3034));
   OR3_X1 i_2168 (.A1(n_3038), .A2(n_3036), .A3(n_3037), .ZN(n_3035));
   NOR2_X1 i_2169 (.A1(n_1803), .A2(n_1816), .ZN(n_3036));
   NOR2_X1 i_2170 (.A1(n_1787), .A2(n_1802), .ZN(n_3037));
   NOR2_X1 i_2171 (.A1(n_1817), .A2(n_1828), .ZN(n_3038));
   NOR4_X1 i_2172 (.A1(n_3043), .A2(n_3040), .A3(n_3044), .A4(n_3047), .ZN(
      n_3039));
   NOR2_X1 i_2173 (.A1(n_3052), .A2(n_3042), .ZN(n_3040));
   INV_X1 i_2174 (.A(n_3042), .ZN(n_3041));
   NAND2_X1 i_2175 (.A1(n_1727), .A2(n_1748), .ZN(n_3042));
   AND2_X1 i_2176 (.A1(n_1749), .A2(n_1768), .ZN(n_3043));
   AOI21_X1 i_2177 (.A(n_3049), .B1(n_3046), .B2(n_3045), .ZN(n_3044));
   NAND2_X1 i_2178 (.A1(n_1703), .A2(n_1726), .ZN(n_3045));
   NAND2_X1 i_2179 (.A1(n_1677), .A2(n_1702), .ZN(n_3046));
   NOR3_X1 i_2180 (.A1(n_3049), .A2(n_3048), .A3(n_3053), .ZN(n_3047));
   NOR2_X1 i_2181 (.A1(n_1677), .A2(n_1702), .ZN(n_3048));
   OR3_X1 i_2182 (.A1(n_3052), .A2(n_3050), .A3(n_3051), .ZN(n_3049));
   NOR2_X1 i_2183 (.A1(n_1727), .A2(n_1748), .ZN(n_3050));
   NOR2_X1 i_2184 (.A1(n_1703), .A2(n_1726), .ZN(n_3051));
   NOR2_X1 i_2185 (.A1(n_1749), .A2(n_1768), .ZN(n_3052));
   NOR3_X1 i_2186 (.A1(n_3075), .A2(n_3054), .A3(n_3082), .ZN(n_3053));
   OAI221_X1 i_2187 (.A(n_3061), .B1(n_3103), .B2(n_3055), .C1(n_3093), .C2(
      n_3069), .ZN(n_3054));
   AOI221_X1 i_2188 (.A(n_3057), .B1(n_1517), .B2(n_1552), .C1(n_3101), .C2(
      n_3056), .ZN(n_3055));
   AND2_X1 i_2189 (.A1(n_1479), .A2(n_1516), .ZN(n_3056));
   AOI21_X1 i_2190 (.A(n_3096), .B1(n_3060), .B2(n_3059), .ZN(n_3057));
   INV_X1 i_2191 (.A(n_3059), .ZN(n_3058));
   NAND2_X1 i_2192 (.A1(n_1439), .A2(n_1478), .ZN(n_3059));
   NAND2_X1 i_2193 (.A1(n_1397), .A2(n_1438), .ZN(n_3060));
   AOI21_X1 i_2194 (.A(n_3062), .B1(n_1649), .B2(n_1676), .ZN(n_3061));
   OAI21_X1 i_2195 (.A(n_3065), .B1(n_3108), .B2(n_3064), .ZN(n_3062));
   INV_X1 i_2196 (.A(n_3064), .ZN(n_3063));
   NAND2_X1 i_2197 (.A1(n_1619), .A2(n_1648), .ZN(n_3064));
   OAI21_X1 i_2198 (.A(n_3104), .B1(n_3067), .B2(n_3066), .ZN(n_3065));
   AND2_X1 i_2199 (.A1(n_1587), .A2(n_1618), .ZN(n_3066));
   INV_X1 i_2200 (.A(n_3068), .ZN(n_3067));
   NAND2_X1 i_2201 (.A1(n_1553), .A2(n_1586), .ZN(n_3068));
   AOI221_X1 i_2202 (.A(n_3071), .B1(n_1353), .B2(n_1396), .C1(n_3115), .C2(
      n_3070), .ZN(n_3069));
   AND2_X1 i_2203 (.A1(n_1307), .A2(n_1352), .ZN(n_3070));
   AOI21_X1 i_2204 (.A(n_3110), .B1(n_3074), .B2(n_3073), .ZN(n_3071));
   INV_X1 i_2205 (.A(n_3073), .ZN(n_3072));
   NAND2_X1 i_2206 (.A1(n_1259), .A2(n_1306), .ZN(n_3073));
   NAND2_X1 i_2207 (.A1(n_1209), .A2(n_1258), .ZN(n_3074));
   NOR2_X1 i_2208 (.A1(n_3092), .A2(n_3076), .ZN(n_3075));
   AOI221_X1 i_2209 (.A(n_3078), .B1(n_1157), .B2(n_1208), .C1(n_3090), .C2(
      n_3077), .ZN(n_3076));
   AND2_X1 i_2210 (.A1(n_1103), .A2(n_1156), .ZN(n_3077));
   AOI21_X1 i_2211 (.A(n_3085), .B1(n_3081), .B2(n_3080), .ZN(n_3078));
   INV_X1 i_2212 (.A(n_3080), .ZN(n_3079));
   NAND2_X1 i_2213 (.A1(n_1047), .A2(n_1102), .ZN(n_3080));
   NAND2_X1 i_2214 (.A1(n_989), .A2(n_1046), .ZN(n_3081));
   NOR3_X1 i_2215 (.A1(n_3092), .A2(n_3083), .A3(n_3118), .ZN(n_3082));
   OR2_X1 i_2216 (.A1(n_3085), .A2(n_3084), .ZN(n_3083));
   NOR2_X1 i_2217 (.A1(n_989), .A2(n_1046), .ZN(n_3084));
   NAND3_X1 i_2218 (.A1(n_3090), .A2(n_3086), .A3(n_3088), .ZN(n_3085));
   INV_X1 i_2219 (.A(n_3087), .ZN(n_3086));
   NOR2_X1 i_2220 (.A1(n_1103), .A2(n_1156), .ZN(n_3087));
   INV_X1 i_2221 (.A(n_3089), .ZN(n_3088));
   NOR2_X1 i_2222 (.A1(n_1047), .A2(n_1102), .ZN(n_3089));
   INV_X1 i_2223 (.A(n_3091), .ZN(n_3090));
   NOR2_X1 i_2224 (.A1(n_1157), .A2(n_1208), .ZN(n_3091));
   OR2_X1 i_2225 (.A1(n_3109), .A2(n_3093), .ZN(n_3092));
   OR2_X1 i_2226 (.A1(n_3103), .A2(n_3094), .ZN(n_3093));
   OR2_X1 i_2227 (.A1(n_3096), .A2(n_3095), .ZN(n_3094));
   NOR2_X1 i_2228 (.A1(n_1397), .A2(n_1438), .ZN(n_3095));
   NAND3_X1 i_2229 (.A1(n_3101), .A2(n_3097), .A3(n_3099), .ZN(n_3096));
   INV_X1 i_2230 (.A(n_3098), .ZN(n_3097));
   NOR2_X1 i_2231 (.A1(n_1479), .A2(n_1516), .ZN(n_3098));
   INV_X1 i_2232 (.A(n_3100), .ZN(n_3099));
   NOR2_X1 i_2233 (.A1(n_1439), .A2(n_1478), .ZN(n_3100));
   INV_X1 i_2234 (.A(n_3102), .ZN(n_3101));
   NOR2_X1 i_2235 (.A1(n_1517), .A2(n_1552), .ZN(n_3102));
   OAI21_X1 i_2236 (.A(n_3104), .B1(n_1553), .B2(n_1586), .ZN(n_3103));
   NOR3_X1 i_2237 (.A1(n_3108), .A2(n_3106), .A3(n_3107), .ZN(n_3104));
   NOR2_X1 i_2238 (.A1(n_3107), .A2(n_3106), .ZN(n_3105));
   NOR2_X1 i_2239 (.A1(n_1619), .A2(n_1648), .ZN(n_3106));
   NOR2_X1 i_2240 (.A1(n_1587), .A2(n_1618), .ZN(n_3107));
   NOR2_X1 i_2241 (.A1(n_1649), .A2(n_1676), .ZN(n_3108));
   OR2_X1 i_2242 (.A1(n_3117), .A2(n_3110), .ZN(n_3109));
   NAND3_X1 i_2243 (.A1(n_3115), .A2(n_3111), .A3(n_3113), .ZN(n_3110));
   INV_X1 i_2244 (.A(n_3112), .ZN(n_3111));
   NOR2_X1 i_2245 (.A1(n_1307), .A2(n_1352), .ZN(n_3112));
   INV_X1 i_2246 (.A(n_3114), .ZN(n_3113));
   NOR2_X1 i_2247 (.A1(n_1259), .A2(n_1306), .ZN(n_3114));
   INV_X1 i_2248 (.A(n_3116), .ZN(n_3115));
   NOR2_X1 i_2249 (.A1(n_1353), .A2(n_1396), .ZN(n_3116));
   NOR2_X1 i_2250 (.A1(n_1209), .A2(n_1258), .ZN(n_3117));
   NOR3_X1 i_2251 (.A1(n_3126), .A2(n_3119), .A3(n_3144), .ZN(n_3118));
   OAI222_X1 i_2252 (.A1(n_3154), .A2(n_3138), .B1(n_3155), .B2(n_3120), 
      .C1(n_3165), .C2(n_3132), .ZN(n_3119));
   AOI221_X1 i_2253 (.A(n_3122), .B1(n_505), .B2(n_550), .C1(n_3180), .C2(n_3121), 
      .ZN(n_3120));
   AND2_X1 i_2254 (.A1(n_461), .A2(n_504), .ZN(n_3121));
   AOI21_X1 i_2255 (.A(n_3175), .B1(n_3125), .B2(n_3124), .ZN(n_3122));
   INV_X1 i_2256 (.A(n_3124), .ZN(n_3123));
   NAND2_X1 i_2257 (.A1(n_419), .A2(n_460), .ZN(n_3124));
   NAND2_X1 i_2258 (.A1(n_379), .A2(n_418), .ZN(n_3125));
   OAI222_X1 i_2259 (.A1(n_3167), .A2(n_3129), .B1(n_3173), .B2(n_3128), 
      .C1(n_3245), .C2(n_3244), .ZN(n_3126));
   INV_X1 i_2260 (.A(n_3128), .ZN(n_3127));
   NAND2_X1 i_2261 (.A1(n_869), .A2(n_928), .ZN(n_3128));
   AOI21_X1 i_2262 (.A(n_3130), .B1(n_755), .B2(n_810), .ZN(n_3129));
   AND2_X1 i_2263 (.A1(n_811), .A2(n_868), .ZN(n_3130));
   NAND2_X1 i_2264 (.A1(n_755), .A2(n_810), .ZN(n_3131));
   AOI221_X1 i_2265 (.A(n_3134), .B1(n_701), .B2(n_754), .C1(n_3163), .C2(n_3133), 
      .ZN(n_3132));
   AND2_X1 i_2266 (.A1(n_649), .A2(n_700), .ZN(n_3133));
   AOI21_X1 i_2267 (.A(n_3158), .B1(n_3137), .B2(n_3136), .ZN(n_3134));
   INV_X1 i_2268 (.A(n_3136), .ZN(n_3135));
   NAND2_X1 i_2269 (.A1(n_599), .A2(n_648), .ZN(n_3136));
   NAND2_X1 i_2270 (.A1(n_596), .A2(n_598), .ZN(n_3137));
   AOI221_X1 i_2271 (.A(n_3140), .B1(n_376), .B2(n_378), .C1(n_3152), .C2(n_3139), 
      .ZN(n_3138));
   AND2_X1 i_2272 (.A1(n_305), .A2(n_340), .ZN(n_3139));
   AOI21_X1 i_2273 (.A(n_3147), .B1(n_3143), .B2(n_3142), .ZN(n_3140));
   INV_X1 i_2274 (.A(n_3142), .ZN(n_3141));
   NAND2_X1 i_2275 (.A1(n_271), .A2(n_304), .ZN(n_3142));
   NAND2_X1 i_2276 (.A1(n_268), .A2(n_270), .ZN(n_3143));
   NOR3_X1 i_2277 (.A1(n_3154), .A2(n_3145), .A3(n_3183), .ZN(n_3144));
   OR2_X1 i_2278 (.A1(n_3147), .A2(n_3146), .ZN(n_3145));
   NOR2_X1 i_2279 (.A1(n_268), .A2(n_270), .ZN(n_3146));
   NAND3_X1 i_2280 (.A1(n_3152), .A2(n_3148), .A3(n_3150), .ZN(n_3147));
   INV_X1 i_2281 (.A(n_3149), .ZN(n_3148));
   NOR2_X1 i_2282 (.A1(n_305), .A2(n_340), .ZN(n_3149));
   INV_X1 i_2283 (.A(n_3151), .ZN(n_3150));
   NOR2_X1 i_2284 (.A1(n_271), .A2(n_304), .ZN(n_3151));
   INV_X1 i_2285 (.A(n_3153), .ZN(n_3152));
   NOR2_X1 i_2286 (.A1(n_376), .A2(n_378), .ZN(n_3153));
   OR2_X1 i_2287 (.A1(n_3174), .A2(n_3155), .ZN(n_3154));
   OR2_X1 i_2288 (.A1(n_3165), .A2(n_3156), .ZN(n_3155));
   OR2_X1 i_2289 (.A1(n_3158), .A2(n_3157), .ZN(n_3156));
   NOR2_X1 i_2290 (.A1(n_596), .A2(n_598), .ZN(n_3157));
   NAND3_X1 i_2291 (.A1(n_3163), .A2(n_3159), .A3(n_3161), .ZN(n_3158));
   INV_X1 i_2292 (.A(n_3160), .ZN(n_3159));
   NOR2_X1 i_2293 (.A1(n_649), .A2(n_700), .ZN(n_3160));
   INV_X1 i_2294 (.A(n_3162), .ZN(n_3161));
   NOR2_X1 i_2295 (.A1(n_599), .A2(n_648), .ZN(n_3162));
   INV_X1 i_2296 (.A(n_3164), .ZN(n_3163));
   NOR2_X1 i_2297 (.A1(n_701), .A2(n_754), .ZN(n_3164));
   OR2_X1 i_2298 (.A1(n_3167), .A2(n_3166), .ZN(n_3165));
   NOR2_X1 i_2299 (.A1(n_755), .A2(n_810), .ZN(n_3166));
   NAND3_X1 i_2300 (.A1(n_3172), .A2(n_3168), .A3(n_3170), .ZN(n_3167));
   INV_X1 i_2301 (.A(n_3169), .ZN(n_3168));
   NOR2_X1 i_2302 (.A1(n_869), .A2(n_928), .ZN(n_3169));
   INV_X1 i_2303 (.A(n_3171), .ZN(n_3170));
   NOR2_X1 i_2304 (.A1(n_811), .A2(n_868), .ZN(n_3171));
   INV_X1 i_2305 (.A(n_3173), .ZN(n_3172));
   NOR2_X1 i_2306 (.A1(n_929), .A2(n_988), .ZN(n_3173));
   OR2_X1 i_2307 (.A1(n_3182), .A2(n_3175), .ZN(n_3174));
   NAND3_X1 i_2308 (.A1(n_3180), .A2(n_3176), .A3(n_3178), .ZN(n_3175));
   INV_X1 i_2309 (.A(n_3177), .ZN(n_3176));
   NOR2_X1 i_2310 (.A1(n_461), .A2(n_504), .ZN(n_3177));
   INV_X1 i_2311 (.A(n_3179), .ZN(n_3178));
   NOR2_X1 i_2312 (.A1(n_419), .A2(n_460), .ZN(n_3179));
   INV_X1 i_2313 (.A(n_3181), .ZN(n_3180));
   NOR2_X1 i_2314 (.A1(n_505), .A2(n_550), .ZN(n_3181));
   NOR2_X1 i_2315 (.A1(n_379), .A2(n_418), .ZN(n_3182));
   NOR4_X1 i_2316 (.A1(n_3187), .A2(n_3184), .A3(n_3188), .A4(n_3191), .ZN(
      n_3183));
   NOR2_X1 i_2317 (.A1(n_3196), .A2(n_3186), .ZN(n_3184));
   INV_X1 i_2318 (.A(n_3186), .ZN(n_3185));
   NAND2_X1 i_2319 (.A1(n_206), .A2(n_208), .ZN(n_3186));
   AND2_X1 i_2320 (.A1(n_236), .A2(n_238), .ZN(n_3187));
   AOI21_X1 i_2321 (.A(n_3193), .B1(n_3190), .B2(n_3189), .ZN(n_3188));
   NAND2_X1 i_2322 (.A1(n_178), .A2(n_180), .ZN(n_3189));
   NAND2_X1 i_2323 (.A1(n_152), .A2(n_154), .ZN(n_3190));
   NOR3_X1 i_2324 (.A1(n_3193), .A2(n_3192), .A3(n_3197), .ZN(n_3191));
   NOR2_X1 i_2325 (.A1(n_152), .A2(n_154), .ZN(n_3192));
   OR3_X1 i_2326 (.A1(n_3196), .A2(n_3194), .A3(n_3195), .ZN(n_3193));
   NOR2_X1 i_2327 (.A1(n_206), .A2(n_208), .ZN(n_3194));
   NOR2_X1 i_2328 (.A1(n_178), .A2(n_180), .ZN(n_3195));
   NOR2_X1 i_2329 (.A1(n_236), .A2(n_238), .ZN(n_3196));
   NOR4_X1 i_2330 (.A1(n_3201), .A2(n_3198), .A3(n_3202), .A4(n_3205), .ZN(
      n_3197));
   NOR2_X1 i_2331 (.A1(n_3210), .A2(n_3200), .ZN(n_3198));
   INV_X1 i_2332 (.A(n_3200), .ZN(n_3199));
   NAND2_X1 i_2333 (.A1(n_106), .A2(n_108), .ZN(n_3200));
   AND2_X1 i_2334 (.A1(n_128), .A2(n_130), .ZN(n_3201));
   AOI21_X1 i_2335 (.A(n_3207), .B1(n_3204), .B2(n_3203), .ZN(n_3202));
   NAND2_X1 i_2336 (.A1(n_86), .A2(n_88), .ZN(n_3203));
   NAND2_X1 i_2337 (.A1(n_68), .A2(n_70), .ZN(n_3204));
   NOR3_X1 i_2338 (.A1(n_3207), .A2(n_3206), .A3(n_3211), .ZN(n_3205));
   NOR2_X1 i_2339 (.A1(n_68), .A2(n_70), .ZN(n_3206));
   OR3_X1 i_2340 (.A1(n_3210), .A2(n_3208), .A3(n_3209), .ZN(n_3207));
   NOR2_X1 i_2341 (.A1(n_106), .A2(n_108), .ZN(n_3208));
   NOR2_X1 i_2342 (.A1(n_86), .A2(n_88), .ZN(n_3209));
   NOR2_X1 i_2343 (.A1(n_128), .A2(n_130), .ZN(n_3210));
   NOR4_X1 i_2344 (.A1(n_3215), .A2(n_3212), .A3(n_3216), .A4(n_3219), .ZN(
      n_3211));
   NOR2_X1 i_2345 (.A1(n_3224), .A2(n_3214), .ZN(n_3212));
   INV_X1 i_2346 (.A(n_3214), .ZN(n_3213));
   NAND2_X1 i_2347 (.A1(n_38), .A2(n_40), .ZN(n_3214));
   AND2_X1 i_2348 (.A1(n_52), .A2(n_54), .ZN(n_3215));
   AOI21_X1 i_2349 (.A(n_3221), .B1(n_3218), .B2(n_3217), .ZN(n_3216));
   NAND2_X1 i_2350 (.A1(n_26), .A2(n_28), .ZN(n_3217));
   NAND2_X1 i_2351 (.A1(n_16), .A2(n_18), .ZN(n_3218));
   NOR3_X1 i_2352 (.A1(n_3221), .A2(n_3220), .A3(n_3225), .ZN(n_3219));
   NOR2_X1 i_2353 (.A1(n_16), .A2(n_18), .ZN(n_3220));
   OR3_X1 i_2354 (.A1(n_3224), .A2(n_3222), .A3(n_3223), .ZN(n_3221));
   NOR2_X1 i_2355 (.A1(n_38), .A2(n_40), .ZN(n_3222));
   NOR2_X1 i_2356 (.A1(n_26), .A2(n_28), .ZN(n_3223));
   NOR2_X1 i_2357 (.A1(n_52), .A2(n_54), .ZN(n_3224));
   OAI22_X1 i_2358 (.A1(n_6), .A2(n_10), .B1(n_3237), .B2(n_3226), .ZN(n_3225));
   NAND2_X1 i_2359 (.A1(n_3236), .A2(n_3227), .ZN(n_3226));
   OAI21_X1 i_2360 (.A(n_3228), .B1(n_2), .B2(n_4), .ZN(n_3227));
   AOI21_X1 i_2361 (.A(n_3234), .B1(n_3230), .B2(n_3229), .ZN(n_3228));
   NAND2_X1 i_2362 (.A1(n_0), .A2(n_3235), .ZN(n_3229));
   NAND2_X1 i_2363 (.A1(p_0[0]), .A2(n_3231), .ZN(n_3230));
   NOR2_X1 i_2364 (.A1(n_3279), .A2(n_3247), .ZN(n_3231));
   NOR2_X1 i_2365 (.A1(n_3278), .A2(n_3246), .ZN(p_0[0]));
   NOR2_X1 i_2366 (.A1(n_3278), .A2(n_3247), .ZN(n_3232));
   NOR2_X1 i_2367 (.A1(n_3279), .A2(n_3246), .ZN(n_3233));
   NOR2_X1 i_2368 (.A1(n_0), .A2(n_3235), .ZN(n_3234));
   NOR2_X1 i_2369 (.A1(n_3278), .A2(n_3248), .ZN(n_3235));
   NAND2_X1 i_2370 (.A1(n_2), .A2(n_4), .ZN(n_3236));
   AND2_X1 i_2371 (.A1(n_6), .A2(n_10), .ZN(n_3237));
   NOR2_X1 i_2372 (.A1(n_3243), .A2(n_3242), .ZN(n_3238));
   NAND2_X1 i_2373 (.A1(n_1859), .A2(n_3241), .ZN(n_3239));
   NOR2_X1 i_2374 (.A1(n_1859), .A2(n_3241), .ZN(n_3240));
   NOR2_X1 i_2375 (.A1(n_3309), .A2(n_3277), .ZN(n_3241));
   INV_X1 i_2376 (.A(n_1858), .ZN(n_3242));
   INV_X1 i_2377 (.A(n_1857), .ZN(n_3243));
   INV_X1 i_2378 (.A(n_988), .ZN(n_3244));
   INV_X1 i_2379 (.A(n_929), .ZN(n_3245));
   INV_X1 i_2380 (.A(a[0]), .ZN(n_3246));
   INV_X1 i_2381 (.A(a[1]), .ZN(n_3247));
   INV_X1 i_2382 (.A(a[2]), .ZN(n_3248));
   INV_X1 i_2383 (.A(a[3]), .ZN(n_3249));
   INV_X1 i_2384 (.A(a[4]), .ZN(n_3250));
   INV_X1 i_2385 (.A(a[5]), .ZN(n_3251));
   INV_X1 i_2386 (.A(a[6]), .ZN(n_3252));
   INV_X1 i_2387 (.A(a[7]), .ZN(n_3253));
   INV_X1 i_2388 (.A(a[8]), .ZN(n_3254));
   INV_X1 i_2389 (.A(a[9]), .ZN(n_3255));
   INV_X1 i_2390 (.A(a[10]), .ZN(n_3256));
   INV_X1 i_2391 (.A(a[11]), .ZN(n_3257));
   INV_X1 i_2392 (.A(a[12]), .ZN(n_3258));
   INV_X1 i_2393 (.A(a[13]), .ZN(n_3259));
   INV_X1 i_2394 (.A(a[14]), .ZN(n_3260));
   INV_X1 i_2395 (.A(a[15]), .ZN(n_3261));
   INV_X1 i_2396 (.A(a[16]), .ZN(n_3262));
   INV_X1 i_2397 (.A(a[17]), .ZN(n_3263));
   INV_X1 i_2398 (.A(a[18]), .ZN(n_3264));
   INV_X1 i_2399 (.A(a[19]), .ZN(n_3265));
   INV_X1 i_2400 (.A(a[20]), .ZN(n_3266));
   INV_X1 i_2401 (.A(a[21]), .ZN(n_3267));
   INV_X1 i_2402 (.A(a[22]), .ZN(n_3268));
   INV_X1 i_2403 (.A(a[23]), .ZN(n_3269));
   INV_X1 i_2404 (.A(a[24]), .ZN(n_3270));
   INV_X1 i_2405 (.A(a[25]), .ZN(n_3271));
   INV_X1 i_2406 (.A(a[26]), .ZN(n_3272));
   INV_X1 i_2407 (.A(a[27]), .ZN(n_3273));
   INV_X1 i_2408 (.A(a[28]), .ZN(n_3274));
   INV_X1 i_2409 (.A(a[29]), .ZN(n_3275));
   INV_X1 i_2410 (.A(a[30]), .ZN(n_3276));
   INV_X1 i_2411 (.A(a[31]), .ZN(n_3277));
   INV_X1 i_2412 (.A(b[0]), .ZN(n_3278));
   INV_X1 i_2413 (.A(b[1]), .ZN(n_3279));
   INV_X1 i_2414 (.A(b[2]), .ZN(n_3280));
   INV_X1 i_2415 (.A(b[3]), .ZN(n_3281));
   INV_X1 i_2416 (.A(b[4]), .ZN(n_3282));
   INV_X1 i_2417 (.A(b[5]), .ZN(n_3283));
   INV_X1 i_2418 (.A(b[6]), .ZN(n_3284));
   INV_X1 i_2419 (.A(b[7]), .ZN(n_3285));
   INV_X1 i_2420 (.A(b[8]), .ZN(n_3286));
   INV_X1 i_2421 (.A(b[9]), .ZN(n_3287));
   INV_X1 i_2422 (.A(b[10]), .ZN(n_3288));
   INV_X1 i_2423 (.A(b[11]), .ZN(n_3289));
   INV_X1 i_2424 (.A(b[12]), .ZN(n_3290));
   INV_X1 i_2425 (.A(b[13]), .ZN(n_3291));
   INV_X1 i_2426 (.A(b[14]), .ZN(n_3292));
   INV_X1 i_2427 (.A(b[15]), .ZN(n_3293));
   INV_X1 i_2428 (.A(b[16]), .ZN(n_3294));
   INV_X1 i_2429 (.A(b[17]), .ZN(n_3295));
   INV_X1 i_2430 (.A(b[18]), .ZN(n_3296));
   INV_X1 i_2431 (.A(b[19]), .ZN(n_3297));
   INV_X1 i_2432 (.A(b[20]), .ZN(n_3298));
   INV_X1 i_2433 (.A(b[21]), .ZN(n_3299));
   INV_X1 i_2434 (.A(b[22]), .ZN(n_3300));
   INV_X1 i_2435 (.A(b[23]), .ZN(n_3301));
   INV_X1 i_2436 (.A(b[24]), .ZN(n_3302));
   INV_X1 i_2437 (.A(b[25]), .ZN(n_3303));
   INV_X1 i_2438 (.A(b[26]), .ZN(n_3304));
   INV_X1 i_2439 (.A(b[27]), .ZN(n_3305));
   INV_X1 i_2440 (.A(b[28]), .ZN(n_3306));
   INV_X1 i_2441 (.A(b[29]), .ZN(n_3307));
   INV_X1 i_2442 (.A(b[30]), .ZN(n_3308));
   INV_X1 i_2443 (.A(b[31]), .ZN(n_3309));
endmodule

module multOperator(clk, rst, a, b, c);
   input clk;
   input rst;
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   DFFR_X1 \c_reg[63]  (.D(n_64), .RN(n_0), .CK(clk), .Q(c[63]), .QN());
   INV_X1 i_0_0 (.A(rst), .ZN(n_0));
   DFFR_X1 \c_reg[62]  (.D(n_63), .RN(n_0), .CK(clk), .Q(c[62]), .QN());
   DFFR_X1 \c_reg[61]  (.D(n_62), .RN(n_0), .CK(clk), .Q(c[61]), .QN());
   DFFR_X1 \c_reg[60]  (.D(n_61), .RN(n_0), .CK(clk), .Q(c[60]), .QN());
   DFFR_X1 \c_reg[59]  (.D(n_60), .RN(n_0), .CK(clk), .Q(c[59]), .QN());
   DFFR_X1 \c_reg[58]  (.D(n_59), .RN(n_0), .CK(clk), .Q(c[58]), .QN());
   DFFR_X1 \c_reg[57]  (.D(n_58), .RN(n_0), .CK(clk), .Q(c[57]), .QN());
   DFFR_X1 \c_reg[56]  (.D(n_57), .RN(n_0), .CK(clk), .Q(c[56]), .QN());
   DFFR_X1 \c_reg[55]  (.D(n_56), .RN(n_0), .CK(clk), .Q(c[55]), .QN());
   DFFR_X1 \c_reg[54]  (.D(n_55), .RN(n_0), .CK(clk), .Q(c[54]), .QN());
   DFFR_X1 \c_reg[53]  (.D(n_54), .RN(n_0), .CK(clk), .Q(c[53]), .QN());
   DFFR_X1 \c_reg[52]  (.D(n_53), .RN(n_0), .CK(clk), .Q(c[52]), .QN());
   DFFR_X1 \c_reg[51]  (.D(n_52), .RN(n_0), .CK(clk), .Q(c[51]), .QN());
   DFFR_X1 \c_reg[50]  (.D(n_51), .RN(n_0), .CK(clk), .Q(c[50]), .QN());
   DFFR_X1 \c_reg[49]  (.D(n_50), .RN(n_0), .CK(clk), .Q(c[49]), .QN());
   DFFR_X1 \c_reg[48]  (.D(n_49), .RN(n_0), .CK(clk), .Q(c[48]), .QN());
   DFFR_X1 \c_reg[47]  (.D(n_48), .RN(n_0), .CK(clk), .Q(c[47]), .QN());
   DFFR_X1 \c_reg[46]  (.D(n_47), .RN(n_0), .CK(clk), .Q(c[46]), .QN());
   DFFR_X1 \c_reg[45]  (.D(n_46), .RN(n_0), .CK(clk), .Q(c[45]), .QN());
   DFFR_X1 \c_reg[44]  (.D(n_45), .RN(n_0), .CK(clk), .Q(c[44]), .QN());
   DFFR_X1 \c_reg[43]  (.D(n_44), .RN(n_0), .CK(clk), .Q(c[43]), .QN());
   DFFR_X1 \c_reg[42]  (.D(n_43), .RN(n_0), .CK(clk), .Q(c[42]), .QN());
   DFFR_X1 \c_reg[41]  (.D(n_42), .RN(n_0), .CK(clk), .Q(c[41]), .QN());
   DFFR_X1 \c_reg[40]  (.D(n_41), .RN(n_0), .CK(clk), .Q(c[40]), .QN());
   DFFR_X1 \c_reg[39]  (.D(n_40), .RN(n_0), .CK(clk), .Q(c[39]), .QN());
   DFFR_X1 \c_reg[38]  (.D(n_39), .RN(n_0), .CK(clk), .Q(c[38]), .QN());
   DFFR_X1 \c_reg[37]  (.D(n_38), .RN(n_0), .CK(clk), .Q(c[37]), .QN());
   DFFR_X1 \c_reg[36]  (.D(n_37), .RN(n_0), .CK(clk), .Q(c[36]), .QN());
   DFFR_X1 \c_reg[35]  (.D(n_36), .RN(n_0), .CK(clk), .Q(c[35]), .QN());
   DFFR_X1 \c_reg[34]  (.D(n_35), .RN(n_0), .CK(clk), .Q(c[34]), .QN());
   DFFR_X1 \c_reg[33]  (.D(n_34), .RN(n_0), .CK(clk), .Q(c[33]), .QN());
   DFFR_X1 \c_reg[32]  (.D(n_33), .RN(n_0), .CK(clk), .Q(c[32]), .QN());
   DFFR_X1 \c_reg[31]  (.D(n_32), .RN(n_0), .CK(clk), .Q(c[31]), .QN());
   DFFR_X1 \c_reg[30]  (.D(n_31), .RN(n_0), .CK(clk), .Q(c[30]), .QN());
   DFFR_X1 \c_reg[29]  (.D(n_30), .RN(n_0), .CK(clk), .Q(c[29]), .QN());
   DFFR_X1 \c_reg[28]  (.D(n_29), .RN(n_0), .CK(clk), .Q(c[28]), .QN());
   DFFR_X1 \c_reg[27]  (.D(n_28), .RN(n_0), .CK(clk), .Q(c[27]), .QN());
   DFFR_X1 \c_reg[26]  (.D(n_27), .RN(n_0), .CK(clk), .Q(c[26]), .QN());
   DFFR_X1 \c_reg[25]  (.D(n_26), .RN(n_0), .CK(clk), .Q(c[25]), .QN());
   DFFR_X1 \c_reg[24]  (.D(n_25), .RN(n_0), .CK(clk), .Q(c[24]), .QN());
   DFFR_X1 \c_reg[23]  (.D(n_24), .RN(n_0), .CK(clk), .Q(c[23]), .QN());
   DFFR_X1 \c_reg[22]  (.D(n_23), .RN(n_0), .CK(clk), .Q(c[22]), .QN());
   DFFR_X1 \c_reg[21]  (.D(n_22), .RN(n_0), .CK(clk), .Q(c[21]), .QN());
   DFFR_X1 \c_reg[20]  (.D(n_21), .RN(n_0), .CK(clk), .Q(c[20]), .QN());
   DFFR_X1 \c_reg[19]  (.D(n_20), .RN(n_0), .CK(clk), .Q(c[19]), .QN());
   DFFR_X1 \c_reg[18]  (.D(n_19), .RN(n_0), .CK(clk), .Q(c[18]), .QN());
   DFFR_X1 \c_reg[17]  (.D(n_18), .RN(n_0), .CK(clk), .Q(c[17]), .QN());
   DFFR_X1 \c_reg[16]  (.D(n_17), .RN(n_0), .CK(clk), .Q(c[16]), .QN());
   DFFR_X1 \c_reg[15]  (.D(n_16), .RN(n_0), .CK(clk), .Q(c[15]), .QN());
   DFFR_X1 \c_reg[14]  (.D(n_15), .RN(n_0), .CK(clk), .Q(c[14]), .QN());
   DFFR_X1 \c_reg[13]  (.D(n_14), .RN(n_0), .CK(clk), .Q(c[13]), .QN());
   DFFR_X1 \c_reg[12]  (.D(n_13), .RN(n_0), .CK(clk), .Q(c[12]), .QN());
   DFFR_X1 \c_reg[11]  (.D(n_12), .RN(n_0), .CK(clk), .Q(c[11]), .QN());
   DFFR_X1 \c_reg[10]  (.D(n_11), .RN(n_0), .CK(clk), .Q(c[10]), .QN());
   DFFR_X1 \c_reg[9]  (.D(n_10), .RN(n_0), .CK(clk), .Q(c[9]), .QN());
   DFFR_X1 \c_reg[8]  (.D(n_9), .RN(n_0), .CK(clk), .Q(c[8]), .QN());
   DFFR_X1 \c_reg[7]  (.D(n_8), .RN(n_0), .CK(clk), .Q(c[7]), .QN());
   DFFR_X1 \c_reg[6]  (.D(n_7), .RN(n_0), .CK(clk), .Q(c[6]), .QN());
   DFFR_X1 \c_reg[5]  (.D(n_6), .RN(n_0), .CK(clk), .Q(c[5]), .QN());
   DFFR_X1 \c_reg[4]  (.D(n_5), .RN(n_0), .CK(clk), .Q(c[4]), .QN());
   DFFR_X1 \c_reg[3]  (.D(n_4), .RN(n_0), .CK(clk), .Q(c[3]), .QN());
   DFFR_X1 \c_reg[2]  (.D(n_3), .RN(n_0), .CK(clk), .Q(c[2]), .QN());
   DFFR_X1 \c_reg[1]  (.D(n_2), .RN(n_0), .CK(clk), .Q(c[1]), .QN());
   DFFR_X1 \c_reg[0]  (.D(n_1), .RN(n_0), .CK(clk), .Q(c[0]), .QN());
   datapath i_1 (.b(b), .a(a), .p_0({n_64, n_63, n_62, n_61, n_60, n_59, n_58, 
      n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, 
      n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, 
      n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, 
      n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, 
      n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1}));
endmodule

module buffer__parameterized0(clk, rst, en, D, Q);
   input clk;
   input rst;
   input en;
   input [63:0]D;
   output [63:0]Q;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[63]  (.D(n_65), .CK(n_0), .Q(Q[63]), .QN());
   DFF_X1 \Q_reg[62]  (.D(n_64), .CK(n_0), .Q(Q[62]), .QN());
   DFF_X1 \Q_reg[61]  (.D(n_63), .CK(n_0), .Q(Q[61]), .QN());
   DFF_X1 \Q_reg[60]  (.D(n_62), .CK(n_0), .Q(Q[60]), .QN());
   DFF_X1 \Q_reg[59]  (.D(n_61), .CK(n_0), .Q(Q[59]), .QN());
   DFF_X1 \Q_reg[58]  (.D(n_60), .CK(n_0), .Q(Q[58]), .QN());
   DFF_X1 \Q_reg[57]  (.D(n_59), .CK(n_0), .Q(Q[57]), .QN());
   DFF_X1 \Q_reg[56]  (.D(n_58), .CK(n_0), .Q(Q[56]), .QN());
   DFF_X1 \Q_reg[55]  (.D(n_57), .CK(n_0), .Q(Q[55]), .QN());
   DFF_X1 \Q_reg[54]  (.D(n_56), .CK(n_0), .Q(Q[54]), .QN());
   DFF_X1 \Q_reg[53]  (.D(n_55), .CK(n_0), .Q(Q[53]), .QN());
   DFF_X1 \Q_reg[52]  (.D(n_54), .CK(n_0), .Q(Q[52]), .QN());
   DFF_X1 \Q_reg[51]  (.D(n_53), .CK(n_0), .Q(Q[51]), .QN());
   DFF_X1 \Q_reg[50]  (.D(n_52), .CK(n_0), .Q(Q[50]), .QN());
   DFF_X1 \Q_reg[49]  (.D(n_51), .CK(n_0), .Q(Q[49]), .QN());
   DFF_X1 \Q_reg[48]  (.D(n_50), .CK(n_0), .Q(Q[48]), .QN());
   DFF_X1 \Q_reg[47]  (.D(n_49), .CK(n_0), .Q(Q[47]), .QN());
   DFF_X1 \Q_reg[46]  (.D(n_48), .CK(n_0), .Q(Q[46]), .QN());
   DFF_X1 \Q_reg[45]  (.D(n_47), .CK(n_0), .Q(Q[45]), .QN());
   DFF_X1 \Q_reg[44]  (.D(n_46), .CK(n_0), .Q(Q[44]), .QN());
   DFF_X1 \Q_reg[43]  (.D(n_45), .CK(n_0), .Q(Q[43]), .QN());
   DFF_X1 \Q_reg[42]  (.D(n_44), .CK(n_0), .Q(Q[42]), .QN());
   DFF_X1 \Q_reg[41]  (.D(n_43), .CK(n_0), .Q(Q[41]), .QN());
   DFF_X1 \Q_reg[40]  (.D(n_42), .CK(n_0), .Q(Q[40]), .QN());
   DFF_X1 \Q_reg[39]  (.D(n_41), .CK(n_0), .Q(Q[39]), .QN());
   DFF_X1 \Q_reg[38]  (.D(n_40), .CK(n_0), .Q(Q[38]), .QN());
   DFF_X1 \Q_reg[37]  (.D(n_39), .CK(n_0), .Q(Q[37]), .QN());
   DFF_X1 \Q_reg[36]  (.D(n_38), .CK(n_0), .Q(Q[36]), .QN());
   DFF_X1 \Q_reg[35]  (.D(n_37), .CK(n_0), .Q(Q[35]), .QN());
   DFF_X1 \Q_reg[34]  (.D(n_36), .CK(n_0), .Q(Q[34]), .QN());
   DFF_X1 \Q_reg[33]  (.D(n_35), .CK(n_0), .Q(Q[33]), .QN());
   DFF_X1 \Q_reg[32]  (.D(n_34), .CK(n_0), .Q(Q[32]), .QN());
   DFF_X1 \Q_reg[31]  (.D(n_33), .CK(n_0), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_32), .CK(n_0), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_31), .CK(n_0), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_30), .CK(n_0), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_29), .CK(n_0), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_28), .CK(n_0), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_27), .CK(n_0), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_26), .CK(n_0), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_25), .CK(n_0), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_24), .CK(n_0), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_23), .CK(n_0), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_22), .CK(n_0), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_21), .CK(n_0), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_20), .CK(n_0), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_19), .CK(n_0), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_18), .CK(n_0), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_17), .CK(n_0), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_16), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_15), .CK(n_0), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_14), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_13), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_12), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_11), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_10), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_9), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_8), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_7), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_6), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_5), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_4), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_3), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_2), .CK(n_0), .Q(Q[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(rst), .ZN(n_1));
   INV_X1 i_0_1 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(D[31]), .ZN(n_33));
   AND2_X1 i_0_34 (.A1(n_0_0), .A2(D[32]), .ZN(n_34));
   AND2_X1 i_0_35 (.A1(n_0_0), .A2(D[33]), .ZN(n_35));
   AND2_X1 i_0_36 (.A1(n_0_0), .A2(D[34]), .ZN(n_36));
   AND2_X1 i_0_37 (.A1(n_0_0), .A2(D[35]), .ZN(n_37));
   AND2_X1 i_0_38 (.A1(n_0_0), .A2(D[36]), .ZN(n_38));
   AND2_X1 i_0_39 (.A1(n_0_0), .A2(D[37]), .ZN(n_39));
   AND2_X1 i_0_40 (.A1(n_0_0), .A2(D[38]), .ZN(n_40));
   AND2_X1 i_0_41 (.A1(n_0_0), .A2(D[39]), .ZN(n_41));
   AND2_X1 i_0_42 (.A1(n_0_0), .A2(D[40]), .ZN(n_42));
   AND2_X1 i_0_43 (.A1(n_0_0), .A2(D[41]), .ZN(n_43));
   AND2_X1 i_0_44 (.A1(n_0_0), .A2(D[42]), .ZN(n_44));
   AND2_X1 i_0_45 (.A1(n_0_0), .A2(D[43]), .ZN(n_45));
   AND2_X1 i_0_46 (.A1(n_0_0), .A2(D[44]), .ZN(n_46));
   AND2_X1 i_0_47 (.A1(n_0_0), .A2(D[45]), .ZN(n_47));
   AND2_X1 i_0_48 (.A1(n_0_0), .A2(D[46]), .ZN(n_48));
   AND2_X1 i_0_49 (.A1(n_0_0), .A2(D[47]), .ZN(n_49));
   AND2_X1 i_0_50 (.A1(n_0_0), .A2(D[48]), .ZN(n_50));
   AND2_X1 i_0_51 (.A1(n_0_0), .A2(D[49]), .ZN(n_51));
   AND2_X1 i_0_52 (.A1(n_0_0), .A2(D[50]), .ZN(n_52));
   AND2_X1 i_0_53 (.A1(n_0_0), .A2(D[51]), .ZN(n_53));
   AND2_X1 i_0_54 (.A1(n_0_0), .A2(D[52]), .ZN(n_54));
   AND2_X1 i_0_55 (.A1(n_0_0), .A2(D[53]), .ZN(n_55));
   AND2_X1 i_0_56 (.A1(n_0_0), .A2(D[54]), .ZN(n_56));
   AND2_X1 i_0_57 (.A1(n_0_0), .A2(D[55]), .ZN(n_57));
   AND2_X1 i_0_58 (.A1(n_0_0), .A2(D[56]), .ZN(n_58));
   AND2_X1 i_0_59 (.A1(n_0_0), .A2(D[57]), .ZN(n_59));
   AND2_X1 i_0_60 (.A1(n_0_0), .A2(D[58]), .ZN(n_60));
   AND2_X1 i_0_61 (.A1(n_0_0), .A2(D[59]), .ZN(n_61));
   AND2_X1 i_0_62 (.A1(n_0_0), .A2(D[60]), .ZN(n_62));
   AND2_X1 i_0_63 (.A1(n_0_0), .A2(D[61]), .ZN(n_63));
   AND2_X1 i_0_64 (.A1(n_0_0), .A2(D[62]), .ZN(n_64));
   AND2_X1 i_0_65 (.A1(n_0_0), .A2(D[63]), .ZN(n_65));
endmodule

module simpleMultiplier(clk, rst, en, a, b, c);
   input clk;
   input rst;
   input en;
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   wire [31:0]a_out;
   wire [31:0]b_out;
   wire [63:0]c_out;

   buffer__0_68 inRegA (.clk(clk), .rst(rst), .en(en), .D(a), .Q(a_out));
   buffer inRegB (.clk(clk), .rst(rst), .en(en), .D(b), .Q(b_out));
   multOperator M64 (.clk(clk), .rst(rst), .a(a_out), .b(b_out), .c(c_out));
   buffer__parameterized0 outReg (.clk(clk), .rst(rst), .en(en), .D(c_out), 
      .Q(c));
endmodule
