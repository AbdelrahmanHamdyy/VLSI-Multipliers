/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 22:58:42 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2254582317 */

module datapath(p_0, a);
   output [31:0]p_0;
   input [31:0]a;

   XOR2_X1 i_0 (.A(a[1]), .B(a[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(a[2]), .B1(a[1]), .B2(a[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(a[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(a[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(a[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(a[6]), .B1(n_27), .B2(a[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(a[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(a[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(a[9]), .B1(n_25), .B2(a[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(a[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(a[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(a[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(a[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(a[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(a[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(a[16]), .B1(n_19), .B2(a[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(a[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(a[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(a[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(a[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(a[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(a[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(a[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(a[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(a[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(a[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(a[27]), .B1(n_9), .B2(a[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(a[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(a[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(a[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(a[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(a[28]), .A3(a[29]), .A4(a[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(a[28]), .A3(a[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(a[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(a[26]), .A3(a[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(a[23]), .A3(a[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(a[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(a[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(a[18]), .A3(a[19]), .A4(a[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(a[18]), .A3(a[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(a[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(a[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(a[15]), .A3(a[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(a[12]), .A3(a[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(a[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(a[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(a[8]), .A3(a[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(a[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(a[5]), .A3(a[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(a[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(a[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(a[2]), .A2(a[1]), .A3(a[0]), .ZN(n_29));
   INV_X1 i_61 (.A(a[11]), .ZN(n_30));
   INV_X1 i_62 (.A(a[14]), .ZN(n_31));
   INV_X1 i_63 (.A(a[21]), .ZN(n_32));
   INV_X1 i_64 (.A(a[25]), .ZN(n_33));
endmodule

module datapath__0_127(A, p_0, multiplicand);
   input [31:0]A;
   output [31:0]p_0;
   input [31:0]multiplicand;

   INV_X1 i_0 (.A(A[0]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_0), .A2(multiplicand[0]), .ZN(n_1));
   OAI21_X1 i_2 (.A(n_1), .B1(multiplicand[0]), .B2(n_0), .ZN(p_0[0]));
   XNOR2_X1 i_3 (.A(A[1]), .B(multiplicand[1]), .ZN(n_2));
   XOR2_X1 i_4 (.A(n_2), .B(n_1), .Z(p_0[1]));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   INV_X1 i_6 (.A(A[1]), .ZN(n_4));
   AOI22_X1 i_7 (.A1(n_2), .A2(n_3), .B1(n_4), .B2(multiplicand[1]), .ZN(n_5));
   XOR2_X1 i_8 (.A(multiplicand[2]), .B(A[2]), .Z(n_6));
   XNOR2_X1 i_9 (.A(n_5), .B(n_6), .ZN(p_0[2]));
   INV_X1 i_10 (.A(multiplicand[2]), .ZN(n_7));
   OAI22_X1 i_11 (.A1(n_5), .A2(n_6), .B1(n_7), .B2(A[2]), .ZN(n_8));
   XNOR2_X1 i_12 (.A(A[3]), .B(multiplicand[3]), .ZN(n_9));
   XNOR2_X1 i_13 (.A(n_8), .B(n_9), .ZN(p_0[3]));
   INV_X1 i_14 (.A(A[3]), .ZN(n_10));
   AOI22_X1 i_15 (.A1(n_8), .A2(n_9), .B1(n_10), .B2(multiplicand[3]), .ZN(n_11));
   XOR2_X1 i_16 (.A(A[4]), .B(multiplicand[4]), .Z(n_12));
   XNOR2_X1 i_17 (.A(n_11), .B(n_12), .ZN(p_0[4]));
   INV_X1 i_18 (.A(multiplicand[4]), .ZN(n_13));
   OAI22_X1 i_19 (.A1(n_11), .A2(n_12), .B1(n_13), .B2(A[4]), .ZN(n_14));
   XNOR2_X1 i_20 (.A(A[5]), .B(multiplicand[5]), .ZN(n_15));
   XNOR2_X1 i_21 (.A(n_14), .B(n_15), .ZN(p_0[5]));
   INV_X1 i_22 (.A(A[5]), .ZN(n_16));
   AOI22_X1 i_23 (.A1(n_14), .A2(n_15), .B1(n_16), .B2(multiplicand[5]), 
      .ZN(n_17));
   XOR2_X1 i_24 (.A(A[6]), .B(multiplicand[6]), .Z(n_18));
   XNOR2_X1 i_25 (.A(n_17), .B(n_18), .ZN(p_0[6]));
   INV_X1 i_26 (.A(multiplicand[6]), .ZN(n_19));
   OAI22_X1 i_27 (.A1(n_17), .A2(n_18), .B1(n_19), .B2(A[6]), .ZN(n_20));
   XNOR2_X1 i_28 (.A(A[7]), .B(multiplicand[7]), .ZN(n_21));
   XNOR2_X1 i_29 (.A(n_20), .B(n_21), .ZN(p_0[7]));
   INV_X1 i_30 (.A(A[7]), .ZN(n_22));
   AOI22_X1 i_31 (.A1(n_20), .A2(n_21), .B1(n_22), .B2(multiplicand[7]), 
      .ZN(n_23));
   XOR2_X1 i_32 (.A(A[8]), .B(multiplicand[8]), .Z(n_24));
   XNOR2_X1 i_33 (.A(n_23), .B(n_24), .ZN(p_0[8]));
   INV_X1 i_34 (.A(multiplicand[8]), .ZN(n_25));
   OAI22_X1 i_35 (.A1(n_23), .A2(n_24), .B1(n_25), .B2(A[8]), .ZN(n_26));
   XNOR2_X1 i_36 (.A(A[9]), .B(multiplicand[9]), .ZN(n_27));
   XNOR2_X1 i_37 (.A(n_26), .B(n_27), .ZN(p_0[9]));
   INV_X1 i_38 (.A(A[9]), .ZN(n_28));
   AOI22_X1 i_39 (.A1(n_26), .A2(n_27), .B1(n_28), .B2(multiplicand[9]), 
      .ZN(n_29));
   XOR2_X1 i_40 (.A(A[10]), .B(multiplicand[10]), .Z(n_30));
   XNOR2_X1 i_41 (.A(n_29), .B(n_30), .ZN(p_0[10]));
   INV_X1 i_42 (.A(multiplicand[10]), .ZN(n_31));
   OAI22_X1 i_43 (.A1(n_29), .A2(n_30), .B1(n_31), .B2(A[10]), .ZN(n_32));
   XNOR2_X1 i_44 (.A(A[11]), .B(multiplicand[11]), .ZN(n_33));
   XNOR2_X1 i_45 (.A(n_32), .B(n_33), .ZN(p_0[11]));
   INV_X1 i_46 (.A(A[11]), .ZN(n_34));
   AOI22_X1 i_47 (.A1(n_32), .A2(n_33), .B1(n_34), .B2(multiplicand[11]), 
      .ZN(n_35));
   XOR2_X1 i_48 (.A(A[12]), .B(multiplicand[12]), .Z(n_36));
   XNOR2_X1 i_49 (.A(n_35), .B(n_36), .ZN(p_0[12]));
   INV_X1 i_50 (.A(multiplicand[12]), .ZN(n_37));
   OAI22_X1 i_51 (.A1(n_35), .A2(n_36), .B1(n_37), .B2(A[12]), .ZN(n_38));
   XNOR2_X1 i_52 (.A(A[13]), .B(multiplicand[13]), .ZN(n_39));
   XNOR2_X1 i_53 (.A(n_38), .B(n_39), .ZN(p_0[13]));
   INV_X1 i_54 (.A(A[13]), .ZN(n_40));
   AOI22_X1 i_55 (.A1(n_38), .A2(n_39), .B1(n_40), .B2(multiplicand[13]), 
      .ZN(n_41));
   XOR2_X1 i_56 (.A(A[14]), .B(multiplicand[14]), .Z(n_42));
   XNOR2_X1 i_57 (.A(n_41), .B(n_42), .ZN(p_0[14]));
   INV_X1 i_58 (.A(multiplicand[14]), .ZN(n_43));
   OAI22_X1 i_59 (.A1(n_41), .A2(n_42), .B1(n_43), .B2(A[14]), .ZN(n_44));
   XNOR2_X1 i_60 (.A(A[15]), .B(multiplicand[15]), .ZN(n_45));
   XNOR2_X1 i_61 (.A(n_44), .B(n_45), .ZN(p_0[15]));
   INV_X1 i_62 (.A(A[15]), .ZN(n_46));
   AOI22_X1 i_63 (.A1(n_44), .A2(n_45), .B1(n_46), .B2(multiplicand[15]), 
      .ZN(n_47));
   XOR2_X1 i_64 (.A(A[16]), .B(multiplicand[16]), .Z(n_48));
   XNOR2_X1 i_65 (.A(n_47), .B(n_48), .ZN(p_0[16]));
   INV_X1 i_66 (.A(multiplicand[16]), .ZN(n_49));
   OAI22_X1 i_67 (.A1(n_47), .A2(n_48), .B1(n_49), .B2(A[16]), .ZN(n_50));
   XNOR2_X1 i_68 (.A(A[17]), .B(multiplicand[17]), .ZN(n_51));
   XNOR2_X1 i_69 (.A(n_50), .B(n_51), .ZN(p_0[17]));
   INV_X1 i_70 (.A(A[17]), .ZN(n_52));
   AOI22_X1 i_71 (.A1(n_50), .A2(n_51), .B1(n_52), .B2(multiplicand[17]), 
      .ZN(n_53));
   XOR2_X1 i_72 (.A(A[18]), .B(multiplicand[18]), .Z(n_54));
   XNOR2_X1 i_73 (.A(n_53), .B(n_54), .ZN(p_0[18]));
   INV_X1 i_74 (.A(multiplicand[18]), .ZN(n_55));
   OAI22_X1 i_75 (.A1(n_53), .A2(n_54), .B1(n_55), .B2(A[18]), .ZN(n_56));
   XNOR2_X1 i_76 (.A(A[19]), .B(multiplicand[19]), .ZN(n_57));
   XNOR2_X1 i_77 (.A(n_56), .B(n_57), .ZN(p_0[19]));
   INV_X1 i_78 (.A(A[19]), .ZN(n_58));
   AOI22_X1 i_79 (.A1(n_56), .A2(n_57), .B1(n_58), .B2(multiplicand[19]), 
      .ZN(n_59));
   XOR2_X1 i_80 (.A(A[20]), .B(multiplicand[20]), .Z(n_60));
   XNOR2_X1 i_81 (.A(n_59), .B(n_60), .ZN(p_0[20]));
   INV_X1 i_82 (.A(multiplicand[20]), .ZN(n_61));
   OAI22_X1 i_83 (.A1(n_59), .A2(n_60), .B1(n_61), .B2(A[20]), .ZN(n_62));
   XNOR2_X1 i_84 (.A(A[21]), .B(multiplicand[21]), .ZN(n_63));
   XNOR2_X1 i_85 (.A(n_62), .B(n_63), .ZN(p_0[21]));
   INV_X1 i_86 (.A(A[21]), .ZN(n_64));
   AOI22_X1 i_87 (.A1(n_62), .A2(n_63), .B1(n_64), .B2(multiplicand[21]), 
      .ZN(n_65));
   XOR2_X1 i_88 (.A(A[22]), .B(multiplicand[22]), .Z(n_66));
   XNOR2_X1 i_89 (.A(n_65), .B(n_66), .ZN(p_0[22]));
   INV_X1 i_90 (.A(multiplicand[22]), .ZN(n_67));
   OAI22_X1 i_91 (.A1(n_65), .A2(n_66), .B1(n_67), .B2(A[22]), .ZN(n_68));
   XNOR2_X1 i_92 (.A(A[23]), .B(multiplicand[23]), .ZN(n_69));
   XNOR2_X1 i_93 (.A(n_68), .B(n_69), .ZN(p_0[23]));
   INV_X1 i_94 (.A(A[23]), .ZN(n_70));
   AOI22_X1 i_95 (.A1(n_68), .A2(n_69), .B1(n_70), .B2(multiplicand[23]), 
      .ZN(n_71));
   XOR2_X1 i_96 (.A(A[24]), .B(multiplicand[24]), .Z(n_72));
   XNOR2_X1 i_97 (.A(n_71), .B(n_72), .ZN(p_0[24]));
   INV_X1 i_98 (.A(multiplicand[24]), .ZN(n_73));
   OAI22_X1 i_99 (.A1(n_71), .A2(n_72), .B1(n_73), .B2(A[24]), .ZN(n_74));
   XNOR2_X1 i_100 (.A(A[25]), .B(multiplicand[25]), .ZN(n_75));
   XNOR2_X1 i_101 (.A(n_74), .B(n_75), .ZN(p_0[25]));
   INV_X1 i_102 (.A(A[25]), .ZN(n_76));
   AOI22_X1 i_103 (.A1(n_74), .A2(n_75), .B1(n_76), .B2(multiplicand[25]), 
      .ZN(n_77));
   XOR2_X1 i_104 (.A(A[26]), .B(multiplicand[26]), .Z(n_78));
   XNOR2_X1 i_105 (.A(n_77), .B(n_78), .ZN(p_0[26]));
   INV_X1 i_106 (.A(multiplicand[26]), .ZN(n_79));
   OAI22_X1 i_107 (.A1(n_77), .A2(n_78), .B1(n_79), .B2(A[26]), .ZN(n_80));
   XNOR2_X1 i_108 (.A(A[27]), .B(multiplicand[27]), .ZN(n_81));
   XNOR2_X1 i_109 (.A(n_80), .B(n_81), .ZN(p_0[27]));
   INV_X1 i_110 (.A(A[27]), .ZN(n_82));
   AOI22_X1 i_111 (.A1(n_80), .A2(n_81), .B1(n_82), .B2(multiplicand[27]), 
      .ZN(n_83));
   XOR2_X1 i_112 (.A(A[28]), .B(multiplicand[28]), .Z(n_84));
   XNOR2_X1 i_113 (.A(n_83), .B(n_84), .ZN(p_0[28]));
   INV_X1 i_114 (.A(multiplicand[28]), .ZN(n_85));
   OAI22_X1 i_115 (.A1(n_83), .A2(n_84), .B1(n_85), .B2(A[28]), .ZN(n_86));
   XNOR2_X1 i_116 (.A(A[29]), .B(multiplicand[29]), .ZN(n_87));
   XNOR2_X1 i_117 (.A(n_86), .B(n_87), .ZN(p_0[29]));
   INV_X1 i_118 (.A(A[29]), .ZN(n_88));
   AOI22_X1 i_119 (.A1(n_86), .A2(n_87), .B1(n_88), .B2(multiplicand[29]), 
      .ZN(n_89));
   INV_X1 i_120 (.A(A[31]), .ZN(n_90));
   INV_X1 i_121 (.A(multiplicand[30]), .ZN(n_91));
   AOI22_X1 i_122 (.A1(n_90), .A2(n_91), .B1(A[31]), .B2(multiplicand[30]), 
      .ZN(n_92));
   XNOR2_X1 i_123 (.A(n_89), .B(n_92), .ZN(p_0[30]));
   INV_X1 i_124 (.A(n_89), .ZN(n_93));
   OAI33_X1 i_125 (.A1(n_93), .A2(A[31]), .A3(multiplicand[30]), .B1(n_89), 
      .B2(n_90), .B3(n_91), .ZN(n_94));
   XNOR2_X1 i_126 (.A(n_94), .B(multiplicand[31]), .ZN(p_0[31]));
endmodule

module datapath__0_128(multiplicand, A, p_0);
   input [31:0]multiplicand;
   input [31:0]A;
   output [31:0]p_0;

   HA_X1 i_0 (.A(multiplicand[0]), .B(A[0]), .CO(n_0), .S(p_0[0]));
   FA_X1 i_1 (.A(multiplicand[1]), .B(A[1]), .CI(n_0), .CO(n_1), .S(p_0[1]));
   FA_X1 i_2 (.A(multiplicand[2]), .B(A[2]), .CI(n_1), .CO(n_2), .S(p_0[2]));
   FA_X1 i_3 (.A(multiplicand[3]), .B(A[3]), .CI(n_2), .CO(n_3), .S(p_0[3]));
   FA_X1 i_4 (.A(multiplicand[4]), .B(A[4]), .CI(n_3), .CO(n_4), .S(p_0[4]));
   FA_X1 i_5 (.A(multiplicand[5]), .B(A[5]), .CI(n_4), .CO(n_5), .S(p_0[5]));
   FA_X1 i_6 (.A(multiplicand[6]), .B(A[6]), .CI(n_5), .CO(n_6), .S(p_0[6]));
   FA_X1 i_7 (.A(multiplicand[7]), .B(A[7]), .CI(n_6), .CO(n_7), .S(p_0[7]));
   FA_X1 i_8 (.A(multiplicand[8]), .B(A[8]), .CI(n_7), .CO(n_8), .S(p_0[8]));
   FA_X1 i_9 (.A(multiplicand[9]), .B(A[9]), .CI(n_8), .CO(n_9), .S(p_0[9]));
   FA_X1 i_10 (.A(multiplicand[10]), .B(A[10]), .CI(n_9), .CO(n_10), .S(p_0[10]));
   FA_X1 i_11 (.A(multiplicand[11]), .B(A[11]), .CI(n_10), .CO(n_11), .S(p_0[11]));
   FA_X1 i_12 (.A(multiplicand[12]), .B(A[12]), .CI(n_11), .CO(n_12), .S(p_0[12]));
   FA_X1 i_13 (.A(multiplicand[13]), .B(A[13]), .CI(n_12), .CO(n_13), .S(p_0[13]));
   FA_X1 i_14 (.A(multiplicand[14]), .B(A[14]), .CI(n_13), .CO(n_14), .S(p_0[14]));
   FA_X1 i_15 (.A(multiplicand[15]), .B(A[15]), .CI(n_14), .CO(n_15), .S(p_0[15]));
   FA_X1 i_16 (.A(multiplicand[16]), .B(A[16]), .CI(n_15), .CO(n_16), .S(p_0[16]));
   FA_X1 i_17 (.A(multiplicand[17]), .B(A[17]), .CI(n_16), .CO(n_17), .S(p_0[17]));
   FA_X1 i_18 (.A(multiplicand[18]), .B(A[18]), .CI(n_17), .CO(n_18), .S(p_0[18]));
   FA_X1 i_19 (.A(multiplicand[19]), .B(A[19]), .CI(n_18), .CO(n_19), .S(p_0[19]));
   FA_X1 i_20 (.A(multiplicand[20]), .B(A[20]), .CI(n_19), .CO(n_20), .S(p_0[20]));
   FA_X1 i_21 (.A(multiplicand[21]), .B(A[21]), .CI(n_20), .CO(n_21), .S(p_0[21]));
   FA_X1 i_22 (.A(multiplicand[22]), .B(A[22]), .CI(n_21), .CO(n_22), .S(p_0[22]));
   FA_X1 i_23 (.A(multiplicand[23]), .B(A[23]), .CI(n_22), .CO(n_23), .S(p_0[23]));
   FA_X1 i_24 (.A(multiplicand[24]), .B(A[24]), .CI(n_23), .CO(n_24), .S(p_0[24]));
   FA_X1 i_25 (.A(multiplicand[25]), .B(A[25]), .CI(n_24), .CO(n_25), .S(p_0[25]));
   FA_X1 i_26 (.A(multiplicand[26]), .B(A[26]), .CI(n_25), .CO(n_26), .S(p_0[26]));
   FA_X1 i_27 (.A(multiplicand[27]), .B(A[27]), .CI(n_26), .CO(n_27), .S(p_0[27]));
   FA_X1 i_28 (.A(multiplicand[28]), .B(A[28]), .CI(n_27), .CO(n_28), .S(p_0[28]));
   FA_X1 i_29 (.A(multiplicand[29]), .B(A[29]), .CI(n_28), .CO(n_29), .S(p_0[29]));
   FA_X1 i_30 (.A(multiplicand[30]), .B(A[31]), .CI(n_29), .CO(n_30), .S(p_0[30]));
   XNOR2_X1 i_31 (.A(multiplicand[31]), .B(A[31]), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(p_0[31]));
endmodule

module datapath__0_129(p_0, b);
   output [31:0]p_0;
   input [31:0]b;

   XOR2_X1 i_0 (.A(b[1]), .B(b[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(b[2]), .B1(b[1]), .B2(b[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(b[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(b[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(b[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(b[6]), .B1(n_27), .B2(b[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(b[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(b[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(b[9]), .B1(n_25), .B2(b[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(b[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(b[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(b[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(b[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(b[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(b[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(b[16]), .B1(n_19), .B2(b[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(b[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(b[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(b[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(b[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(b[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(b[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(b[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(b[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(b[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(b[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(b[27]), .B1(n_9), .B2(b[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(b[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(b[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(b[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(b[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(b[28]), .A3(b[29]), .A4(b[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(b[28]), .A3(b[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(b[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(b[26]), .A3(b[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(b[23]), .A3(b[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(b[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(b[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(b[18]), .A3(b[19]), .A4(b[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(b[18]), .A3(b[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(b[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(b[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(b[15]), .A3(b[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(b[12]), .A3(b[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(b[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(b[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(b[8]), .A3(b[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(b[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(b[5]), .A3(b[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(b[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(b[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(b[2]), .A2(b[1]), .A3(b[0]), .ZN(n_29));
   INV_X1 i_61 (.A(b[11]), .ZN(n_30));
   INV_X1 i_62 (.A(b[14]), .ZN(n_31));
   INV_X1 i_63 (.A(b[21]), .ZN(n_32));
   INV_X1 i_64 (.A(b[25]), .ZN(n_33));
endmodule

module datapath__0_132(p_0, p_1);
   output [63:0]p_0;
   input [63:0]p_1;

   XOR2_X1 i_0 (.A(p_1[1]), .B(p_1[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_60), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(p_1[2]), .B1(p_1[1]), .B2(p_1[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_1[3]), .B(n_60), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(p_1[4]), .B(n_59), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(p_1[5]), .B(n_58), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_57), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(p_1[6]), .B1(n_58), .B2(p_1[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_1[7]), .B(n_57), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(p_1[8]), .B(n_56), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_55), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(p_1[9]), .B1(n_56), .B2(p_1[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_1[10]), .B(n_55), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(p_1[11]), .B(n_54), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(p_1[12]), .B(n_53), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(p_1[13]), .B(n_52), .ZN(p_0[13]));
   XOR2_X1 i_16 (.A(p_1[14]), .B(n_51), .Z(p_0[14]));
   AND2_X1 i_17 (.A1(n_50), .A2(n_3), .ZN(p_0[15]));
   OAI21_X1 i_18 (.A(p_1[15]), .B1(n_51), .B2(p_1[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(p_1[16]), .B(n_50), .Z(p_0[16]));
   XOR2_X1 i_20 (.A(p_1[17]), .B(n_49), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(p_1[18]), .B(n_48), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(p_1[19]), .B(n_47), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(p_1[20]), .B(n_46), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(p_1[21]), .B(n_45), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(p_1[22]), .B(n_44), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(p_1[23]), .B(n_43), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(p_1[24]), .B(n_42), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(p_1[25]), .B(n_41), .ZN(p_0[25]));
   XNOR2_X1 i_29 (.A(p_1[26]), .B(n_40), .ZN(p_0[26]));
   XOR2_X1 i_30 (.A(p_1[27]), .B(n_39), .Z(p_0[27]));
   XOR2_X1 i_31 (.A(p_1[28]), .B(n_38), .Z(p_0[28]));
   XNOR2_X1 i_32 (.A(p_1[29]), .B(n_37), .ZN(p_0[29]));
   XNOR2_X1 i_33 (.A(p_1[30]), .B(n_36), .ZN(p_0[30]));
   XNOR2_X1 i_34 (.A(p_1[31]), .B(n_35), .ZN(p_0[31]));
   XOR2_X1 i_35 (.A(p_1[32]), .B(n_34), .Z(p_0[32]));
   XOR2_X1 i_36 (.A(p_1[33]), .B(n_33), .Z(p_0[33]));
   XNOR2_X1 i_37 (.A(p_1[34]), .B(n_32), .ZN(p_0[34]));
   XNOR2_X1 i_38 (.A(p_1[35]), .B(n_31), .ZN(p_0[35]));
   XNOR2_X1 i_39 (.A(p_1[36]), .B(n_30), .ZN(p_0[36]));
   XOR2_X1 i_40 (.A(p_1[37]), .B(n_29), .Z(p_0[37]));
   XOR2_X1 i_41 (.A(p_1[38]), .B(n_28), .Z(p_0[38]));
   XNOR2_X1 i_42 (.A(p_1[39]), .B(n_27), .ZN(p_0[39]));
   XNOR2_X1 i_43 (.A(p_1[40]), .B(n_26), .ZN(p_0[40]));
   XOR2_X1 i_44 (.A(p_1[41]), .B(n_25), .Z(p_0[41]));
   XNOR2_X1 i_45 (.A(p_1[42]), .B(n_24), .ZN(p_0[42]));
   XOR2_X1 i_46 (.A(p_1[43]), .B(n_23), .Z(p_0[43]));
   AND2_X1 i_47 (.A1(n_22), .A2(n_4), .ZN(p_0[44]));
   OAI21_X1 i_48 (.A(p_1[44]), .B1(n_23), .B2(p_1[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(p_1[45]), .B(n_22), .Z(p_0[45]));
   XOR2_X1 i_50 (.A(p_1[46]), .B(n_21), .Z(p_0[46]));
   XOR2_X1 i_51 (.A(p_1[47]), .B(n_20), .Z(p_0[47]));
   XOR2_X1 i_52 (.A(p_1[48]), .B(n_19), .Z(p_0[48]));
   XNOR2_X1 i_53 (.A(p_1[49]), .B(n_18), .ZN(p_0[49]));
   XNOR2_X1 i_54 (.A(p_1[50]), .B(n_17), .ZN(p_0[50]));
   XNOR2_X1 i_55 (.A(p_1[51]), .B(n_16), .ZN(p_0[51]));
   XOR2_X1 i_56 (.A(p_1[52]), .B(n_15), .Z(p_0[52]));
   XNOR2_X1 i_57 (.A(p_1[53]), .B(n_14), .ZN(p_0[53]));
   XNOR2_X1 i_58 (.A(p_1[54]), .B(n_13), .ZN(p_0[54]));
   XNOR2_X1 i_59 (.A(p_1[55]), .B(n_12), .ZN(p_0[55]));
   XOR2_X1 i_60 (.A(p_1[56]), .B(n_11), .Z(p_0[56]));
   AND2_X1 i_61 (.A1(n_10), .A2(n_5), .ZN(p_0[57]));
   OAI21_X1 i_62 (.A(p_1[57]), .B1(n_11), .B2(p_1[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(p_1[58]), .B(n_10), .Z(p_0[58]));
   XNOR2_X1 i_64 (.A(p_1[59]), .B(n_9), .ZN(p_0[59]));
   XNOR2_X1 i_65 (.A(p_1[60]), .B(n_8), .ZN(p_0[60]));
   XOR2_X1 i_66 (.A(p_1[61]), .B(n_7), .Z(p_0[61]));
   XNOR2_X1 i_67 (.A(p_1[62]), .B(n_6), .ZN(p_0[62]));
   NAND2_X1 i_68 (.A1(n_6), .A2(n_72), .ZN(p_0[63]));
   NOR2_X1 i_69 (.A1(n_7), .A2(p_1[61]), .ZN(n_6));
   NAND2_X1 i_70 (.A1(n_8), .A2(n_71), .ZN(n_7));
   NOR3_X1 i_71 (.A1(n_10), .A2(p_1[58]), .A3(p_1[59]), .ZN(n_8));
   NOR2_X1 i_72 (.A1(n_10), .A2(p_1[58]), .ZN(n_9));
   OR3_X1 i_73 (.A1(n_11), .A2(p_1[56]), .A3(p_1[57]), .ZN(n_10));
   NAND2_X1 i_74 (.A1(n_12), .A2(n_70), .ZN(n_11));
   NOR4_X1 i_75 (.A1(n_15), .A2(p_1[52]), .A3(p_1[53]), .A4(p_1[54]), .ZN(n_12));
   NOR3_X1 i_76 (.A1(n_15), .A2(p_1[52]), .A3(p_1[53]), .ZN(n_13));
   NOR2_X1 i_77 (.A1(n_15), .A2(p_1[52]), .ZN(n_14));
   NAND2_X1 i_78 (.A1(n_16), .A2(n_69), .ZN(n_15));
   NOR4_X1 i_79 (.A1(n_19), .A2(p_1[48]), .A3(p_1[49]), .A4(p_1[50]), .ZN(n_16));
   NOR3_X1 i_80 (.A1(n_19), .A2(p_1[48]), .A3(p_1[49]), .ZN(n_17));
   NOR2_X1 i_81 (.A1(n_19), .A2(p_1[48]), .ZN(n_18));
   OR2_X1 i_82 (.A1(n_20), .A2(p_1[47]), .ZN(n_19));
   OR2_X1 i_83 (.A1(n_21), .A2(p_1[46]), .ZN(n_20));
   OR2_X1 i_84 (.A1(n_22), .A2(p_1[45]), .ZN(n_21));
   OR3_X1 i_85 (.A1(n_23), .A2(p_1[43]), .A3(p_1[44]), .ZN(n_22));
   NAND2_X1 i_86 (.A1(n_24), .A2(n_68), .ZN(n_23));
   NOR2_X1 i_87 (.A1(n_25), .A2(p_1[41]), .ZN(n_24));
   NAND2_X1 i_88 (.A1(n_26), .A2(n_67), .ZN(n_25));
   NOR3_X1 i_89 (.A1(n_28), .A2(p_1[38]), .A3(p_1[39]), .ZN(n_26));
   NOR2_X1 i_90 (.A1(n_28), .A2(p_1[38]), .ZN(n_27));
   OR2_X1 i_91 (.A1(n_29), .A2(p_1[37]), .ZN(n_28));
   NAND2_X1 i_92 (.A1(n_30), .A2(n_66), .ZN(n_29));
   NOR4_X1 i_93 (.A1(n_33), .A2(p_1[33]), .A3(p_1[34]), .A4(p_1[35]), .ZN(n_30));
   NOR3_X1 i_94 (.A1(n_33), .A2(p_1[33]), .A3(p_1[34]), .ZN(n_31));
   NOR2_X1 i_95 (.A1(n_33), .A2(p_1[33]), .ZN(n_32));
   OR2_X1 i_96 (.A1(n_34), .A2(p_1[32]), .ZN(n_33));
   NAND2_X1 i_97 (.A1(n_35), .A2(n_65), .ZN(n_34));
   NOR4_X1 i_98 (.A1(n_38), .A2(p_1[28]), .A3(p_1[29]), .A4(p_1[30]), .ZN(n_35));
   NOR3_X1 i_99 (.A1(n_38), .A2(p_1[28]), .A3(p_1[29]), .ZN(n_36));
   NOR2_X1 i_100 (.A1(n_38), .A2(p_1[28]), .ZN(n_37));
   OR2_X1 i_101 (.A1(n_39), .A2(p_1[27]), .ZN(n_38));
   NAND2_X1 i_102 (.A1(n_40), .A2(n_64), .ZN(n_39));
   NOR4_X1 i_103 (.A1(n_43), .A2(p_1[23]), .A3(p_1[24]), .A4(p_1[25]), .ZN(n_40));
   NOR3_X1 i_104 (.A1(n_43), .A2(p_1[23]), .A3(p_1[24]), .ZN(n_41));
   NOR2_X1 i_105 (.A1(n_43), .A2(p_1[23]), .ZN(n_42));
   OR2_X1 i_106 (.A1(n_44), .A2(p_1[22]), .ZN(n_43));
   NAND2_X1 i_107 (.A1(n_45), .A2(n_63), .ZN(n_44));
   NOR4_X1 i_108 (.A1(n_48), .A2(p_1[18]), .A3(p_1[19]), .A4(p_1[20]), .ZN(n_45));
   NOR3_X1 i_109 (.A1(n_48), .A2(p_1[18]), .A3(p_1[19]), .ZN(n_46));
   NOR2_X1 i_110 (.A1(n_48), .A2(p_1[18]), .ZN(n_47));
   OR2_X1 i_111 (.A1(n_49), .A2(p_1[17]), .ZN(n_48));
   OR2_X1 i_112 (.A1(n_50), .A2(p_1[16]), .ZN(n_49));
   OR3_X1 i_113 (.A1(n_51), .A2(p_1[14]), .A3(p_1[15]), .ZN(n_50));
   NAND2_X1 i_114 (.A1(n_52), .A2(n_62), .ZN(n_51));
   NOR2_X1 i_115 (.A1(n_53), .A2(p_1[12]), .ZN(n_52));
   NAND2_X1 i_116 (.A1(n_54), .A2(n_61), .ZN(n_53));
   NOR2_X1 i_117 (.A1(n_55), .A2(p_1[10]), .ZN(n_54));
   OR3_X1 i_118 (.A1(n_56), .A2(p_1[8]), .A3(p_1[9]), .ZN(n_55));
   OR2_X1 i_119 (.A1(n_57), .A2(p_1[7]), .ZN(n_56));
   OR3_X1 i_120 (.A1(n_58), .A2(p_1[5]), .A3(p_1[6]), .ZN(n_57));
   OR2_X1 i_121 (.A1(n_59), .A2(p_1[4]), .ZN(n_58));
   OR2_X1 i_122 (.A1(n_60), .A2(p_1[3]), .ZN(n_59));
   OR3_X1 i_123 (.A1(p_1[2]), .A2(p_1[1]), .A3(p_1[0]), .ZN(n_60));
   INV_X1 i_124 (.A(p_1[11]), .ZN(n_61));
   INV_X1 i_125 (.A(p_1[13]), .ZN(n_62));
   INV_X1 i_126 (.A(p_1[21]), .ZN(n_63));
   INV_X1 i_127 (.A(p_1[26]), .ZN(n_64));
   INV_X1 i_128 (.A(p_1[31]), .ZN(n_65));
   INV_X1 i_129 (.A(p_1[36]), .ZN(n_66));
   INV_X1 i_130 (.A(p_1[40]), .ZN(n_67));
   INV_X1 i_131 (.A(p_1[42]), .ZN(n_68));
   INV_X1 i_132 (.A(p_1[51]), .ZN(n_69));
   INV_X1 i_133 (.A(p_1[55]), .ZN(n_70));
   INV_X1 i_134 (.A(p_1[60]), .ZN(n_71));
   INV_X1 i_135 (.A(p_1[62]), .ZN(n_72));
endmodule

module booth_multiplier(clk, rst, en, a, b, c);
   input clk;
   input rst;
   input en;
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   wire n_64_0;
   wire n_64_3;
   wire n_64_4;
   wire n_64_5;
   wire n_64_6;
   wire n_64_7;
   wire n_64_8;
   wire n_64_9;
   wire n_64_10;
   wire n_64_11;
   wire n_64_12;
   wire n_64_13;
   wire n_64_14;
   wire n_64_15;
   wire n_64_16;
   wire n_64_17;
   wire n_64_18;
   wire n_64_19;
   wire n_64_20;
   wire n_64_21;
   wire n_64_22;
   wire n_64_23;
   wire n_64_24;
   wire n_64_25;
   wire n_64_26;
   wire n_64_27;
   wire n_64_28;
   wire n_64_29;
   wire n_64_30;
   wire n_64_31;
   wire n_64_32;
   wire n_64_33;
   wire n_64_34;
   wire n_64_35;
   wire n_64_36;
   wire n_64_37;
   wire n_64_38;
   wire n_64_39;
   wire n_64_40;
   wire n_64_41;
   wire n_64_42;
   wire n_64_43;
   wire n_64_44;
   wire n_64_45;
   wire n_64_46;
   wire n_64_47;
   wire n_64_48;
   wire n_64_49;
   wire n_64_50;
   wire n_64_51;
   wire n_64_52;
   wire n_64_53;
   wire n_64_54;
   wire n_64_55;
   wire n_64_56;
   wire n_64_57;
   wire n_64_58;
   wire n_64_59;
   wire n_64_60;
   wire n_64_61;
   wire n_64_62;
   wire n_64_63;
   wire n_64_64;
   wire n_64_65;
   wire n_64_66;
   wire n_64_67;
   wire n_64_68;
   wire n_64_69;
   wire n_64_70;
   wire n_64_71;
   wire n_64_72;
   wire n_64_73;
   wire n_64_74;
   wire n_64_75;
   wire n_64_76;
   wire n_64_77;
   wire n_64_78;
   wire n_64_79;
   wire n_64_80;
   wire n_64_81;
   wire n_64_82;
   wire n_64_83;
   wire n_64_84;
   wire n_64_85;
   wire n_64_86;
   wire n_64_87;
   wire n_64_88;
   wire n_64_89;
   wire n_64_90;
   wire n_64_91;
   wire n_64_92;
   wire n_64_93;
   wire n_64_94;
   wire n_64_95;
   wire n_64_96;
   wire n_64_97;
   wire n_64_98;
   wire n_64_99;
   wire n_64_100;
   wire n_64_101;
   wire n_64_102;
   wire n_64_103;
   wire n_64_104;
   wire n_64_105;
   wire n_64_106;
   wire n_64_107;
   wire n_64_108;
   wire n_64_109;
   wire n_64_110;
   wire n_64_111;
   wire n_64_112;
   wire n_64_113;
   wire n_64_114;
   wire n_64_115;
   wire n_64_116;
   wire n_64_117;
   wire n_64_118;
   wire n_64_119;
   wire n_64_120;
   wire n_64_121;
   wire n_64_122;
   wire n_64_123;
   wire n_64_124;
   wire n_64_125;
   wire n_64_126;
   wire n_64_127;
   wire n_64_128;
   wire n_64_129;
   wire n_64_130;
   wire n_64_131;
   wire n_64_132;
   wire n_64_133;
   wire n_64_134;
   wire n_64_135;
   wire n_64_136;
   wire n_64_137;
   wire n_64_138;
   wire n_64_139;
   wire n_64_140;
   wire n_64_141;
   wire n_64_142;
   wire n_64_143;
   wire n_64_144;
   wire n_64_145;
   wire n_64_146;
   wire n_64_147;
   wire n_64_148;
   wire n_64_149;
   wire n_64_150;
   wire n_64_151;
   wire n_64_152;
   wire n_64_153;
   wire n_64_154;
   wire n_64_155;
   wire n_64_156;
   wire n_64_157;
   wire n_64_158;
   wire n_64_159;
   wire n_64_160;
   wire n_64_161;
   wire n_64_162;
   wire n_64_163;
   wire n_64_164;
   wire n_64_165;
   wire n_64_166;
   wire n_64_167;
   wire n_64_168;
   wire n_64_169;
   wire n_64_170;
   wire n_64_171;
   wire n_64_172;
   wire n_64_173;
   wire n_64_174;
   wire n_64_175;
   wire n_64_176;
   wire n_64_177;
   wire n_64_178;
   wire n_64_179;
   wire n_64_180;
   wire n_64_181;
   wire n_64_182;
   wire n_64_183;
   wire n_64_184;
   wire n_64_185;
   wire n_64_186;
   wire n_64_187;
   wire n_64_188;
   wire n_64_189;
   wire n_64_190;
   wire n_64_191;
   wire n_64_192;
   wire [6:0]SC;
   wire [31:0]A;
   wire [31:0]multiplicand;
   wire [32:0]Q;
   wire out_sign;
   wire n_64_193;
   wire n_64_1;
   wire n_64_2;
   wire n_64_2_5;
   wire n_64_2_0;
   wire n_64_2_6;
   wire n_64_2_1;
   wire n_64_2_7;
   wire n_64_2_2;
   wire n_64_2_8;
   wire n_64_2_3;
   wire n_64_2_9;
   wire n_64_2_4;
   wire n_64_194;
   wire n_64_195;
   wire n_64_196;
   wire n_64_197;
   wire n_64_198;
   wire n_64_199;
   wire n_64_200;
   wire n_64_2_10;
   wire n_64_201;
   wire n_64_2_11;
   wire n_64_2_12;
   wire n_64_2_13;
   wire n_64_202;
   wire n_64_2_14;
   wire n_64_203;
   wire n_64_2_15;
   wire n_64_204;
   wire n_64_2_16;
   wire n_64_205;
   wire n_64_2_17;
   wire n_64_206;
   wire n_64_2_18;
   wire n_64_207;
   wire n_64_2_19;
   wire n_64_208;
   wire n_64_2_20;
   wire n_64_209;
   wire n_64_2_21;
   wire n_64_210;
   wire n_64_2_22;
   wire n_64_211;
   wire n_64_2_23;
   wire n_64_212;
   wire n_64_2_24;
   wire n_64_213;
   wire n_64_2_25;
   wire n_64_214;
   wire n_64_2_26;
   wire n_64_215;
   wire n_64_2_27;
   wire n_64_216;
   wire n_64_2_28;
   wire n_64_217;
   wire n_64_2_29;
   wire n_64_218;
   wire n_64_2_30;
   wire n_64_219;
   wire n_64_2_31;
   wire n_64_220;
   wire n_64_2_32;
   wire n_64_221;
   wire n_64_2_33;
   wire n_64_222;
   wire n_64_2_34;
   wire n_64_223;
   wire n_64_2_35;
   wire n_64_224;
   wire n_64_2_36;
   wire n_64_225;
   wire n_64_2_37;
   wire n_64_226;
   wire n_64_2_38;
   wire n_64_227;
   wire n_64_2_39;
   wire n_64_228;
   wire n_64_2_40;
   wire n_64_229;
   wire n_64_2_41;
   wire n_64_230;
   wire n_64_2_42;
   wire n_64_231;
   wire n_64_2_43;
   wire n_64_232;
   wire n_64_233;
   wire n_64_234;
   wire n_64_235;
   wire n_64_236;
   wire n_64_237;
   wire n_64_238;
   wire n_64_239;
   wire n_64_240;
   wire n_64_241;
   wire n_64_242;
   wire n_64_243;
   wire n_64_244;
   wire n_64_245;
   wire n_64_246;
   wire n_64_247;
   wire n_64_248;
   wire n_64_249;
   wire n_64_250;
   wire n_64_251;
   wire n_64_252;
   wire n_64_253;
   wire n_64_254;
   wire n_64_255;
   wire n_64_256;
   wire n_64_257;
   wire n_64_258;
   wire n_64_259;
   wire n_64_260;
   wire n_64_261;
   wire n_64_262;
   wire n_64_263;
   wire n_64_264;
   wire n_64_2_44;
   wire n_64_265;
   wire n_64_267;
   wire n_64_2_45;
   wire n_64_268;
   wire n_64_2_46;
   wire n_64_269;
   wire n_64_2_47;
   wire n_64_270;
   wire n_64_2_48;
   wire n_64_271;
   wire n_64_2_49;
   wire n_64_272;
   wire n_64_2_50;
   wire n_64_273;
   wire n_64_2_51;
   wire n_64_274;
   wire n_64_2_52;
   wire n_64_275;
   wire n_64_2_53;
   wire n_64_276;
   wire n_64_2_54;
   wire n_64_277;
   wire n_64_2_55;
   wire n_64_278;
   wire n_64_2_56;
   wire n_64_279;
   wire n_64_2_57;
   wire n_64_280;
   wire n_64_2_58;
   wire n_64_281;
   wire n_64_2_59;
   wire n_64_282;
   wire n_64_2_60;
   wire n_64_283;
   wire n_64_2_61;
   wire n_64_284;
   wire n_64_2_62;
   wire n_64_285;
   wire n_64_2_63;
   wire n_64_286;
   wire n_64_2_64;
   wire n_64_287;
   wire n_64_2_65;
   wire n_64_288;
   wire n_64_2_66;
   wire n_64_289;
   wire n_64_2_67;
   wire n_64_290;
   wire n_64_2_68;
   wire n_64_291;
   wire n_64_2_69;
   wire n_64_292;
   wire n_64_2_70;
   wire n_64_293;
   wire n_64_2_71;
   wire n_64_294;
   wire n_64_2_72;
   wire n_64_295;
   wire n_64_2_73;
   wire n_64_296;
   wire n_64_2_74;
   wire n_64_2_75;
   wire n_64_297;
   wire n_64_2_76;
   wire n_64_2_77;
   wire n_64_2_78;
   wire n_64_298;
   wire n_64_2_79;
   wire n_64_2_80;
   wire n_64_299;
   wire n_64_2_81;
   wire n_64_2_82;
   wire n_64_300;
   wire n_64_2_83;
   wire n_64_2_84;
   wire n_64_301;
   wire n_64_2_85;
   wire n_64_2_86;
   wire n_64_302;
   wire n_64_2_87;
   wire n_64_2_88;
   wire n_64_303;
   wire n_64_2_89;
   wire n_64_2_90;
   wire n_64_304;
   wire n_64_2_91;
   wire n_64_2_92;
   wire n_64_305;
   wire n_64_2_93;
   wire n_64_2_94;
   wire n_64_306;
   wire n_64_2_95;
   wire n_64_2_96;
   wire n_64_307;
   wire n_64_2_97;
   wire n_64_2_98;
   wire n_64_308;
   wire n_64_2_99;
   wire n_64_2_100;
   wire n_64_309;
   wire n_64_2_101;
   wire n_64_2_102;
   wire n_64_310;
   wire n_64_2_103;
   wire n_64_2_104;
   wire n_64_311;
   wire n_64_2_105;
   wire n_64_2_106;
   wire n_64_312;
   wire n_64_2_107;
   wire n_64_2_108;
   wire n_64_313;
   wire n_64_2_109;
   wire n_64_2_110;
   wire n_64_314;
   wire n_64_2_111;
   wire n_64_2_112;
   wire n_64_315;
   wire n_64_2_113;
   wire n_64_2_114;
   wire n_64_316;
   wire n_64_2_115;
   wire n_64_2_116;
   wire n_64_317;
   wire n_64_2_117;
   wire n_64_2_118;
   wire n_64_318;
   wire n_64_2_119;
   wire n_64_2_120;
   wire n_64_319;
   wire n_64_2_121;
   wire n_64_2_122;
   wire n_64_320;
   wire n_64_2_123;
   wire n_64_2_124;
   wire n_64_321;
   wire n_64_2_125;
   wire n_64_2_126;
   wire n_64_322;
   wire n_64_2_127;
   wire n_64_2_128;
   wire n_64_323;
   wire n_64_2_129;
   wire n_64_2_130;
   wire n_64_324;
   wire n_64_2_131;
   wire n_64_2_132;
   wire n_64_325;
   wire n_64_2_133;
   wire n_64_2_134;
   wire n_64_326;
   wire n_64_2_135;
   wire n_64_2_136;
   wire n_64_327;
   wire n_64_2_137;
   wire n_64_2_138;
   wire n_64_328;
   wire n_64_2_139;
   wire n_64_329;
   wire n_64_2_140;
   wire n_64_2_141;
   wire n_64_2_142;
   wire n_64_2_143;
   wire n_64_2_144;
   wire n_64_266;
   wire n_64_330;
   wire n_64_331;
   wire n_64_2_145;
   wire n_64_332;
   wire n_64_2_146;
   wire n_64_333;
   wire n_64_2_147;
   wire n_64_334;
   wire n_64_2_148;
   wire n_64_335;
   wire n_64_2_149;
   wire n_64_336;
   wire n_64_2_150;
   wire n_64_337;
   wire n_64_2_151;
   wire n_64_338;
   wire n_64_2_152;
   wire n_64_339;
   wire n_64_2_153;
   wire n_64_340;
   wire n_64_2_154;
   wire n_64_341;
   wire n_64_2_155;
   wire n_64_342;
   wire n_64_2_156;
   wire n_64_343;
   wire n_64_2_157;
   wire n_64_344;
   wire n_64_2_158;
   wire n_64_345;
   wire n_64_2_159;
   wire n_64_346;
   wire n_64_2_160;
   wire n_64_347;
   wire n_64_2_161;
   wire n_64_348;
   wire n_64_2_162;
   wire n_64_349;
   wire n_64_2_163;
   wire n_64_350;
   wire n_64_2_164;
   wire n_64_351;
   wire n_64_2_165;
   wire n_64_352;
   wire n_64_2_166;
   wire n_64_353;
   wire n_64_2_167;
   wire n_64_354;
   wire n_64_2_168;
   wire n_64_355;
   wire n_64_2_169;
   wire n_64_356;
   wire n_64_2_170;
   wire n_64_357;
   wire n_64_2_171;
   wire n_64_358;
   wire n_64_2_172;
   wire n_64_359;
   wire n_64_2_173;
   wire n_64_360;
   wire n_64_2_174;
   wire n_64_2_175;
   wire n_64_361;
   wire n_64_2_176;
   wire n_64_2_177;
   wire n_64_2_178;
   wire n_64_2_179;
   wire n_64_2_180;
   wire n_64_362;
   wire n_64_2_181;
   wire n_64_363;
   wire n_64_2_182;
   wire n_64_2_183;
   wire n_64_2_184;
   wire n_64_2_185;
   wire n_64_2_186;
   wire n_64_2_187;
   wire n_64_2_188;

   TBUF_X1 i_0 (.A(n_64), .EN(n_0), .Z(c[0]));
   TBUF_X1 i_1 (.A(n_63), .EN(n_0), .Z(c[1]));
   TBUF_X1 i_2 (.A(n_62), .EN(n_0), .Z(c[2]));
   TBUF_X1 i_3 (.A(n_61), .EN(n_0), .Z(c[3]));
   TBUF_X1 i_4 (.A(n_60), .EN(n_0), .Z(c[4]));
   TBUF_X1 i_5 (.A(n_59), .EN(n_0), .Z(c[5]));
   TBUF_X1 i_6 (.A(n_58), .EN(n_0), .Z(c[6]));
   TBUF_X1 i_7 (.A(n_57), .EN(n_0), .Z(c[7]));
   TBUF_X1 i_8 (.A(n_56), .EN(n_0), .Z(c[8]));
   TBUF_X1 i_9 (.A(n_55), .EN(n_0), .Z(c[9]));
   TBUF_X1 i_10 (.A(n_54), .EN(n_0), .Z(c[10]));
   TBUF_X1 i_11 (.A(n_53), .EN(n_0), .Z(c[11]));
   TBUF_X1 i_12 (.A(n_52), .EN(n_0), .Z(c[12]));
   TBUF_X1 i_13 (.A(n_51), .EN(n_0), .Z(c[13]));
   TBUF_X1 i_14 (.A(n_50), .EN(n_0), .Z(c[14]));
   TBUF_X1 i_15 (.A(n_49), .EN(n_0), .Z(c[15]));
   TBUF_X1 i_16 (.A(n_48), .EN(n_0), .Z(c[16]));
   TBUF_X1 i_17 (.A(n_47), .EN(n_0), .Z(c[17]));
   TBUF_X1 i_18 (.A(n_46), .EN(n_0), .Z(c[18]));
   TBUF_X1 i_19 (.A(n_45), .EN(n_0), .Z(c[19]));
   TBUF_X1 i_20 (.A(n_44), .EN(n_0), .Z(c[20]));
   TBUF_X1 i_21 (.A(n_43), .EN(n_0), .Z(c[21]));
   TBUF_X1 i_22 (.A(n_42), .EN(n_0), .Z(c[22]));
   TBUF_X1 i_23 (.A(n_41), .EN(n_0), .Z(c[23]));
   TBUF_X1 i_24 (.A(n_40), .EN(n_0), .Z(c[24]));
   TBUF_X1 i_25 (.A(n_39), .EN(n_0), .Z(c[25]));
   TBUF_X1 i_26 (.A(n_38), .EN(n_0), .Z(c[26]));
   TBUF_X1 i_27 (.A(n_37), .EN(n_0), .Z(c[27]));
   TBUF_X1 i_28 (.A(n_36), .EN(n_0), .Z(c[28]));
   TBUF_X1 i_29 (.A(n_35), .EN(n_0), .Z(c[29]));
   TBUF_X1 i_30 (.A(n_34), .EN(n_0), .Z(c[30]));
   TBUF_X1 i_31 (.A(n_33), .EN(n_0), .Z(c[31]));
   TBUF_X1 i_32 (.A(n_32), .EN(n_0), .Z(c[32]));
   TBUF_X1 i_33 (.A(n_31), .EN(n_0), .Z(c[33]));
   TBUF_X1 i_34 (.A(n_30), .EN(n_0), .Z(c[34]));
   TBUF_X1 i_35 (.A(n_29), .EN(n_0), .Z(c[35]));
   TBUF_X1 i_36 (.A(n_28), .EN(n_0), .Z(c[36]));
   TBUF_X1 i_37 (.A(n_27), .EN(n_0), .Z(c[37]));
   TBUF_X1 i_38 (.A(n_26), .EN(n_0), .Z(c[38]));
   TBUF_X1 i_39 (.A(n_25), .EN(n_0), .Z(c[39]));
   TBUF_X1 i_40 (.A(n_24), .EN(n_0), .Z(c[40]));
   TBUF_X1 i_41 (.A(n_23), .EN(n_0), .Z(c[41]));
   TBUF_X1 i_42 (.A(n_22), .EN(n_0), .Z(c[42]));
   TBUF_X1 i_43 (.A(n_21), .EN(n_0), .Z(c[43]));
   TBUF_X1 i_44 (.A(n_20), .EN(n_0), .Z(c[44]));
   TBUF_X1 i_45 (.A(n_19), .EN(n_0), .Z(c[45]));
   TBUF_X1 i_46 (.A(n_18), .EN(n_0), .Z(c[46]));
   TBUF_X1 i_47 (.A(n_17), .EN(n_0), .Z(c[47]));
   TBUF_X1 i_48 (.A(n_16), .EN(n_0), .Z(c[48]));
   TBUF_X1 i_49 (.A(n_15), .EN(n_0), .Z(c[49]));
   TBUF_X1 i_50 (.A(n_14), .EN(n_0), .Z(c[50]));
   TBUF_X1 i_51 (.A(n_13), .EN(n_0), .Z(c[51]));
   TBUF_X1 i_52 (.A(n_12), .EN(n_0), .Z(c[52]));
   TBUF_X1 i_53 (.A(n_11), .EN(n_0), .Z(c[53]));
   TBUF_X1 i_54 (.A(n_10), .EN(n_0), .Z(c[54]));
   TBUF_X1 i_55 (.A(n_9), .EN(n_0), .Z(c[55]));
   TBUF_X1 i_56 (.A(n_8), .EN(n_0), .Z(c[56]));
   TBUF_X1 i_57 (.A(n_7), .EN(n_0), .Z(c[57]));
   TBUF_X1 i_58 (.A(n_6), .EN(n_0), .Z(c[58]));
   TBUF_X1 i_59 (.A(n_5), .EN(n_0), .Z(c[59]));
   TBUF_X1 i_60 (.A(n_4), .EN(n_0), .Z(c[60]));
   TBUF_X1 i_61 (.A(n_3), .EN(n_0), .Z(c[61]));
   TBUF_X1 i_62 (.A(n_2), .EN(n_0), .Z(c[62]));
   TBUF_X1 i_63 (.A(n_1), .EN(n_0), .Z(c[63]));
   INV_X1 i_64_0 (.A(n_64_3), .ZN(n_0));
   CLKGATETST_X1 clk_gate_c_reg (.CK(clk), .E(n_64_362), .SE(1'b0), .GCK(n_64_0));
   DFF_X1 \c_reg[63]  (.D(n_64_264), .CK(n_64_0), .Q(n_1), .QN());
   DFF_X1 \c_reg[62]  (.D(n_64_263), .CK(n_64_0), .Q(n_2), .QN());
   DFF_X1 \c_reg[61]  (.D(n_64_262), .CK(n_64_0), .Q(n_3), .QN());
   DFF_X1 \c_reg[60]  (.D(n_64_261), .CK(n_64_0), .Q(n_4), .QN());
   DFF_X1 \c_reg[59]  (.D(n_64_260), .CK(n_64_0), .Q(n_5), .QN());
   DFF_X1 \c_reg[58]  (.D(n_64_259), .CK(n_64_0), .Q(n_6), .QN());
   DFF_X1 \c_reg[57]  (.D(n_64_258), .CK(n_64_0), .Q(n_7), .QN());
   DFF_X1 \c_reg[56]  (.D(n_64_257), .CK(n_64_0), .Q(n_8), .QN());
   DFF_X1 \c_reg[55]  (.D(n_64_256), .CK(n_64_0), .Q(n_9), .QN());
   DFF_X1 \c_reg[54]  (.D(n_64_255), .CK(n_64_0), .Q(n_10), .QN());
   DFF_X1 \c_reg[53]  (.D(n_64_254), .CK(n_64_0), .Q(n_11), .QN());
   DFF_X1 \c_reg[52]  (.D(n_64_253), .CK(n_64_0), .Q(n_12), .QN());
   DFF_X1 \c_reg[51]  (.D(n_64_252), .CK(n_64_0), .Q(n_13), .QN());
   DFF_X1 \c_reg[50]  (.D(n_64_251), .CK(n_64_0), .Q(n_14), .QN());
   DFF_X1 \c_reg[49]  (.D(n_64_250), .CK(n_64_0), .Q(n_15), .QN());
   DFF_X1 \c_reg[48]  (.D(n_64_249), .CK(n_64_0), .Q(n_16), .QN());
   DFF_X1 \c_reg[47]  (.D(n_64_248), .CK(n_64_0), .Q(n_17), .QN());
   DFF_X1 \c_reg[46]  (.D(n_64_247), .CK(n_64_0), .Q(n_18), .QN());
   DFF_X1 \c_reg[45]  (.D(n_64_246), .CK(n_64_0), .Q(n_19), .QN());
   DFF_X1 \c_reg[44]  (.D(n_64_245), .CK(n_64_0), .Q(n_20), .QN());
   DFF_X1 \c_reg[43]  (.D(n_64_244), .CK(n_64_0), .Q(n_21), .QN());
   DFF_X1 \c_reg[42]  (.D(n_64_243), .CK(n_64_0), .Q(n_22), .QN());
   DFF_X1 \c_reg[41]  (.D(n_64_242), .CK(n_64_0), .Q(n_23), .QN());
   DFF_X1 \c_reg[40]  (.D(n_64_241), .CK(n_64_0), .Q(n_24), .QN());
   DFF_X1 \c_reg[39]  (.D(n_64_240), .CK(n_64_0), .Q(n_25), .QN());
   DFF_X1 \c_reg[38]  (.D(n_64_239), .CK(n_64_0), .Q(n_26), .QN());
   DFF_X1 \c_reg[37]  (.D(n_64_238), .CK(n_64_0), .Q(n_27), .QN());
   DFF_X1 \c_reg[36]  (.D(n_64_237), .CK(n_64_0), .Q(n_28), .QN());
   DFF_X1 \c_reg[35]  (.D(n_64_236), .CK(n_64_0), .Q(n_29), .QN());
   DFF_X1 \c_reg[34]  (.D(n_64_235), .CK(n_64_0), .Q(n_30), .QN());
   DFF_X1 \c_reg[33]  (.D(n_64_234), .CK(n_64_0), .Q(n_31), .QN());
   DFF_X1 \c_reg[32]  (.D(n_64_233), .CK(n_64_0), .Q(n_32), .QN());
   DFF_X1 \c_reg[31]  (.D(n_64_232), .CK(n_64_0), .Q(n_33), .QN());
   DFF_X1 \c_reg[30]  (.D(n_64_231), .CK(n_64_0), .Q(n_34), .QN());
   DFF_X1 \c_reg[29]  (.D(n_64_230), .CK(n_64_0), .Q(n_35), .QN());
   DFF_X1 \c_reg[28]  (.D(n_64_229), .CK(n_64_0), .Q(n_36), .QN());
   DFF_X1 \c_reg[27]  (.D(n_64_228), .CK(n_64_0), .Q(n_37), .QN());
   DFF_X1 \c_reg[26]  (.D(n_64_227), .CK(n_64_0), .Q(n_38), .QN());
   DFF_X1 \c_reg[25]  (.D(n_64_226), .CK(n_64_0), .Q(n_39), .QN());
   DFF_X1 \c_reg[24]  (.D(n_64_225), .CK(n_64_0), .Q(n_40), .QN());
   DFF_X1 \c_reg[23]  (.D(n_64_224), .CK(n_64_0), .Q(n_41), .QN());
   DFF_X1 \c_reg[22]  (.D(n_64_223), .CK(n_64_0), .Q(n_42), .QN());
   DFF_X1 \c_reg[21]  (.D(n_64_222), .CK(n_64_0), .Q(n_43), .QN());
   DFF_X1 \c_reg[20]  (.D(n_64_221), .CK(n_64_0), .Q(n_44), .QN());
   DFF_X1 \c_reg[19]  (.D(n_64_220), .CK(n_64_0), .Q(n_45), .QN());
   DFF_X1 \c_reg[18]  (.D(n_64_219), .CK(n_64_0), .Q(n_46), .QN());
   DFF_X1 \c_reg[17]  (.D(n_64_218), .CK(n_64_0), .Q(n_47), .QN());
   DFF_X1 \c_reg[16]  (.D(n_64_217), .CK(n_64_0), .Q(n_48), .QN());
   DFF_X1 \c_reg[15]  (.D(n_64_216), .CK(n_64_0), .Q(n_49), .QN());
   DFF_X1 \c_reg[14]  (.D(n_64_215), .CK(n_64_0), .Q(n_50), .QN());
   DFF_X1 \c_reg[13]  (.D(n_64_214), .CK(n_64_0), .Q(n_51), .QN());
   DFF_X1 \c_reg[12]  (.D(n_64_213), .CK(n_64_0), .Q(n_52), .QN());
   DFF_X1 \c_reg[11]  (.D(n_64_212), .CK(n_64_0), .Q(n_53), .QN());
   DFF_X1 \c_reg[10]  (.D(n_64_211), .CK(n_64_0), .Q(n_54), .QN());
   DFF_X1 \c_reg[9]  (.D(n_64_210), .CK(n_64_0), .Q(n_55), .QN());
   DFF_X1 \c_reg[8]  (.D(n_64_209), .CK(n_64_0), .Q(n_56), .QN());
   DFF_X1 \c_reg[7]  (.D(n_64_208), .CK(n_64_0), .Q(n_57), .QN());
   DFF_X1 \c_reg[6]  (.D(n_64_207), .CK(n_64_0), .Q(n_58), .QN());
   DFF_X1 \c_reg[5]  (.D(n_64_206), .CK(n_64_0), .Q(n_59), .QN());
   DFF_X1 \c_reg[4]  (.D(n_64_205), .CK(n_64_0), .Q(n_60), .QN());
   DFF_X1 \c_reg[3]  (.D(n_64_204), .CK(n_64_0), .Q(n_61), .QN());
   DFF_X1 \c_reg[2]  (.D(n_64_203), .CK(n_64_0), .Q(n_62), .QN());
   DFF_X1 \c_reg[1]  (.D(n_64_202), .CK(n_64_0), .Q(n_63), .QN());
   DFF_X1 \c_reg[0]  (.D(n_64_267), .CK(n_64_0), .Q(n_64), .QN());
   DFFR_X1 i_64_64 (.D(n_64_363), .RN(n_64_193), .CK(clk), .Q(n_64_3), .QN());
   datapath i_64_194 (.p_0({n_64_34, n_64_33, n_64_32, n_64_31, n_64_30, n_64_29, 
      n_64_28, n_64_27, n_64_26, n_64_25, n_64_24, n_64_23, n_64_22, n_64_21, 
      n_64_20, n_64_19, n_64_18, n_64_17, n_64_16, n_64_15, n_64_14, n_64_13, 
      n_64_12, n_64_11, n_64_10, n_64_9, n_64_8, n_64_7, n_64_6, n_64_5, n_64_4, 
      uc_0}), .a(a));
   datapath__0_127 i_64_196 (.A({A[31], uc_1, A[29], A[28], A[27], A[26], A[25], 
      A[24], A[23], A[22], A[21], A[20], A[19], A[18], A[17], A[16], A[15], 
      A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], 
      A[3], A[2], A[1], A[0]}), .p_0({n_64_66, n_64_65, n_64_64, n_64_63, 
      n_64_62, n_64_61, n_64_60, n_64_59, n_64_58, n_64_57, n_64_56, n_64_55, 
      n_64_54, n_64_53, n_64_52, n_64_51, n_64_50, n_64_49, n_64_48, n_64_47, 
      n_64_46, n_64_45, n_64_44, n_64_43, n_64_42, n_64_41, n_64_40, n_64_39, 
      n_64_38, n_64_37, n_64_36, n_64_35}), .multiplicand({n_64_361, n_64_360, 
      n_64_359, n_64_358, n_64_357, n_64_356, n_64_355, n_64_354, n_64_353, 
      n_64_352, n_64_351, n_64_350, n_64_349, n_64_348, n_64_347, n_64_346, 
      n_64_345, n_64_344, n_64_343, n_64_342, n_64_341, n_64_340, n_64_339, 
      n_64_338, n_64_337, n_64_336, n_64_335, n_64_334, n_64_333, n_64_332, 
      n_64_331, n_64_330}));
   datapath__0_128 i_64_197 (.multiplicand({n_64_361, n_64_360, n_64_359, 
      n_64_358, n_64_357, n_64_356, n_64_355, n_64_354, n_64_353, n_64_352, 
      n_64_351, n_64_350, n_64_349, n_64_348, n_64_347, n_64_346, n_64_345, 
      n_64_344, n_64_343, n_64_342, n_64_341, n_64_340, n_64_339, n_64_338, 
      n_64_337, n_64_336, n_64_335, n_64_334, n_64_333, n_64_332, n_64_331, 
      n_64_330}), .A({A[31], uc_2, A[29], A[28], A[27], A[26], A[25], A[24], 
      A[23], A[22], A[21], A[20], A[19], A[18], A[17], A[16], A[15], A[14], 
      A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], 
      A[1], A[0]}), .p_0({n_64_98, n_64_97, n_64_96, n_64_95, n_64_94, n_64_93, 
      n_64_92, n_64_91, n_64_90, n_64_89, n_64_88, n_64_87, n_64_86, n_64_85, 
      n_64_84, n_64_83, n_64_82, n_64_81, n_64_80, n_64_79, n_64_78, n_64_77, 
      n_64_76, n_64_75, n_64_74, n_64_73, n_64_72, n_64_71, n_64_70, n_64_69, 
      n_64_68, n_64_67}));
   datapath__0_129 i_64_198 (.p_0({n_64_129, n_64_128, n_64_127, n_64_126, 
      n_64_125, n_64_124, n_64_123, n_64_122, n_64_121, n_64_120, n_64_119, 
      n_64_118, n_64_117, n_64_116, n_64_115, n_64_114, n_64_113, n_64_112, 
      n_64_111, n_64_110, n_64_109, n_64_108, n_64_107, n_64_106, n_64_105, 
      n_64_104, n_64_103, n_64_102, n_64_101, n_64_100, n_64_99, uc_3}), 
      .b(b));
   datapath__0_132 i_64_201 (.p_0({n_64_192, n_64_191, n_64_190, n_64_189, 
      n_64_188, n_64_187, n_64_186, n_64_185, n_64_184, n_64_183, n_64_182, 
      n_64_181, n_64_180, n_64_179, n_64_178, n_64_177, n_64_176, n_64_175, 
      n_64_174, n_64_173, n_64_172, n_64_171, n_64_170, n_64_169, n_64_168, 
      n_64_167, n_64_166, n_64_165, n_64_164, n_64_163, n_64_162, n_64_161, 
      n_64_160, n_64_159, n_64_158, n_64_157, n_64_156, n_64_155, n_64_154, 
      n_64_153, n_64_152, n_64_151, n_64_150, n_64_149, n_64_148, n_64_147, 
      n_64_146, n_64_145, n_64_144, n_64_143, n_64_142, n_64_141, n_64_140, 
      n_64_139, n_64_138, n_64_137, n_64_136, n_64_135, n_64_134, n_64_133, 
      n_64_132, n_64_131, n_64_130, uc_4}), .p_1({1'b0, n_64_329, n_64_328, 
      n_64_327, n_64_326, n_64_325, n_64_324, n_64_323, n_64_322, n_64_321, 
      n_64_320, n_64_319, n_64_318, n_64_317, n_64_316, n_64_315, n_64_314, 
      n_64_313, n_64_312, n_64_311, n_64_310, n_64_309, n_64_308, n_64_307, 
      n_64_306, n_64_305, n_64_304, n_64_303, n_64_302, n_64_301, n_64_300, 
      n_64_299, n_64_298, n_64_297, n_64_296, n_64_295, n_64_294, n_64_293, 
      n_64_292, n_64_291, n_64_290, n_64_289, n_64_288, n_64_287, n_64_286, 
      n_64_285, n_64_284, n_64_283, n_64_282, n_64_281, n_64_280, n_64_279, 
      n_64_278, n_64_277, n_64_276, n_64_275, n_64_274, n_64_273, n_64_272, 
      n_64_271, n_64_270, n_64_269, n_64_268, n_64_267}));
   DFFR_X1 \SC_reg[6]  (.D(n_64_200), .RN(n_64_193), .CK(n_64_1), .Q(SC[6]), 
      .QN());
   DFFR_X1 \SC_reg[5]  (.D(n_64_199), .RN(n_64_193), .CK(n_64_1), .Q(SC[5]), 
      .QN());
   DFFR_X1 \SC_reg[4]  (.D(n_64_198), .RN(n_64_193), .CK(n_64_1), .Q(SC[4]), 
      .QN());
   DFFR_X1 \SC_reg[3]  (.D(n_64_197), .RN(n_64_193), .CK(n_64_1), .Q(SC[3]), 
      .QN());
   DFFR_X1 \SC_reg[2]  (.D(n_64_196), .RN(n_64_193), .CK(n_64_1), .Q(SC[2]), 
      .QN());
   DFFR_X1 \SC_reg[1]  (.D(n_64_195), .RN(n_64_193), .CK(n_64_1), .Q(SC[1]), 
      .QN());
   DFFR_X1 \SC_reg[0]  (.D(n_64_194), .RN(n_64_193), .CK(n_64_1), .Q(SC[0]), 
      .QN());
   DFFR_X1 \A_reg[31]  (.D(n_64_329), .RN(n_64_193), .CK(n_64_1), .Q(A[31]), 
      .QN());
   DFFR_X1 \A_reg[29]  (.D(n_64_328), .RN(n_64_193), .CK(n_64_1), .Q(A[29]), 
      .QN());
   DFFR_X1 \A_reg[28]  (.D(n_64_327), .RN(n_64_193), .CK(n_64_1), .Q(A[28]), 
      .QN());
   DFFR_X1 \A_reg[27]  (.D(n_64_326), .RN(n_64_193), .CK(n_64_1), .Q(A[27]), 
      .QN());
   DFFR_X1 \A_reg[26]  (.D(n_64_325), .RN(n_64_193), .CK(n_64_1), .Q(A[26]), 
      .QN());
   DFFR_X1 \A_reg[25]  (.D(n_64_324), .RN(n_64_193), .CK(n_64_1), .Q(A[25]), 
      .QN());
   DFFR_X1 \A_reg[24]  (.D(n_64_323), .RN(n_64_193), .CK(n_64_1), .Q(A[24]), 
      .QN());
   DFFR_X1 \A_reg[23]  (.D(n_64_322), .RN(n_64_193), .CK(n_64_1), .Q(A[23]), 
      .QN());
   DFFR_X1 \A_reg[22]  (.D(n_64_321), .RN(n_64_193), .CK(n_64_1), .Q(A[22]), 
      .QN());
   DFFR_X1 \A_reg[21]  (.D(n_64_320), .RN(n_64_193), .CK(n_64_1), .Q(A[21]), 
      .QN());
   DFFR_X1 \A_reg[20]  (.D(n_64_319), .RN(n_64_193), .CK(n_64_1), .Q(A[20]), 
      .QN());
   DFFR_X1 \A_reg[19]  (.D(n_64_318), .RN(n_64_193), .CK(n_64_1), .Q(A[19]), 
      .QN());
   DFFR_X1 \A_reg[18]  (.D(n_64_317), .RN(n_64_193), .CK(n_64_1), .Q(A[18]), 
      .QN());
   DFFR_X1 \A_reg[17]  (.D(n_64_316), .RN(n_64_193), .CK(n_64_1), .Q(A[17]), 
      .QN());
   DFFR_X1 \A_reg[16]  (.D(n_64_315), .RN(n_64_193), .CK(n_64_1), .Q(A[16]), 
      .QN());
   DFFR_X1 \A_reg[15]  (.D(n_64_314), .RN(n_64_193), .CK(n_64_1), .Q(A[15]), 
      .QN());
   DFFR_X1 \A_reg[14]  (.D(n_64_313), .RN(n_64_193), .CK(n_64_1), .Q(A[14]), 
      .QN());
   DFFR_X1 \A_reg[13]  (.D(n_64_312), .RN(n_64_193), .CK(n_64_1), .Q(A[13]), 
      .QN());
   DFFR_X1 \A_reg[12]  (.D(n_64_311), .RN(n_64_193), .CK(n_64_1), .Q(A[12]), 
      .QN());
   DFFR_X1 \A_reg[11]  (.D(n_64_310), .RN(n_64_193), .CK(n_64_1), .Q(A[11]), 
      .QN());
   DFFR_X1 \A_reg[10]  (.D(n_64_309), .RN(n_64_193), .CK(n_64_1), .Q(A[10]), 
      .QN());
   DFFR_X1 \A_reg[9]  (.D(n_64_308), .RN(n_64_193), .CK(n_64_1), .Q(A[9]), .QN());
   DFFR_X1 \A_reg[8]  (.D(n_64_307), .RN(n_64_193), .CK(n_64_1), .Q(A[8]), .QN());
   DFFR_X1 \A_reg[7]  (.D(n_64_306), .RN(n_64_193), .CK(n_64_1), .Q(A[7]), .QN());
   DFFR_X1 \A_reg[6]  (.D(n_64_305), .RN(n_64_193), .CK(n_64_1), .Q(A[6]), .QN());
   DFFR_X1 \A_reg[5]  (.D(n_64_304), .RN(n_64_193), .CK(n_64_1), .Q(A[5]), .QN());
   DFFR_X1 \A_reg[4]  (.D(n_64_303), .RN(n_64_193), .CK(n_64_1), .Q(A[4]), .QN());
   DFFR_X1 \A_reg[3]  (.D(n_64_302), .RN(n_64_193), .CK(n_64_1), .Q(A[3]), .QN());
   DFFR_X1 \A_reg[2]  (.D(n_64_301), .RN(n_64_193), .CK(n_64_1), .Q(A[2]), .QN());
   DFFR_X1 \A_reg[1]  (.D(n_64_300), .RN(n_64_193), .CK(n_64_1), .Q(A[1]), .QN());
   DFFR_X1 \A_reg[0]  (.D(n_64_299), .RN(n_64_193), .CK(n_64_1), .Q(A[0]), .QN());
   DFF_X1 \multiplicand_reg[31]  (.D(n_64_361), .CK(n_64_2), .Q(multiplicand[31]), 
      .QN());
   DFF_X1 \multiplicand_reg[30]  (.D(n_64_360), .CK(n_64_2), .Q(multiplicand[30]), 
      .QN());
   DFF_X1 \multiplicand_reg[29]  (.D(n_64_359), .CK(n_64_2), .Q(multiplicand[29]), 
      .QN());
   DFF_X1 \multiplicand_reg[28]  (.D(n_64_358), .CK(n_64_2), .Q(multiplicand[28]), 
      .QN());
   DFF_X1 \multiplicand_reg[27]  (.D(n_64_357), .CK(n_64_2), .Q(multiplicand[27]), 
      .QN());
   DFF_X1 \multiplicand_reg[26]  (.D(n_64_356), .CK(n_64_2), .Q(multiplicand[26]), 
      .QN());
   DFF_X1 \multiplicand_reg[25]  (.D(n_64_355), .CK(n_64_2), .Q(multiplicand[25]), 
      .QN());
   DFF_X1 \multiplicand_reg[24]  (.D(n_64_354), .CK(n_64_2), .Q(multiplicand[24]), 
      .QN());
   DFF_X1 \multiplicand_reg[23]  (.D(n_64_353), .CK(n_64_2), .Q(multiplicand[23]), 
      .QN());
   DFF_X1 \multiplicand_reg[22]  (.D(n_64_352), .CK(n_64_2), .Q(multiplicand[22]), 
      .QN());
   DFF_X1 \multiplicand_reg[21]  (.D(n_64_351), .CK(n_64_2), .Q(multiplicand[21]), 
      .QN());
   DFF_X1 \multiplicand_reg[20]  (.D(n_64_350), .CK(n_64_2), .Q(multiplicand[20]), 
      .QN());
   DFF_X1 \multiplicand_reg[19]  (.D(n_64_349), .CK(n_64_2), .Q(multiplicand[19]), 
      .QN());
   DFF_X1 \multiplicand_reg[18]  (.D(n_64_348), .CK(n_64_2), .Q(multiplicand[18]), 
      .QN());
   DFF_X1 \multiplicand_reg[17]  (.D(n_64_347), .CK(n_64_2), .Q(multiplicand[17]), 
      .QN());
   DFF_X1 \multiplicand_reg[16]  (.D(n_64_346), .CK(n_64_2), .Q(multiplicand[16]), 
      .QN());
   DFF_X1 \multiplicand_reg[15]  (.D(n_64_345), .CK(n_64_2), .Q(multiplicand[15]), 
      .QN());
   DFF_X1 \multiplicand_reg[14]  (.D(n_64_344), .CK(n_64_2), .Q(multiplicand[14]), 
      .QN());
   DFF_X1 \multiplicand_reg[13]  (.D(n_64_343), .CK(n_64_2), .Q(multiplicand[13]), 
      .QN());
   DFF_X1 \multiplicand_reg[12]  (.D(n_64_342), .CK(n_64_2), .Q(multiplicand[12]), 
      .QN());
   DFF_X1 \multiplicand_reg[11]  (.D(n_64_341), .CK(n_64_2), .Q(multiplicand[11]), 
      .QN());
   DFF_X1 \multiplicand_reg[10]  (.D(n_64_340), .CK(n_64_2), .Q(multiplicand[10]), 
      .QN());
   DFF_X1 \multiplicand_reg[9]  (.D(n_64_339), .CK(n_64_2), .Q(multiplicand[9]), 
      .QN());
   DFF_X1 \multiplicand_reg[8]  (.D(n_64_338), .CK(n_64_2), .Q(multiplicand[8]), 
      .QN());
   DFF_X1 \multiplicand_reg[7]  (.D(n_64_337), .CK(n_64_2), .Q(multiplicand[7]), 
      .QN());
   DFF_X1 \multiplicand_reg[6]  (.D(n_64_336), .CK(n_64_2), .Q(multiplicand[6]), 
      .QN());
   DFF_X1 \multiplicand_reg[5]  (.D(n_64_335), .CK(n_64_2), .Q(multiplicand[5]), 
      .QN());
   DFF_X1 \multiplicand_reg[4]  (.D(n_64_334), .CK(n_64_2), .Q(multiplicand[4]), 
      .QN());
   DFF_X1 \multiplicand_reg[3]  (.D(n_64_333), .CK(n_64_2), .Q(multiplicand[3]), 
      .QN());
   DFF_X1 \multiplicand_reg[2]  (.D(n_64_332), .CK(n_64_2), .Q(multiplicand[2]), 
      .QN());
   DFF_X1 \multiplicand_reg[1]  (.D(n_64_331), .CK(n_64_2), .Q(multiplicand[1]), 
      .QN());
   DFF_X1 \multiplicand_reg[0]  (.D(n_64_330), .CK(n_64_2), .Q(multiplicand[0]), 
      .QN());
   DFF_X1 \Q_reg[32]  (.D(n_64_298), .CK(n_64_2), .Q(Q[32]), .QN());
   DFF_X1 \Q_reg[31]  (.D(n_64_297), .CK(n_64_2), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_64_296), .CK(n_64_2), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_64_295), .CK(n_64_2), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_64_294), .CK(n_64_2), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_64_293), .CK(n_64_2), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_64_292), .CK(n_64_2), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_64_291), .CK(n_64_2), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_64_290), .CK(n_64_2), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_64_289), .CK(n_64_2), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_64_288), .CK(n_64_2), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_64_287), .CK(n_64_2), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_64_286), .CK(n_64_2), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_64_285), .CK(n_64_2), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_64_284), .CK(n_64_2), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_64_283), .CK(n_64_2), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_64_282), .CK(n_64_2), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_64_281), .CK(n_64_2), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_64_280), .CK(n_64_2), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_64_279), .CK(n_64_2), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_64_278), .CK(n_64_2), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_64_277), .CK(n_64_2), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_64_276), .CK(n_64_2), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_64_275), .CK(n_64_2), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_64_274), .CK(n_64_2), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_64_273), .CK(n_64_2), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_64_272), .CK(n_64_2), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_64_271), .CK(n_64_2), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_64_270), .CK(n_64_2), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_64_269), .CK(n_64_2), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_64_268), .CK(n_64_2), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_64_267), .CK(n_64_2), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_64_266), .CK(n_64_2), .Q(Q[0]), .QN());
   DFF_X1 out_sign_reg (.D(n_64_201), .CK(n_64_2), .Q(out_sign), .QN());
   INV_X1 i_64_1_0 (.A(rst), .ZN(n_64_193));
   CLKGATETST_X1 clk_gate_SC_reg (.CK(clk), .E(en), .SE(1'b0), .GCK(n_64_1));
   CLKGATETST_X1 clk_gate_out_sign_reg (.CK(clk), .E(n_64_265), .SE(1'b0), 
      .GCK(n_64_2));
   HA_X1 i_64_2_0 (.A(SC[1]), .B(SC[0]), .CO(n_64_2_0), .S(n_64_2_5));
   HA_X1 i_64_2_1 (.A(SC[2]), .B(n_64_2_0), .CO(n_64_2_1), .S(n_64_2_6));
   HA_X1 i_64_2_2 (.A(SC[3]), .B(n_64_2_1), .CO(n_64_2_2), .S(n_64_2_7));
   HA_X1 i_64_2_3 (.A(SC[4]), .B(n_64_2_2), .CO(n_64_2_3), .S(n_64_2_8));
   HA_X1 i_64_2_4 (.A(SC[5]), .B(n_64_2_3), .CO(n_64_2_4), .S(n_64_2_9));
   NOR2_X1 i_64_2_5 (.A1(n_64_2_187), .A2(SC[0]), .ZN(n_64_194));
   AND2_X1 i_64_2_6 (.A1(n_64_2_5), .A2(n_64_2_181), .ZN(n_64_195));
   AND2_X1 i_64_2_7 (.A1(n_64_2_6), .A2(n_64_2_181), .ZN(n_64_196));
   AND2_X1 i_64_2_8 (.A1(n_64_2_7), .A2(n_64_2_181), .ZN(n_64_197));
   AND2_X1 i_64_2_9 (.A1(n_64_2_8), .A2(n_64_2_181), .ZN(n_64_198));
   AND2_X1 i_64_2_10 (.A1(n_64_2_9), .A2(n_64_2_181), .ZN(n_64_199));
   NOR2_X1 i_64_2_11 (.A1(n_64_362), .A2(n_64_2_10), .ZN(n_64_200));
   XNOR2_X1 i_64_2_12 (.A(SC[6]), .B(n_64_2_4), .ZN(n_64_2_10));
   AOI21_X1 i_64_2_13 (.A(n_64_2_13), .B1(n_64_2_11), .B2(en), .ZN(n_64_201));
   OAI21_X1 i_64_2_14 (.A(n_64_2_12), .B1(n_64_2_75), .B2(a[31]), .ZN(n_64_2_11));
   NAND2_X1 i_64_2_15 (.A1(b[31]), .A2(n_64_2_177), .ZN(n_64_2_12));
   AOI21_X1 i_64_2_16 (.A(out_sign), .B1(n_64_2_188), .B2(en), .ZN(n_64_2_13));
   OAI21_X1 i_64_2_17 (.A(n_64_2_14), .B1(n_64_2_44), .B2(n_64_2_46), .ZN(
      n_64_202));
   NAND2_X1 i_64_2_18 (.A1(n_64_2_44), .A2(n_64_130), .ZN(n_64_2_14));
   OAI21_X1 i_64_2_19 (.A(n_64_2_15), .B1(n_64_2_44), .B2(n_64_2_47), .ZN(
      n_64_203));
   NAND2_X1 i_64_2_20 (.A1(n_64_2_44), .A2(n_64_131), .ZN(n_64_2_15));
   OAI21_X1 i_64_2_21 (.A(n_64_2_16), .B1(n_64_2_44), .B2(n_64_2_48), .ZN(
      n_64_204));
   NAND2_X1 i_64_2_22 (.A1(n_64_2_44), .A2(n_64_132), .ZN(n_64_2_16));
   OAI21_X1 i_64_2_23 (.A(n_64_2_17), .B1(n_64_2_44), .B2(n_64_2_49), .ZN(
      n_64_205));
   NAND2_X1 i_64_2_24 (.A1(n_64_2_44), .A2(n_64_133), .ZN(n_64_2_17));
   OAI21_X1 i_64_2_25 (.A(n_64_2_18), .B1(n_64_2_44), .B2(n_64_2_50), .ZN(
      n_64_206));
   NAND2_X1 i_64_2_26 (.A1(n_64_2_44), .A2(n_64_134), .ZN(n_64_2_18));
   OAI21_X1 i_64_2_27 (.A(n_64_2_19), .B1(n_64_2_44), .B2(n_64_2_51), .ZN(
      n_64_207));
   NAND2_X1 i_64_2_28 (.A1(n_64_2_44), .A2(n_64_135), .ZN(n_64_2_19));
   OAI21_X1 i_64_2_29 (.A(n_64_2_20), .B1(n_64_2_44), .B2(n_64_2_52), .ZN(
      n_64_208));
   NAND2_X1 i_64_2_30 (.A1(n_64_2_44), .A2(n_64_136), .ZN(n_64_2_20));
   OAI21_X1 i_64_2_31 (.A(n_64_2_21), .B1(n_64_2_44), .B2(n_64_2_53), .ZN(
      n_64_209));
   NAND2_X1 i_64_2_32 (.A1(n_64_2_44), .A2(n_64_137), .ZN(n_64_2_21));
   OAI21_X1 i_64_2_33 (.A(n_64_2_22), .B1(n_64_2_44), .B2(n_64_2_54), .ZN(
      n_64_210));
   NAND2_X1 i_64_2_34 (.A1(n_64_2_44), .A2(n_64_138), .ZN(n_64_2_22));
   OAI21_X1 i_64_2_35 (.A(n_64_2_23), .B1(n_64_2_44), .B2(n_64_2_55), .ZN(
      n_64_211));
   NAND2_X1 i_64_2_36 (.A1(n_64_2_44), .A2(n_64_139), .ZN(n_64_2_23));
   OAI21_X1 i_64_2_37 (.A(n_64_2_24), .B1(n_64_2_44), .B2(n_64_2_56), .ZN(
      n_64_212));
   NAND2_X1 i_64_2_38 (.A1(n_64_2_44), .A2(n_64_140), .ZN(n_64_2_24));
   OAI21_X1 i_64_2_39 (.A(n_64_2_25), .B1(n_64_2_44), .B2(n_64_2_57), .ZN(
      n_64_213));
   NAND2_X1 i_64_2_40 (.A1(n_64_2_44), .A2(n_64_141), .ZN(n_64_2_25));
   OAI21_X1 i_64_2_41 (.A(n_64_2_26), .B1(n_64_2_44), .B2(n_64_2_58), .ZN(
      n_64_214));
   NAND2_X1 i_64_2_42 (.A1(n_64_2_44), .A2(n_64_142), .ZN(n_64_2_26));
   OAI21_X1 i_64_2_43 (.A(n_64_2_27), .B1(n_64_2_44), .B2(n_64_2_59), .ZN(
      n_64_215));
   NAND2_X1 i_64_2_44 (.A1(n_64_2_44), .A2(n_64_143), .ZN(n_64_2_27));
   OAI21_X1 i_64_2_45 (.A(n_64_2_28), .B1(n_64_2_44), .B2(n_64_2_60), .ZN(
      n_64_216));
   NAND2_X1 i_64_2_46 (.A1(n_64_2_44), .A2(n_64_144), .ZN(n_64_2_28));
   OAI21_X1 i_64_2_47 (.A(n_64_2_29), .B1(n_64_2_44), .B2(n_64_2_61), .ZN(
      n_64_217));
   NAND2_X1 i_64_2_48 (.A1(n_64_2_44), .A2(n_64_145), .ZN(n_64_2_29));
   OAI21_X1 i_64_2_49 (.A(n_64_2_30), .B1(n_64_2_44), .B2(n_64_2_62), .ZN(
      n_64_218));
   NAND2_X1 i_64_2_50 (.A1(n_64_2_44), .A2(n_64_146), .ZN(n_64_2_30));
   OAI21_X1 i_64_2_51 (.A(n_64_2_31), .B1(n_64_2_44), .B2(n_64_2_63), .ZN(
      n_64_219));
   NAND2_X1 i_64_2_52 (.A1(n_64_2_44), .A2(n_64_147), .ZN(n_64_2_31));
   OAI21_X1 i_64_2_53 (.A(n_64_2_32), .B1(n_64_2_44), .B2(n_64_2_64), .ZN(
      n_64_220));
   NAND2_X1 i_64_2_54 (.A1(n_64_2_44), .A2(n_64_148), .ZN(n_64_2_32));
   OAI21_X1 i_64_2_55 (.A(n_64_2_33), .B1(n_64_2_44), .B2(n_64_2_65), .ZN(
      n_64_221));
   NAND2_X1 i_64_2_56 (.A1(n_64_2_44), .A2(n_64_149), .ZN(n_64_2_33));
   OAI21_X1 i_64_2_57 (.A(n_64_2_34), .B1(n_64_2_44), .B2(n_64_2_66), .ZN(
      n_64_222));
   NAND2_X1 i_64_2_58 (.A1(n_64_2_44), .A2(n_64_150), .ZN(n_64_2_34));
   OAI21_X1 i_64_2_59 (.A(n_64_2_35), .B1(n_64_2_44), .B2(n_64_2_67), .ZN(
      n_64_223));
   NAND2_X1 i_64_2_60 (.A1(n_64_2_44), .A2(n_64_151), .ZN(n_64_2_35));
   OAI21_X1 i_64_2_61 (.A(n_64_2_36), .B1(n_64_2_44), .B2(n_64_2_68), .ZN(
      n_64_224));
   NAND2_X1 i_64_2_62 (.A1(n_64_2_44), .A2(n_64_152), .ZN(n_64_2_36));
   OAI21_X1 i_64_2_63 (.A(n_64_2_37), .B1(n_64_2_44), .B2(n_64_2_69), .ZN(
      n_64_225));
   NAND2_X1 i_64_2_64 (.A1(n_64_2_44), .A2(n_64_153), .ZN(n_64_2_37));
   OAI21_X1 i_64_2_65 (.A(n_64_2_38), .B1(n_64_2_44), .B2(n_64_2_70), .ZN(
      n_64_226));
   NAND2_X1 i_64_2_66 (.A1(n_64_2_44), .A2(n_64_154), .ZN(n_64_2_38));
   OAI21_X1 i_64_2_67 (.A(n_64_2_39), .B1(n_64_2_44), .B2(n_64_2_71), .ZN(
      n_64_227));
   NAND2_X1 i_64_2_68 (.A1(n_64_2_44), .A2(n_64_155), .ZN(n_64_2_39));
   OAI21_X1 i_64_2_69 (.A(n_64_2_40), .B1(n_64_2_44), .B2(n_64_2_72), .ZN(
      n_64_228));
   NAND2_X1 i_64_2_70 (.A1(n_64_2_44), .A2(n_64_156), .ZN(n_64_2_40));
   OAI21_X1 i_64_2_71 (.A(n_64_2_41), .B1(n_64_2_44), .B2(n_64_2_73), .ZN(
      n_64_229));
   NAND2_X1 i_64_2_72 (.A1(n_64_2_44), .A2(n_64_157), .ZN(n_64_2_41));
   OAI21_X1 i_64_2_73 (.A(n_64_2_42), .B1(n_64_2_44), .B2(n_64_2_74), .ZN(
      n_64_230));
   NAND2_X1 i_64_2_74 (.A1(n_64_2_44), .A2(n_64_158), .ZN(n_64_2_42));
   OAI21_X1 i_64_2_75 (.A(n_64_2_43), .B1(n_64_2_44), .B2(n_64_2_76), .ZN(
      n_64_231));
   NAND2_X1 i_64_2_76 (.A1(n_64_2_44), .A2(n_64_159), .ZN(n_64_2_43));
   MUX2_X1 i_64_2_77 (.A(n_64_298), .B(n_64_160), .S(n_64_2_44), .Z(n_64_232));
   MUX2_X1 i_64_2_78 (.A(n_64_299), .B(n_64_161), .S(n_64_2_44), .Z(n_64_233));
   MUX2_X1 i_64_2_79 (.A(n_64_300), .B(n_64_162), .S(n_64_2_44), .Z(n_64_234));
   MUX2_X1 i_64_2_80 (.A(n_64_301), .B(n_64_163), .S(n_64_2_44), .Z(n_64_235));
   MUX2_X1 i_64_2_81 (.A(n_64_302), .B(n_64_164), .S(n_64_2_44), .Z(n_64_236));
   MUX2_X1 i_64_2_82 (.A(n_64_303), .B(n_64_165), .S(n_64_2_44), .Z(n_64_237));
   MUX2_X1 i_64_2_83 (.A(n_64_304), .B(n_64_166), .S(n_64_2_44), .Z(n_64_238));
   MUX2_X1 i_64_2_84 (.A(n_64_305), .B(n_64_167), .S(n_64_2_44), .Z(n_64_239));
   MUX2_X1 i_64_2_85 (.A(n_64_306), .B(n_64_168), .S(n_64_2_44), .Z(n_64_240));
   MUX2_X1 i_64_2_86 (.A(n_64_307), .B(n_64_169), .S(n_64_2_44), .Z(n_64_241));
   MUX2_X1 i_64_2_87 (.A(n_64_308), .B(n_64_170), .S(n_64_2_44), .Z(n_64_242));
   MUX2_X1 i_64_2_88 (.A(n_64_309), .B(n_64_171), .S(n_64_2_44), .Z(n_64_243));
   MUX2_X1 i_64_2_89 (.A(n_64_310), .B(n_64_172), .S(n_64_2_44), .Z(n_64_244));
   MUX2_X1 i_64_2_90 (.A(n_64_311), .B(n_64_173), .S(n_64_2_44), .Z(n_64_245));
   MUX2_X1 i_64_2_91 (.A(n_64_312), .B(n_64_174), .S(n_64_2_44), .Z(n_64_246));
   MUX2_X1 i_64_2_92 (.A(n_64_313), .B(n_64_175), .S(n_64_2_44), .Z(n_64_247));
   MUX2_X1 i_64_2_93 (.A(n_64_314), .B(n_64_176), .S(n_64_2_44), .Z(n_64_248));
   MUX2_X1 i_64_2_94 (.A(n_64_315), .B(n_64_177), .S(n_64_2_44), .Z(n_64_249));
   MUX2_X1 i_64_2_95 (.A(n_64_316), .B(n_64_178), .S(n_64_2_44), .Z(n_64_250));
   MUX2_X1 i_64_2_96 (.A(n_64_317), .B(n_64_179), .S(n_64_2_44), .Z(n_64_251));
   MUX2_X1 i_64_2_97 (.A(n_64_318), .B(n_64_180), .S(n_64_2_44), .Z(n_64_252));
   MUX2_X1 i_64_2_98 (.A(n_64_319), .B(n_64_181), .S(n_64_2_44), .Z(n_64_253));
   MUX2_X1 i_64_2_99 (.A(n_64_320), .B(n_64_182), .S(n_64_2_44), .Z(n_64_254));
   MUX2_X1 i_64_2_100 (.A(n_64_321), .B(n_64_183), .S(n_64_2_44), .Z(n_64_255));
   MUX2_X1 i_64_2_101 (.A(n_64_322), .B(n_64_184), .S(n_64_2_44), .Z(n_64_256));
   MUX2_X1 i_64_2_102 (.A(n_64_323), .B(n_64_185), .S(n_64_2_44), .Z(n_64_257));
   MUX2_X1 i_64_2_103 (.A(n_64_324), .B(n_64_186), .S(n_64_2_44), .Z(n_64_258));
   MUX2_X1 i_64_2_104 (.A(n_64_325), .B(n_64_187), .S(n_64_2_44), .Z(n_64_259));
   MUX2_X1 i_64_2_105 (.A(n_64_326), .B(n_64_188), .S(n_64_2_44), .Z(n_64_260));
   MUX2_X1 i_64_2_106 (.A(n_64_327), .B(n_64_189), .S(n_64_2_44), .Z(n_64_261));
   MUX2_X1 i_64_2_107 (.A(n_64_328), .B(n_64_190), .S(n_64_2_44), .Z(n_64_262));
   MUX2_X1 i_64_2_108 (.A(n_64_329), .B(n_64_191), .S(n_64_2_44), .Z(n_64_263));
   AND2_X1 i_64_2_109 (.A1(n_64_2_44), .A2(n_64_192), .ZN(n_64_264));
   OR2_X1 i_64_2_110 (.A1(n_64_2_182), .A2(out_sign), .ZN(n_64_2_44));
   NOR2_X1 i_64_2_111 (.A1(n_64_2_187), .A2(rst), .ZN(n_64_265));
   INV_X1 i_64_2_112 (.A(n_64_2_45), .ZN(n_64_267));
   OAI222_X1 i_64_2_113 (.A1(n_64_2_75), .A2(b[1]), .B1(n_64_2_78), .B2(n_64_99), 
      .C1(Q[2]), .C2(n_64_2_188), .ZN(n_64_2_45));
   INV_X1 i_64_2_114 (.A(n_64_2_46), .ZN(n_64_268));
   OAI222_X1 i_64_2_115 (.A1(n_64_2_75), .A2(b[2]), .B1(n_64_2_78), .B2(n_64_100), 
      .C1(Q[3]), .C2(n_64_2_188), .ZN(n_64_2_46));
   INV_X1 i_64_2_116 (.A(n_64_2_47), .ZN(n_64_269));
   OAI222_X1 i_64_2_117 (.A1(n_64_2_75), .A2(b[3]), .B1(n_64_2_78), .B2(n_64_101), 
      .C1(Q[4]), .C2(n_64_2_188), .ZN(n_64_2_47));
   INV_X1 i_64_2_118 (.A(n_64_2_48), .ZN(n_64_270));
   OAI222_X1 i_64_2_119 (.A1(n_64_2_75), .A2(b[4]), .B1(n_64_2_78), .B2(n_64_102), 
      .C1(Q[5]), .C2(n_64_2_188), .ZN(n_64_2_48));
   INV_X1 i_64_2_120 (.A(n_64_2_49), .ZN(n_64_271));
   OAI222_X1 i_64_2_121 (.A1(n_64_2_75), .A2(b[5]), .B1(n_64_2_78), .B2(n_64_103), 
      .C1(Q[6]), .C2(n_64_2_188), .ZN(n_64_2_49));
   INV_X1 i_64_2_122 (.A(n_64_2_50), .ZN(n_64_272));
   OAI222_X1 i_64_2_123 (.A1(n_64_2_75), .A2(b[6]), .B1(n_64_2_78), .B2(n_64_104), 
      .C1(Q[7]), .C2(n_64_2_188), .ZN(n_64_2_50));
   INV_X1 i_64_2_124 (.A(n_64_2_51), .ZN(n_64_273));
   OAI222_X1 i_64_2_125 (.A1(n_64_2_75), .A2(b[7]), .B1(n_64_2_78), .B2(n_64_105), 
      .C1(Q[8]), .C2(n_64_2_188), .ZN(n_64_2_51));
   INV_X1 i_64_2_126 (.A(n_64_2_52), .ZN(n_64_274));
   OAI222_X1 i_64_2_127 (.A1(n_64_2_75), .A2(b[8]), .B1(n_64_2_78), .B2(n_64_106), 
      .C1(Q[9]), .C2(n_64_2_188), .ZN(n_64_2_52));
   INV_X1 i_64_2_128 (.A(n_64_2_53), .ZN(n_64_275));
   OAI222_X1 i_64_2_129 (.A1(n_64_2_75), .A2(b[9]), .B1(n_64_2_78), .B2(n_64_107), 
      .C1(Q[10]), .C2(n_64_2_188), .ZN(n_64_2_53));
   INV_X1 i_64_2_130 (.A(n_64_2_54), .ZN(n_64_276));
   OAI222_X1 i_64_2_131 (.A1(n_64_2_75), .A2(b[10]), .B1(n_64_2_78), .B2(
      n_64_108), .C1(Q[11]), .C2(n_64_2_188), .ZN(n_64_2_54));
   INV_X1 i_64_2_132 (.A(n_64_2_55), .ZN(n_64_277));
   OAI222_X1 i_64_2_133 (.A1(n_64_2_75), .A2(b[11]), .B1(n_64_2_78), .B2(
      n_64_109), .C1(Q[12]), .C2(n_64_2_188), .ZN(n_64_2_55));
   INV_X1 i_64_2_134 (.A(n_64_2_56), .ZN(n_64_278));
   OAI222_X1 i_64_2_135 (.A1(n_64_2_75), .A2(b[12]), .B1(n_64_2_78), .B2(
      n_64_110), .C1(Q[13]), .C2(n_64_2_188), .ZN(n_64_2_56));
   INV_X1 i_64_2_136 (.A(n_64_2_57), .ZN(n_64_279));
   OAI222_X1 i_64_2_137 (.A1(n_64_2_75), .A2(b[13]), .B1(n_64_2_78), .B2(
      n_64_111), .C1(Q[14]), .C2(n_64_2_188), .ZN(n_64_2_57));
   INV_X1 i_64_2_138 (.A(n_64_2_58), .ZN(n_64_280));
   OAI222_X1 i_64_2_139 (.A1(n_64_2_75), .A2(b[14]), .B1(n_64_2_78), .B2(
      n_64_112), .C1(Q[15]), .C2(n_64_2_188), .ZN(n_64_2_58));
   INV_X1 i_64_2_140 (.A(n_64_2_59), .ZN(n_64_281));
   OAI222_X1 i_64_2_141 (.A1(n_64_2_75), .A2(b[15]), .B1(n_64_2_78), .B2(
      n_64_113), .C1(Q[16]), .C2(n_64_2_188), .ZN(n_64_2_59));
   INV_X1 i_64_2_142 (.A(n_64_2_60), .ZN(n_64_282));
   OAI222_X1 i_64_2_143 (.A1(n_64_2_75), .A2(b[16]), .B1(n_64_2_78), .B2(
      n_64_114), .C1(Q[17]), .C2(n_64_2_188), .ZN(n_64_2_60));
   INV_X1 i_64_2_144 (.A(n_64_2_61), .ZN(n_64_283));
   OAI222_X1 i_64_2_145 (.A1(n_64_2_75), .A2(b[17]), .B1(n_64_2_78), .B2(
      n_64_115), .C1(Q[18]), .C2(n_64_2_188), .ZN(n_64_2_61));
   INV_X1 i_64_2_146 (.A(n_64_2_62), .ZN(n_64_284));
   OAI222_X1 i_64_2_147 (.A1(n_64_2_75), .A2(b[18]), .B1(n_64_2_78), .B2(
      n_64_116), .C1(Q[19]), .C2(n_64_2_188), .ZN(n_64_2_62));
   INV_X1 i_64_2_148 (.A(n_64_2_63), .ZN(n_64_285));
   OAI222_X1 i_64_2_149 (.A1(n_64_2_75), .A2(b[19]), .B1(n_64_2_78), .B2(
      n_64_117), .C1(Q[20]), .C2(n_64_2_188), .ZN(n_64_2_63));
   INV_X1 i_64_2_150 (.A(n_64_2_64), .ZN(n_64_286));
   OAI222_X1 i_64_2_151 (.A1(n_64_2_75), .A2(b[20]), .B1(n_64_2_78), .B2(
      n_64_118), .C1(Q[21]), .C2(n_64_2_188), .ZN(n_64_2_64));
   INV_X1 i_64_2_152 (.A(n_64_2_65), .ZN(n_64_287));
   OAI222_X1 i_64_2_153 (.A1(n_64_2_75), .A2(b[21]), .B1(n_64_2_78), .B2(
      n_64_119), .C1(Q[22]), .C2(n_64_2_188), .ZN(n_64_2_65));
   INV_X1 i_64_2_154 (.A(n_64_2_66), .ZN(n_64_288));
   OAI222_X1 i_64_2_155 (.A1(n_64_2_75), .A2(b[22]), .B1(n_64_2_78), .B2(
      n_64_120), .C1(Q[23]), .C2(n_64_2_188), .ZN(n_64_2_66));
   INV_X1 i_64_2_156 (.A(n_64_2_67), .ZN(n_64_289));
   OAI222_X1 i_64_2_157 (.A1(n_64_2_75), .A2(b[23]), .B1(n_64_2_78), .B2(
      n_64_121), .C1(Q[24]), .C2(n_64_2_188), .ZN(n_64_2_67));
   INV_X1 i_64_2_158 (.A(n_64_2_68), .ZN(n_64_290));
   OAI222_X1 i_64_2_159 (.A1(n_64_2_75), .A2(b[24]), .B1(n_64_2_78), .B2(
      n_64_122), .C1(Q[25]), .C2(n_64_2_188), .ZN(n_64_2_68));
   INV_X1 i_64_2_160 (.A(n_64_2_69), .ZN(n_64_291));
   OAI222_X1 i_64_2_161 (.A1(n_64_2_75), .A2(b[25]), .B1(n_64_2_78), .B2(
      n_64_123), .C1(Q[26]), .C2(n_64_2_188), .ZN(n_64_2_69));
   INV_X1 i_64_2_162 (.A(n_64_2_70), .ZN(n_64_292));
   OAI222_X1 i_64_2_163 (.A1(n_64_2_75), .A2(b[26]), .B1(n_64_2_78), .B2(
      n_64_124), .C1(Q[27]), .C2(n_64_2_188), .ZN(n_64_2_70));
   INV_X1 i_64_2_164 (.A(n_64_2_71), .ZN(n_64_293));
   OAI222_X1 i_64_2_165 (.A1(n_64_2_75), .A2(b[27]), .B1(n_64_2_78), .B2(
      n_64_125), .C1(Q[28]), .C2(n_64_2_188), .ZN(n_64_2_71));
   INV_X1 i_64_2_166 (.A(n_64_2_72), .ZN(n_64_294));
   OAI222_X1 i_64_2_167 (.A1(n_64_2_75), .A2(b[28]), .B1(n_64_2_78), .B2(
      n_64_126), .C1(Q[29]), .C2(n_64_2_188), .ZN(n_64_2_72));
   INV_X1 i_64_2_168 (.A(n_64_2_73), .ZN(n_64_295));
   OAI222_X1 i_64_2_169 (.A1(n_64_2_75), .A2(b[29]), .B1(n_64_2_78), .B2(
      n_64_127), .C1(Q[30]), .C2(n_64_2_188), .ZN(n_64_2_73));
   INV_X1 i_64_2_170 (.A(n_64_2_74), .ZN(n_64_296));
   OAI222_X1 i_64_2_171 (.A1(n_64_2_75), .A2(b[30]), .B1(n_64_2_78), .B2(
      n_64_128), .C1(Q[31]), .C2(n_64_2_188), .ZN(n_64_2_74));
   OR2_X1 i_64_2_172 (.A1(n_64_2_178), .A2(b[31]), .ZN(n_64_2_75));
   INV_X1 i_64_2_173 (.A(n_64_2_76), .ZN(n_64_297));
   AOI22_X1 i_64_2_174 (.A1(n_64_129), .A2(n_64_2_77), .B1(n_64_2_178), .B2(
      Q[32]), .ZN(n_64_2_76));
   INV_X1 i_64_2_175 (.A(n_64_2_78), .ZN(n_64_2_77));
   NAND2_X1 i_64_2_176 (.A1(b[31]), .A2(n_64_2_188), .ZN(n_64_2_78));
   NOR2_X1 i_64_2_177 (.A1(n_64_2_80), .A2(n_64_2_79), .ZN(n_64_298));
   OAI22_X1 i_64_2_178 (.A1(n_64_35), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_67), .ZN(n_64_2_79));
   NOR2_X1 i_64_2_179 (.A1(n_64_2_142), .A2(A[0]), .ZN(n_64_2_80));
   NOR2_X1 i_64_2_180 (.A1(n_64_2_82), .A2(n_64_2_81), .ZN(n_64_299));
   OAI22_X1 i_64_2_181 (.A1(n_64_36), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_68), .ZN(n_64_2_81));
   NOR2_X1 i_64_2_182 (.A1(n_64_2_142), .A2(A[1]), .ZN(n_64_2_82));
   NOR2_X1 i_64_2_183 (.A1(n_64_2_84), .A2(n_64_2_83), .ZN(n_64_300));
   OAI22_X1 i_64_2_184 (.A1(n_64_37), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_69), .ZN(n_64_2_83));
   NOR2_X1 i_64_2_185 (.A1(n_64_2_142), .A2(A[2]), .ZN(n_64_2_84));
   NOR2_X1 i_64_2_186 (.A1(n_64_2_86), .A2(n_64_2_85), .ZN(n_64_301));
   OAI22_X1 i_64_2_187 (.A1(n_64_38), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_70), .ZN(n_64_2_85));
   NOR2_X1 i_64_2_188 (.A1(n_64_2_142), .A2(A[3]), .ZN(n_64_2_86));
   NOR2_X1 i_64_2_189 (.A1(n_64_2_88), .A2(n_64_2_87), .ZN(n_64_302));
   OAI22_X1 i_64_2_190 (.A1(n_64_39), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_71), .ZN(n_64_2_87));
   NOR2_X1 i_64_2_191 (.A1(n_64_2_142), .A2(A[4]), .ZN(n_64_2_88));
   NOR2_X1 i_64_2_192 (.A1(n_64_2_90), .A2(n_64_2_89), .ZN(n_64_303));
   OAI22_X1 i_64_2_193 (.A1(n_64_40), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_72), .ZN(n_64_2_89));
   NOR2_X1 i_64_2_194 (.A1(n_64_2_142), .A2(A[5]), .ZN(n_64_2_90));
   NOR2_X1 i_64_2_195 (.A1(n_64_2_92), .A2(n_64_2_91), .ZN(n_64_304));
   OAI22_X1 i_64_2_196 (.A1(n_64_41), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_73), .ZN(n_64_2_91));
   NOR2_X1 i_64_2_197 (.A1(n_64_2_142), .A2(A[6]), .ZN(n_64_2_92));
   NOR2_X1 i_64_2_198 (.A1(n_64_2_94), .A2(n_64_2_93), .ZN(n_64_305));
   OAI22_X1 i_64_2_199 (.A1(n_64_42), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_74), .ZN(n_64_2_93));
   NOR2_X1 i_64_2_200 (.A1(n_64_2_142), .A2(A[7]), .ZN(n_64_2_94));
   NOR2_X1 i_64_2_201 (.A1(n_64_2_96), .A2(n_64_2_95), .ZN(n_64_306));
   OAI22_X1 i_64_2_202 (.A1(n_64_43), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_75), .ZN(n_64_2_95));
   NOR2_X1 i_64_2_203 (.A1(n_64_2_142), .A2(A[8]), .ZN(n_64_2_96));
   NOR2_X1 i_64_2_204 (.A1(n_64_2_98), .A2(n_64_2_97), .ZN(n_64_307));
   OAI22_X1 i_64_2_205 (.A1(n_64_44), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_76), .ZN(n_64_2_97));
   NOR2_X1 i_64_2_206 (.A1(n_64_2_142), .A2(A[9]), .ZN(n_64_2_98));
   NOR2_X1 i_64_2_207 (.A1(n_64_2_100), .A2(n_64_2_99), .ZN(n_64_308));
   OAI22_X1 i_64_2_208 (.A1(n_64_45), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_77), .ZN(n_64_2_99));
   NOR2_X1 i_64_2_209 (.A1(n_64_2_142), .A2(A[10]), .ZN(n_64_2_100));
   NOR2_X1 i_64_2_210 (.A1(n_64_2_102), .A2(n_64_2_101), .ZN(n_64_309));
   OAI22_X1 i_64_2_211 (.A1(n_64_46), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_78), .ZN(n_64_2_101));
   NOR2_X1 i_64_2_212 (.A1(n_64_2_142), .A2(A[11]), .ZN(n_64_2_102));
   NOR2_X1 i_64_2_213 (.A1(n_64_2_104), .A2(n_64_2_103), .ZN(n_64_310));
   OAI22_X1 i_64_2_214 (.A1(n_64_47), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_79), .ZN(n_64_2_103));
   NOR2_X1 i_64_2_215 (.A1(n_64_2_142), .A2(A[12]), .ZN(n_64_2_104));
   NOR2_X1 i_64_2_216 (.A1(n_64_2_106), .A2(n_64_2_105), .ZN(n_64_311));
   OAI22_X1 i_64_2_217 (.A1(n_64_48), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_80), .ZN(n_64_2_105));
   NOR2_X1 i_64_2_218 (.A1(n_64_2_142), .A2(A[13]), .ZN(n_64_2_106));
   NOR2_X1 i_64_2_219 (.A1(n_64_2_108), .A2(n_64_2_107), .ZN(n_64_312));
   OAI22_X1 i_64_2_220 (.A1(n_64_49), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_81), .ZN(n_64_2_107));
   NOR2_X1 i_64_2_221 (.A1(n_64_2_142), .A2(A[14]), .ZN(n_64_2_108));
   NOR2_X1 i_64_2_222 (.A1(n_64_2_110), .A2(n_64_2_109), .ZN(n_64_313));
   OAI22_X1 i_64_2_223 (.A1(n_64_50), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_82), .ZN(n_64_2_109));
   NOR2_X1 i_64_2_224 (.A1(n_64_2_142), .A2(A[15]), .ZN(n_64_2_110));
   NOR2_X1 i_64_2_225 (.A1(n_64_2_112), .A2(n_64_2_111), .ZN(n_64_314));
   OAI22_X1 i_64_2_226 (.A1(n_64_51), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_83), .ZN(n_64_2_111));
   NOR2_X1 i_64_2_227 (.A1(n_64_2_142), .A2(A[16]), .ZN(n_64_2_112));
   NOR2_X1 i_64_2_228 (.A1(n_64_2_114), .A2(n_64_2_113), .ZN(n_64_315));
   OAI22_X1 i_64_2_229 (.A1(n_64_52), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_84), .ZN(n_64_2_113));
   NOR2_X1 i_64_2_230 (.A1(n_64_2_142), .A2(A[17]), .ZN(n_64_2_114));
   NOR2_X1 i_64_2_231 (.A1(n_64_2_116), .A2(n_64_2_115), .ZN(n_64_316));
   OAI22_X1 i_64_2_232 (.A1(n_64_53), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_85), .ZN(n_64_2_115));
   NOR2_X1 i_64_2_233 (.A1(n_64_2_142), .A2(A[18]), .ZN(n_64_2_116));
   NOR2_X1 i_64_2_234 (.A1(n_64_2_118), .A2(n_64_2_117), .ZN(n_64_317));
   OAI22_X1 i_64_2_235 (.A1(n_64_54), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_86), .ZN(n_64_2_117));
   NOR2_X1 i_64_2_236 (.A1(n_64_2_142), .A2(A[19]), .ZN(n_64_2_118));
   NOR2_X1 i_64_2_237 (.A1(n_64_2_120), .A2(n_64_2_119), .ZN(n_64_318));
   OAI22_X1 i_64_2_238 (.A1(n_64_55), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_87), .ZN(n_64_2_119));
   NOR2_X1 i_64_2_239 (.A1(n_64_2_142), .A2(A[20]), .ZN(n_64_2_120));
   NOR2_X1 i_64_2_240 (.A1(n_64_2_122), .A2(n_64_2_121), .ZN(n_64_319));
   OAI22_X1 i_64_2_241 (.A1(n_64_56), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_88), .ZN(n_64_2_121));
   NOR2_X1 i_64_2_242 (.A1(n_64_2_142), .A2(A[21]), .ZN(n_64_2_122));
   NOR2_X1 i_64_2_243 (.A1(n_64_2_124), .A2(n_64_2_123), .ZN(n_64_320));
   OAI22_X1 i_64_2_244 (.A1(n_64_57), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_89), .ZN(n_64_2_123));
   NOR2_X1 i_64_2_245 (.A1(n_64_2_142), .A2(A[22]), .ZN(n_64_2_124));
   NOR2_X1 i_64_2_246 (.A1(n_64_2_126), .A2(n_64_2_125), .ZN(n_64_321));
   OAI22_X1 i_64_2_247 (.A1(n_64_58), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_90), .ZN(n_64_2_125));
   NOR2_X1 i_64_2_248 (.A1(n_64_2_142), .A2(A[23]), .ZN(n_64_2_126));
   NOR2_X1 i_64_2_249 (.A1(n_64_2_128), .A2(n_64_2_127), .ZN(n_64_322));
   OAI22_X1 i_64_2_250 (.A1(n_64_59), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_91), .ZN(n_64_2_127));
   NOR2_X1 i_64_2_251 (.A1(n_64_2_142), .A2(A[24]), .ZN(n_64_2_128));
   NOR2_X1 i_64_2_252 (.A1(n_64_2_130), .A2(n_64_2_129), .ZN(n_64_323));
   OAI22_X1 i_64_2_253 (.A1(n_64_60), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_92), .ZN(n_64_2_129));
   NOR2_X1 i_64_2_254 (.A1(n_64_2_142), .A2(A[25]), .ZN(n_64_2_130));
   NOR2_X1 i_64_2_255 (.A1(n_64_2_132), .A2(n_64_2_131), .ZN(n_64_324));
   OAI22_X1 i_64_2_256 (.A1(n_64_61), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_93), .ZN(n_64_2_131));
   NOR2_X1 i_64_2_257 (.A1(n_64_2_142), .A2(A[26]), .ZN(n_64_2_132));
   NOR2_X1 i_64_2_258 (.A1(n_64_2_134), .A2(n_64_2_133), .ZN(n_64_325));
   OAI22_X1 i_64_2_259 (.A1(n_64_62), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_94), .ZN(n_64_2_133));
   NOR2_X1 i_64_2_260 (.A1(n_64_2_142), .A2(A[27]), .ZN(n_64_2_134));
   NOR2_X1 i_64_2_261 (.A1(n_64_2_136), .A2(n_64_2_135), .ZN(n_64_326));
   OAI22_X1 i_64_2_262 (.A1(n_64_63), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_95), .ZN(n_64_2_135));
   NOR2_X1 i_64_2_263 (.A1(n_64_2_142), .A2(A[28]), .ZN(n_64_2_136));
   NOR2_X1 i_64_2_264 (.A1(n_64_2_138), .A2(n_64_2_137), .ZN(n_64_327));
   OAI22_X1 i_64_2_265 (.A1(n_64_64), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_96), .ZN(n_64_2_137));
   NOR2_X1 i_64_2_266 (.A1(n_64_2_142), .A2(A[29]), .ZN(n_64_2_138));
   NOR2_X1 i_64_2_267 (.A1(n_64_2_141), .A2(n_64_2_139), .ZN(n_64_328));
   OAI22_X1 i_64_2_268 (.A1(n_64_65), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_97), .ZN(n_64_2_139));
   NOR2_X1 i_64_2_269 (.A1(n_64_2_141), .A2(n_64_2_140), .ZN(n_64_329));
   OAI22_X1 i_64_2_270 (.A1(n_64_66), .A2(n_64_2_144), .B1(n_64_2_143), .B2(
      n_64_98), .ZN(n_64_2_140));
   NOR2_X1 i_64_2_271 (.A1(n_64_2_142), .A2(A[31]), .ZN(n_64_2_141));
   NAND2_X1 i_64_2_272 (.A1(n_64_2_144), .A2(n_64_2_143), .ZN(n_64_2_142));
   OR3_X1 i_64_2_273 (.A1(Q[1]), .A2(n_64_2_188), .A3(n_64_2_185), .ZN(
      n_64_2_143));
   OAI21_X1 i_64_2_274 (.A(n_64_266), .B1(n_64_2_188), .B2(n_64_2_185), .ZN(
      n_64_2_144));
   MUX2_X1 i_64_2_275 (.A(b[0]), .B(Q[1]), .S(n_64_2_178), .Z(n_64_266));
   MUX2_X1 i_64_2_276 (.A(a[0]), .B(multiplicand[0]), .S(n_64_2_178), .Z(
      n_64_330));
   INV_X1 i_64_2_277 (.A(n_64_2_145), .ZN(n_64_331));
   AOI222_X1 i_64_2_278 (.A1(n_64_4), .A2(n_64_2_177), .B1(n_64_2_175), .B2(a[1]), 
      .C1(n_64_2_178), .C2(multiplicand[1]), .ZN(n_64_2_145));
   INV_X1 i_64_2_279 (.A(n_64_2_146), .ZN(n_64_332));
   AOI222_X1 i_64_2_280 (.A1(n_64_5), .A2(n_64_2_177), .B1(n_64_2_175), .B2(a[2]), 
      .C1(n_64_2_178), .C2(multiplicand[2]), .ZN(n_64_2_146));
   INV_X1 i_64_2_281 (.A(n_64_2_147), .ZN(n_64_333));
   AOI222_X1 i_64_2_282 (.A1(n_64_6), .A2(n_64_2_177), .B1(n_64_2_175), .B2(a[3]), 
      .C1(n_64_2_178), .C2(multiplicand[3]), .ZN(n_64_2_147));
   INV_X1 i_64_2_283 (.A(n_64_2_148), .ZN(n_64_334));
   AOI222_X1 i_64_2_284 (.A1(n_64_7), .A2(n_64_2_177), .B1(n_64_2_175), .B2(a[4]), 
      .C1(n_64_2_178), .C2(multiplicand[4]), .ZN(n_64_2_148));
   INV_X1 i_64_2_285 (.A(n_64_2_149), .ZN(n_64_335));
   AOI222_X1 i_64_2_286 (.A1(n_64_8), .A2(n_64_2_177), .B1(n_64_2_175), .B2(a[5]), 
      .C1(n_64_2_178), .C2(multiplicand[5]), .ZN(n_64_2_149));
   INV_X1 i_64_2_287 (.A(n_64_2_150), .ZN(n_64_336));
   AOI222_X1 i_64_2_288 (.A1(n_64_9), .A2(n_64_2_177), .B1(n_64_2_175), .B2(a[6]), 
      .C1(n_64_2_178), .C2(multiplicand[6]), .ZN(n_64_2_150));
   INV_X1 i_64_2_289 (.A(n_64_2_151), .ZN(n_64_337));
   AOI222_X1 i_64_2_290 (.A1(n_64_10), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[7]), .C1(n_64_2_178), .C2(multiplicand[7]), .ZN(n_64_2_151));
   INV_X1 i_64_2_291 (.A(n_64_2_152), .ZN(n_64_338));
   AOI222_X1 i_64_2_292 (.A1(n_64_11), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[8]), .C1(n_64_2_178), .C2(multiplicand[8]), .ZN(n_64_2_152));
   INV_X1 i_64_2_293 (.A(n_64_2_153), .ZN(n_64_339));
   AOI222_X1 i_64_2_294 (.A1(n_64_12), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[9]), .C1(n_64_2_178), .C2(multiplicand[9]), .ZN(n_64_2_153));
   INV_X1 i_64_2_295 (.A(n_64_2_154), .ZN(n_64_340));
   AOI222_X1 i_64_2_296 (.A1(n_64_13), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[10]), .C1(n_64_2_178), .C2(multiplicand[10]), .ZN(n_64_2_154));
   INV_X1 i_64_2_297 (.A(n_64_2_155), .ZN(n_64_341));
   AOI222_X1 i_64_2_298 (.A1(n_64_14), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[11]), .C1(n_64_2_178), .C2(multiplicand[11]), .ZN(n_64_2_155));
   INV_X1 i_64_2_299 (.A(n_64_2_156), .ZN(n_64_342));
   AOI222_X1 i_64_2_300 (.A1(n_64_15), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[12]), .C1(n_64_2_178), .C2(multiplicand[12]), .ZN(n_64_2_156));
   INV_X1 i_64_2_301 (.A(n_64_2_157), .ZN(n_64_343));
   AOI222_X1 i_64_2_302 (.A1(n_64_16), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[13]), .C1(n_64_2_178), .C2(multiplicand[13]), .ZN(n_64_2_157));
   INV_X1 i_64_2_303 (.A(n_64_2_158), .ZN(n_64_344));
   AOI222_X1 i_64_2_304 (.A1(n_64_17), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[14]), .C1(n_64_2_178), .C2(multiplicand[14]), .ZN(n_64_2_158));
   INV_X1 i_64_2_305 (.A(n_64_2_159), .ZN(n_64_345));
   AOI222_X1 i_64_2_306 (.A1(n_64_18), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[15]), .C1(n_64_2_178), .C2(multiplicand[15]), .ZN(n_64_2_159));
   INV_X1 i_64_2_307 (.A(n_64_2_160), .ZN(n_64_346));
   AOI222_X1 i_64_2_308 (.A1(n_64_19), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[16]), .C1(n_64_2_178), .C2(multiplicand[16]), .ZN(n_64_2_160));
   INV_X1 i_64_2_309 (.A(n_64_2_161), .ZN(n_64_347));
   AOI222_X1 i_64_2_310 (.A1(n_64_20), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[17]), .C1(n_64_2_178), .C2(multiplicand[17]), .ZN(n_64_2_161));
   INV_X1 i_64_2_311 (.A(n_64_2_162), .ZN(n_64_348));
   AOI222_X1 i_64_2_312 (.A1(n_64_21), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[18]), .C1(n_64_2_178), .C2(multiplicand[18]), .ZN(n_64_2_162));
   INV_X1 i_64_2_313 (.A(n_64_2_163), .ZN(n_64_349));
   AOI222_X1 i_64_2_314 (.A1(n_64_22), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[19]), .C1(n_64_2_178), .C2(multiplicand[19]), .ZN(n_64_2_163));
   INV_X1 i_64_2_315 (.A(n_64_2_164), .ZN(n_64_350));
   AOI222_X1 i_64_2_316 (.A1(n_64_23), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[20]), .C1(n_64_2_178), .C2(multiplicand[20]), .ZN(n_64_2_164));
   INV_X1 i_64_2_317 (.A(n_64_2_165), .ZN(n_64_351));
   AOI222_X1 i_64_2_318 (.A1(n_64_24), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[21]), .C1(n_64_2_178), .C2(multiplicand[21]), .ZN(n_64_2_165));
   INV_X1 i_64_2_319 (.A(n_64_2_166), .ZN(n_64_352));
   AOI222_X1 i_64_2_320 (.A1(n_64_25), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[22]), .C1(n_64_2_178), .C2(multiplicand[22]), .ZN(n_64_2_166));
   INV_X1 i_64_2_321 (.A(n_64_2_167), .ZN(n_64_353));
   AOI222_X1 i_64_2_322 (.A1(n_64_26), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[23]), .C1(n_64_2_178), .C2(multiplicand[23]), .ZN(n_64_2_167));
   INV_X1 i_64_2_323 (.A(n_64_2_168), .ZN(n_64_354));
   AOI222_X1 i_64_2_324 (.A1(n_64_27), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[24]), .C1(n_64_2_178), .C2(multiplicand[24]), .ZN(n_64_2_168));
   INV_X1 i_64_2_325 (.A(n_64_2_169), .ZN(n_64_355));
   AOI222_X1 i_64_2_326 (.A1(n_64_28), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[25]), .C1(n_64_2_178), .C2(multiplicand[25]), .ZN(n_64_2_169));
   INV_X1 i_64_2_327 (.A(n_64_2_170), .ZN(n_64_356));
   AOI222_X1 i_64_2_328 (.A1(n_64_29), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[26]), .C1(n_64_2_178), .C2(multiplicand[26]), .ZN(n_64_2_170));
   INV_X1 i_64_2_329 (.A(n_64_2_171), .ZN(n_64_357));
   AOI222_X1 i_64_2_330 (.A1(n_64_30), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[27]), .C1(n_64_2_178), .C2(multiplicand[27]), .ZN(n_64_2_171));
   INV_X1 i_64_2_331 (.A(n_64_2_172), .ZN(n_64_358));
   AOI222_X1 i_64_2_332 (.A1(n_64_31), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[28]), .C1(n_64_2_178), .C2(multiplicand[28]), .ZN(n_64_2_172));
   INV_X1 i_64_2_333 (.A(n_64_2_173), .ZN(n_64_359));
   AOI222_X1 i_64_2_334 (.A1(n_64_32), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[29]), .C1(n_64_2_178), .C2(multiplicand[29]), .ZN(n_64_2_173));
   INV_X1 i_64_2_335 (.A(n_64_2_174), .ZN(n_64_360));
   AOI222_X1 i_64_2_336 (.A1(n_64_33), .A2(n_64_2_177), .B1(n_64_2_175), 
      .B2(a[30]), .C1(n_64_2_178), .C2(multiplicand[30]), .ZN(n_64_2_174));
   NOR2_X1 i_64_2_337 (.A1(n_64_2_178), .A2(a[31]), .ZN(n_64_2_175));
   INV_X1 i_64_2_338 (.A(n_64_2_176), .ZN(n_64_361));
   AOI22_X1 i_64_2_339 (.A1(n_64_34), .A2(n_64_2_177), .B1(n_64_2_178), .B2(
      multiplicand[31]), .ZN(n_64_2_176));
   AND2_X1 i_64_2_340 (.A1(a[31]), .A2(n_64_2_188), .ZN(n_64_2_177));
   NAND3_X1 i_64_2_341 (.A1(n_64_2_183), .A2(n_64_2_180), .A3(n_64_2_179), 
      .ZN(n_64_2_178));
   NOR2_X1 i_64_2_342 (.A1(SC[4]), .A2(SC[3]), .ZN(n_64_2_179));
   NOR3_X1 i_64_2_343 (.A1(SC[2]), .A2(SC[1]), .A3(SC[0]), .ZN(n_64_2_180));
   INV_X1 i_64_2_344 (.A(n_64_2_181), .ZN(n_64_362));
   AND2_X1 i_64_2_345 (.A1(n_64_2_182), .A2(en), .ZN(n_64_2_181));
   AOI21_X1 i_64_2_346 (.A(n_64_2_187), .B1(n_64_2_186), .B2(n_64_2_182), 
      .ZN(n_64_363));
   NAND4_X1 i_64_2_347 (.A1(SC[4]), .A2(SC[3]), .A3(n_64_2_184), .A4(n_64_2_183), 
      .ZN(n_64_2_182));
   NOR2_X1 i_64_2_348 (.A1(SC[6]), .A2(SC[5]), .ZN(n_64_2_183));
   AND3_X1 i_64_2_349 (.A1(SC[2]), .A2(SC[1]), .A3(SC[0]), .ZN(n_64_2_184));
   INV_X1 i_64_2_350 (.A(Q[0]), .ZN(n_64_2_185));
   INV_X1 i_64_2_351 (.A(n_64_3), .ZN(n_64_2_186));
   INV_X1 i_64_2_352 (.A(en), .ZN(n_64_2_187));
   INV_X1 i_64_2_353 (.A(n_64_2_178), .ZN(n_64_2_188));
endmodule
