
// 	Thu Dec 22 23:27:55 2022
//	vlsi
//	localhost.localdomain

module buffer__parameterized0 (clk_CTS_0_PP_0, clk, rst, en, D, Q);

output [63:0] Q;
input [63:0] D;
input clk;
input en;
input rst;
input clk_CTS_0_PP_0;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_8;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire hfn_ipo_n5;
wire hfn_ipo_n6;
wire CTS_n_tid1_9;


AND2_X1 i_0_65 (.ZN (n_65), .A1 (hfn_ipo_n6), .A2 (D[63]));
AND2_X1 i_0_64 (.ZN (n_64), .A1 (hfn_ipo_n6), .A2 (D[62]));
AND2_X1 i_0_63 (.ZN (n_63), .A1 (hfn_ipo_n6), .A2 (D[61]));
AND2_X1 i_0_62 (.ZN (n_62), .A1 (hfn_ipo_n6), .A2 (D[60]));
AND2_X1 i_0_61 (.ZN (n_61), .A1 (hfn_ipo_n6), .A2 (D[59]));
AND2_X1 i_0_60 (.ZN (n_60), .A1 (hfn_ipo_n6), .A2 (D[58]));
AND2_X1 i_0_59 (.ZN (n_59), .A1 (hfn_ipo_n6), .A2 (D[57]));
AND2_X1 i_0_58 (.ZN (n_58), .A1 (hfn_ipo_n6), .A2 (D[56]));
AND2_X1 i_0_57 (.ZN (n_57), .A1 (hfn_ipo_n6), .A2 (D[55]));
AND2_X1 i_0_56 (.ZN (n_56), .A1 (hfn_ipo_n6), .A2 (D[54]));
AND2_X1 i_0_55 (.ZN (n_55), .A1 (hfn_ipo_n6), .A2 (D[53]));
AND2_X1 i_0_54 (.ZN (n_54), .A1 (hfn_ipo_n6), .A2 (D[52]));
AND2_X1 i_0_53 (.ZN (n_53), .A1 (hfn_ipo_n6), .A2 (D[51]));
AND2_X1 i_0_52 (.ZN (n_52), .A1 (hfn_ipo_n6), .A2 (D[50]));
AND2_X1 i_0_51 (.ZN (n_51), .A1 (hfn_ipo_n6), .A2 (D[49]));
AND2_X1 i_0_50 (.ZN (n_50), .A1 (hfn_ipo_n5), .A2 (D[48]));
AND2_X1 i_0_49 (.ZN (n_49), .A1 (hfn_ipo_n5), .A2 (D[47]));
AND2_X1 i_0_48 (.ZN (n_48), .A1 (hfn_ipo_n5), .A2 (D[46]));
AND2_X1 i_0_47 (.ZN (n_47), .A1 (hfn_ipo_n5), .A2 (D[45]));
AND2_X1 i_0_46 (.ZN (n_46), .A1 (hfn_ipo_n5), .A2 (D[44]));
AND2_X1 i_0_45 (.ZN (n_45), .A1 (hfn_ipo_n5), .A2 (D[43]));
AND2_X1 i_0_44 (.ZN (n_44), .A1 (hfn_ipo_n5), .A2 (D[42]));
AND2_X1 i_0_43 (.ZN (n_43), .A1 (hfn_ipo_n5), .A2 (D[41]));
AND2_X1 i_0_42 (.ZN (n_42), .A1 (hfn_ipo_n5), .A2 (D[40]));
AND2_X1 i_0_41 (.ZN (n_41), .A1 (hfn_ipo_n5), .A2 (D[39]));
AND2_X1 i_0_40 (.ZN (n_40), .A1 (hfn_ipo_n5), .A2 (D[38]));
AND2_X1 i_0_39 (.ZN (n_39), .A1 (hfn_ipo_n5), .A2 (D[37]));
AND2_X1 i_0_38 (.ZN (n_38), .A1 (hfn_ipo_n5), .A2 (D[36]));
AND2_X1 i_0_37 (.ZN (n_37), .A1 (hfn_ipo_n5), .A2 (D[35]));
AND2_X1 i_0_36 (.ZN (n_36), .A1 (hfn_ipo_n5), .A2 (D[34]));
AND2_X1 i_0_35 (.ZN (n_35), .A1 (hfn_ipo_n5), .A2 (D[33]));
AND2_X1 i_0_34 (.ZN (n_34), .A1 (hfn_ipo_n6), .A2 (D[32]));
AND2_X1 i_0_33 (.ZN (n_33), .A1 (hfn_ipo_n6), .A2 (D[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (hfn_ipo_n6), .A2 (D[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (hfn_ipo_n6), .A2 (D[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (hfn_ipo_n6), .A2 (D[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (hfn_ipo_n6), .A2 (D[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (hfn_ipo_n6), .A2 (D[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (hfn_ipo_n6), .A2 (D[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (hfn_ipo_n6), .A2 (D[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (hfn_ipo_n6), .A2 (D[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (hfn_ipo_n6), .A2 (D[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (hfn_ipo_n6), .A2 (D[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (hfn_ipo_n6), .A2 (D[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (hfn_ipo_n6), .A2 (D[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (hfn_ipo_n6), .A2 (D[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (hfn_ipo_n5), .A2 (D[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (hfn_ipo_n5), .A2 (D[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (hfn_ipo_n5), .A2 (D[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (hfn_ipo_n5), .A2 (D[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (hfn_ipo_n5), .A2 (D[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (hfn_ipo_n5), .A2 (D[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (hfn_ipo_n5), .A2 (D[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (hfn_ipo_n5), .A2 (D[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (hfn_ipo_n5), .A2 (D[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (hfn_ipo_n5), .A2 (D[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (hfn_ipo_n5), .A2 (D[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (hfn_ipo_n5), .A2 (D[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (hfn_ipo_n5), .A2 (D[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (hfn_ipo_n5), .A2 (D[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (hfn_ipo_n5), .A2 (D[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (hfn_ipo_n5), .A2 (D[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (hfn_ipo_n5), .A2 (D[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (hfn_ipo_n5), .A2 (D[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (rst));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (rst));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (CTS_n_tid1_8), .D (n_2));
DFF_X1 \Q_reg[1]  (.Q (Q[1]), .CK (CTS_n_tid1_8), .D (n_3));
DFF_X1 \Q_reg[2]  (.Q (Q[2]), .CK (CTS_n_tid1_8), .D (n_4));
DFF_X1 \Q_reg[3]  (.Q (Q[3]), .CK (CTS_n_tid1_8), .D (n_5));
DFF_X1 \Q_reg[4]  (.Q (Q[4]), .CK (CTS_n_tid1_8), .D (n_6));
DFF_X1 \Q_reg[5]  (.Q (Q[5]), .CK (CTS_n_tid1_8), .D (n_7));
DFF_X1 \Q_reg[6]  (.Q (Q[6]), .CK (CTS_n_tid1_8), .D (n_8));
DFF_X1 \Q_reg[7]  (.Q (Q[7]), .CK (CTS_n_tid1_8), .D (n_9));
DFF_X1 \Q_reg[8]  (.Q (Q[8]), .CK (CTS_n_tid1_8), .D (n_10));
DFF_X1 \Q_reg[9]  (.Q (Q[9]), .CK (CTS_n_tid1_8), .D (n_11));
DFF_X1 \Q_reg[10]  (.Q (Q[10]), .CK (CTS_n_tid1_8), .D (n_12));
DFF_X1 \Q_reg[11]  (.Q (Q[11]), .CK (CTS_n_tid1_8), .D (n_13));
DFF_X1 \Q_reg[12]  (.Q (Q[12]), .CK (CTS_n_tid1_8), .D (n_14));
DFF_X1 \Q_reg[13]  (.Q (Q[13]), .CK (CTS_n_tid1_8), .D (n_15));
DFF_X1 \Q_reg[14]  (.Q (Q[14]), .CK (CTS_n_tid1_8), .D (n_16));
DFF_X1 \Q_reg[15]  (.Q (Q[15]), .CK (CTS_n_tid1_8), .D (n_17));
DFF_X1 \Q_reg[16]  (.Q (Q[16]), .CK (CTS_n_tid1_8), .D (n_18));
DFF_X1 \Q_reg[17]  (.Q (Q[17]), .CK (CTS_n_tid1_8), .D (n_19));
DFF_X1 \Q_reg[18]  (.Q (Q[18]), .CK (CTS_n_tid1_8), .D (n_20));
DFF_X1 \Q_reg[19]  (.Q (Q[19]), .CK (CTS_n_tid1_8), .D (n_21));
DFF_X1 \Q_reg[20]  (.Q (Q[20]), .CK (CTS_n_tid1_8), .D (n_22));
DFF_X1 \Q_reg[21]  (.Q (Q[21]), .CK (CTS_n_tid1_8), .D (n_23));
DFF_X1 \Q_reg[22]  (.Q (Q[22]), .CK (CTS_n_tid1_8), .D (n_24));
DFF_X1 \Q_reg[23]  (.Q (Q[23]), .CK (CTS_n_tid1_8), .D (n_25));
DFF_X1 \Q_reg[24]  (.Q (Q[24]), .CK (CTS_n_tid1_8), .D (n_26));
DFF_X1 \Q_reg[25]  (.Q (Q[25]), .CK (CTS_n_tid1_8), .D (n_27));
DFF_X1 \Q_reg[26]  (.Q (Q[26]), .CK (CTS_n_tid1_8), .D (n_28));
DFF_X1 \Q_reg[27]  (.Q (Q[27]), .CK (CTS_n_tid1_8), .D (n_29));
DFF_X1 \Q_reg[28]  (.Q (Q[28]), .CK (CTS_n_tid1_8), .D (n_30));
DFF_X1 \Q_reg[29]  (.Q (Q[29]), .CK (CTS_n_tid1_8), .D (n_31));
DFF_X1 \Q_reg[30]  (.Q (Q[30]), .CK (CTS_n_tid1_8), .D (n_32));
DFF_X1 \Q_reg[31]  (.Q (Q[31]), .CK (CTS_n_tid1_8), .D (n_33));
DFF_X1 \Q_reg[32]  (.Q (Q[32]), .CK (CTS_n_tid1_8), .D (n_34));
DFF_X1 \Q_reg[33]  (.Q (Q[33]), .CK (CTS_n_tid1_8), .D (n_35));
DFF_X1 \Q_reg[34]  (.Q (Q[34]), .CK (CTS_n_tid1_8), .D (n_36));
DFF_X1 \Q_reg[35]  (.Q (Q[35]), .CK (CTS_n_tid1_8), .D (n_37));
DFF_X1 \Q_reg[36]  (.Q (Q[36]), .CK (CTS_n_tid1_8), .D (n_38));
DFF_X1 \Q_reg[37]  (.Q (Q[37]), .CK (CTS_n_tid1_8), .D (n_39));
DFF_X1 \Q_reg[38]  (.Q (Q[38]), .CK (CTS_n_tid1_8), .D (n_40));
DFF_X1 \Q_reg[39]  (.Q (Q[39]), .CK (CTS_n_tid1_8), .D (n_41));
DFF_X1 \Q_reg[40]  (.Q (Q[40]), .CK (CTS_n_tid1_8), .D (n_42));
DFF_X1 \Q_reg[41]  (.Q (Q[41]), .CK (CTS_n_tid1_8), .D (n_43));
DFF_X1 \Q_reg[42]  (.Q (Q[42]), .CK (CTS_n_tid1_8), .D (n_44));
DFF_X1 \Q_reg[43]  (.Q (Q[43]), .CK (CTS_n_tid1_8), .D (n_45));
DFF_X1 \Q_reg[44]  (.Q (Q[44]), .CK (CTS_n_tid1_8), .D (n_46));
DFF_X1 \Q_reg[45]  (.Q (Q[45]), .CK (CTS_n_tid1_8), .D (n_47));
DFF_X1 \Q_reg[46]  (.Q (Q[46]), .CK (CTS_n_tid1_8), .D (n_48));
DFF_X1 \Q_reg[47]  (.Q (Q[47]), .CK (CTS_n_tid1_8), .D (n_49));
DFF_X1 \Q_reg[48]  (.Q (Q[48]), .CK (CTS_n_tid1_8), .D (n_50));
DFF_X1 \Q_reg[49]  (.Q (Q[49]), .CK (CTS_n_tid1_8), .D (n_51));
DFF_X1 \Q_reg[50]  (.Q (Q[50]), .CK (CTS_n_tid1_8), .D (n_52));
DFF_X1 \Q_reg[51]  (.Q (Q[51]), .CK (CTS_n_tid1_8), .D (n_53));
DFF_X1 \Q_reg[52]  (.Q (Q[52]), .CK (CTS_n_tid1_8), .D (n_54));
DFF_X1 \Q_reg[53]  (.Q (Q[53]), .CK (CTS_n_tid1_8), .D (n_55));
DFF_X1 \Q_reg[54]  (.Q (Q[54]), .CK (CTS_n_tid1_8), .D (n_56));
DFF_X1 \Q_reg[55]  (.Q (Q[55]), .CK (CTS_n_tid1_8), .D (n_57));
DFF_X1 \Q_reg[56]  (.Q (Q[56]), .CK (CTS_n_tid1_8), .D (n_58));
DFF_X1 \Q_reg[57]  (.Q (Q[57]), .CK (CTS_n_tid1_8), .D (n_59));
DFF_X1 \Q_reg[58]  (.Q (Q[58]), .CK (CTS_n_tid1_8), .D (n_60));
DFF_X1 \Q_reg[59]  (.Q (Q[59]), .CK (CTS_n_tid1_8), .D (n_61));
DFF_X1 \Q_reg[60]  (.Q (Q[60]), .CK (CTS_n_tid1_8), .D (n_62));
DFF_X1 \Q_reg[61]  (.Q (Q[61]), .CK (CTS_n_tid1_8), .D (n_63));
DFF_X1 \Q_reg[62]  (.Q (Q[62]), .CK (CTS_n_tid1_8), .D (n_64));
DFF_X1 \Q_reg[63]  (.Q (Q[63]), .CK (CTS_n_tid1_8), .D (n_65));
CLKGATETST_X8 clk_gate_Q_reg (.GCK (CTS_n_tid1_9), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
BUF_X2 hfn_ipo_c5 (.Z (hfn_ipo_n5), .A (n_0_0));
CLKBUF_X1 hfn_ipo_c6 (.Z (hfn_ipo_n6), .A (n_0_0));
CLKBUF_X3 CTS_L3_c_tid1_9 (.Z (CTS_n_tid1_8), .A (CTS_n_tid1_9));

endmodule //buffer__parameterized0

module datapath (b, a, p_0);

output [63:0] p_0;
input [31:0] a;
input [31:0] b;
wire n_2818;
wire n_3231;
wire n_1;
wire n_0;
wire n_2786;
wire n_2817;
wire n_2848;
wire n_3;
wire n_2;
wire n_2877;
wire n_5;
wire n_4;
wire n_2754;
wire n_2785;
wire n_2816;
wire n_7;
wire n_6;
wire n_2847;
wire n_2876;
wire n_9;
wire n_8;
wire n_11;
wire n_10;
wire n_2722;
wire n_2753;
wire n_2784;
wire n_13;
wire n_12;
wire n_2815;
wire n_2846;
wire n_2875;
wire n_15;
wire n_14;
wire n_17;
wire n_16;
wire n_19;
wire n_18;
wire n_2690;
wire n_2721;
wire n_2752;
wire n_21;
wire n_20;
wire n_2783;
wire n_2814;
wire n_2845;
wire n_23;
wire n_22;
wire n_2874;
wire n_25;
wire n_24;
wire n_27;
wire n_26;
wire n_29;
wire n_28;
wire n_2658;
wire n_2689;
wire n_2720;
wire n_31;
wire n_30;
wire n_2751;
wire n_2782;
wire n_2813;
wire n_33;
wire n_32;
wire n_2844;
wire n_2873;
wire n_35;
wire n_34;
wire n_37;
wire n_36;
wire n_39;
wire n_38;
wire n_41;
wire n_40;
wire n_2626;
wire n_2657;
wire n_2688;
wire n_43;
wire n_42;
wire n_2719;
wire n_2750;
wire n_2781;
wire n_45;
wire n_44;
wire n_2812;
wire n_2843;
wire n_2872;
wire n_47;
wire n_46;
wire n_49;
wire n_48;
wire n_51;
wire n_50;
wire n_53;
wire n_52;
wire n_55;
wire n_54;
wire n_2594;
wire n_2625;
wire n_2656;
wire n_57;
wire n_56;
wire n_2687;
wire n_2718;
wire n_2749;
wire n_59;
wire n_58;
wire n_2780;
wire n_2811;
wire n_2842;
wire n_61;
wire n_60;
wire n_2871;
wire n_63;
wire n_62;
wire n_65;
wire n_64;
wire n_67;
wire n_66;
wire n_69;
wire n_68;
wire n_71;
wire n_70;
wire n_2562;
wire n_2593;
wire n_2624;
wire n_73;
wire n_72;
wire n_2655;
wire n_2686;
wire n_2717;
wire n_75;
wire n_74;
wire n_2748;
wire n_2779;
wire n_2810;
wire n_77;
wire n_76;
wire n_2841;
wire n_2870;
wire n_79;
wire n_78;
wire n_81;
wire n_80;
wire n_83;
wire n_82;
wire n_85;
wire n_84;
wire n_87;
wire n_86;
wire n_89;
wire n_88;
wire n_2530;
wire n_2561;
wire n_2592;
wire n_91;
wire n_90;
wire n_2623;
wire n_2654;
wire n_2685;
wire n_93;
wire n_92;
wire n_2716;
wire n_2747;
wire n_2778;
wire n_95;
wire n_94;
wire n_2809;
wire n_2840;
wire n_2869;
wire n_97;
wire n_96;
wire n_99;
wire n_98;
wire n_101;
wire n_100;
wire n_103;
wire n_102;
wire n_105;
wire n_104;
wire n_107;
wire n_106;
wire n_109;
wire n_108;
wire n_2498;
wire n_2529;
wire n_2560;
wire n_111;
wire n_110;
wire n_2591;
wire n_2622;
wire n_2653;
wire n_113;
wire n_112;
wire n_2684;
wire n_2715;
wire n_2746;
wire n_115;
wire n_114;
wire n_2777;
wire n_2808;
wire n_2839;
wire n_117;
wire n_116;
wire n_2868;
wire n_119;
wire n_118;
wire n_121;
wire n_120;
wire n_123;
wire n_122;
wire n_125;
wire n_124;
wire n_127;
wire n_126;
wire n_129;
wire n_128;
wire n_131;
wire n_130;
wire n_2466;
wire n_2497;
wire n_2528;
wire n_133;
wire n_132;
wire n_2559;
wire n_2590;
wire n_2621;
wire n_135;
wire n_134;
wire n_2652;
wire n_2683;
wire n_2714;
wire n_137;
wire n_136;
wire n_2745;
wire n_2776;
wire n_2807;
wire n_139;
wire n_138;
wire n_2838;
wire n_2867;
wire n_141;
wire n_140;
wire n_143;
wire n_142;
wire n_145;
wire n_144;
wire n_147;
wire n_146;
wire n_149;
wire n_148;
wire n_151;
wire n_150;
wire n_153;
wire n_152;
wire n_155;
wire n_154;
wire n_2434;
wire n_2465;
wire n_2496;
wire n_157;
wire n_156;
wire n_2527;
wire n_2558;
wire n_2589;
wire n_159;
wire n_158;
wire n_2620;
wire n_2651;
wire n_2682;
wire n_161;
wire n_160;
wire n_2713;
wire n_2744;
wire n_2775;
wire n_163;
wire n_162;
wire n_2806;
wire n_2837;
wire n_2866;
wire n_165;
wire n_164;
wire n_167;
wire n_166;
wire n_169;
wire n_168;
wire n_171;
wire n_170;
wire n_173;
wire n_172;
wire n_175;
wire n_174;
wire n_177;
wire n_176;
wire n_179;
wire n_178;
wire n_181;
wire n_180;
wire n_2402;
wire n_2433;
wire n_2464;
wire n_183;
wire n_182;
wire n_2495;
wire n_2526;
wire n_2557;
wire n_185;
wire n_184;
wire n_2588;
wire n_2619;
wire n_2650;
wire n_187;
wire n_186;
wire n_2681;
wire n_2712;
wire n_2743;
wire n_189;
wire n_188;
wire n_2774;
wire n_2805;
wire n_2836;
wire n_191;
wire n_190;
wire n_2865;
wire n_193;
wire n_192;
wire n_195;
wire n_194;
wire n_197;
wire n_196;
wire n_199;
wire n_198;
wire n_201;
wire n_200;
wire n_203;
wire n_202;
wire n_205;
wire n_204;
wire n_207;
wire n_206;
wire n_209;
wire n_208;
wire n_2370;
wire n_2401;
wire n_2432;
wire n_211;
wire n_210;
wire n_2463;
wire n_2494;
wire n_2525;
wire n_213;
wire n_212;
wire n_2556;
wire n_2587;
wire n_2618;
wire n_215;
wire n_214;
wire n_2649;
wire n_2680;
wire n_2711;
wire n_217;
wire n_216;
wire n_2742;
wire n_2773;
wire n_2804;
wire n_219;
wire n_218;
wire n_2835;
wire n_2864;
wire n_221;
wire n_220;
wire n_223;
wire n_222;
wire n_225;
wire n_224;
wire n_227;
wire n_226;
wire n_229;
wire n_228;
wire n_231;
wire n_230;
wire n_233;
wire n_232;
wire n_235;
wire n_234;
wire n_237;
wire n_236;
wire n_239;
wire n_238;
wire n_2338;
wire n_2369;
wire n_2400;
wire n_241;
wire n_240;
wire n_2431;
wire n_2462;
wire n_2493;
wire n_243;
wire n_242;
wire n_2524;
wire n_2555;
wire n_2586;
wire n_245;
wire n_244;
wire n_2617;
wire n_2648;
wire n_2679;
wire n_247;
wire n_246;
wire n_2710;
wire n_2741;
wire n_2772;
wire n_249;
wire n_248;
wire n_2803;
wire n_2834;
wire n_2863;
wire n_251;
wire n_250;
wire n_253;
wire n_252;
wire n_255;
wire n_254;
wire n_257;
wire n_256;
wire n_259;
wire n_258;
wire n_261;
wire n_260;
wire n_263;
wire n_262;
wire n_265;
wire n_264;
wire n_267;
wire n_266;
wire n_269;
wire n_268;
wire n_271;
wire n_270;
wire n_2306;
wire n_2337;
wire n_2368;
wire n_273;
wire n_272;
wire n_2399;
wire n_2430;
wire n_2461;
wire n_275;
wire n_274;
wire n_2492;
wire n_2523;
wire n_2554;
wire n_277;
wire n_276;
wire n_2585;
wire n_2616;
wire n_2647;
wire n_279;
wire n_278;
wire n_2678;
wire n_2709;
wire n_2740;
wire n_281;
wire n_280;
wire n_2771;
wire n_2802;
wire n_2833;
wire n_283;
wire n_282;
wire n_2862;
wire n_285;
wire n_284;
wire n_287;
wire n_286;
wire n_289;
wire n_288;
wire n_291;
wire n_290;
wire n_293;
wire n_292;
wire n_295;
wire n_294;
wire n_297;
wire n_296;
wire n_299;
wire n_298;
wire n_301;
wire n_300;
wire n_303;
wire n_302;
wire n_305;
wire n_304;
wire n_2274;
wire n_2305;
wire n_2336;
wire n_307;
wire n_306;
wire n_2367;
wire n_2398;
wire n_2429;
wire n_309;
wire n_308;
wire n_2460;
wire n_2491;
wire n_2522;
wire n_311;
wire n_310;
wire n_2553;
wire n_2584;
wire n_2615;
wire n_313;
wire n_312;
wire n_2646;
wire n_2677;
wire n_2708;
wire n_315;
wire n_314;
wire n_2739;
wire n_2770;
wire n_2801;
wire n_317;
wire n_316;
wire n_2832;
wire n_2861;
wire n_319;
wire n_318;
wire n_321;
wire n_320;
wire n_323;
wire n_322;
wire n_325;
wire n_324;
wire n_327;
wire n_326;
wire n_329;
wire n_328;
wire n_331;
wire n_330;
wire n_333;
wire n_332;
wire n_335;
wire n_334;
wire n_337;
wire n_336;
wire n_339;
wire n_338;
wire n_341;
wire n_340;
wire n_2242;
wire n_2273;
wire n_2304;
wire n_343;
wire n_342;
wire n_2335;
wire n_2366;
wire n_2397;
wire n_345;
wire n_344;
wire n_2428;
wire n_2459;
wire n_2490;
wire n_347;
wire n_346;
wire n_2521;
wire n_2552;
wire n_2583;
wire n_349;
wire n_348;
wire n_2614;
wire n_2645;
wire n_2676;
wire n_351;
wire n_350;
wire n_2707;
wire n_2738;
wire n_2769;
wire n_353;
wire n_352;
wire n_2800;
wire n_2831;
wire n_2860;
wire n_355;
wire n_354;
wire n_357;
wire n_356;
wire n_359;
wire n_358;
wire n_361;
wire n_360;
wire n_363;
wire n_362;
wire n_365;
wire n_364;
wire n_367;
wire n_366;
wire n_369;
wire n_368;
wire n_371;
wire n_370;
wire n_373;
wire n_372;
wire n_375;
wire n_374;
wire n_377;
wire n_376;
wire n_379;
wire n_378;
wire n_2210;
wire n_2241;
wire n_2272;
wire n_381;
wire n_380;
wire n_2303;
wire n_2334;
wire n_2365;
wire n_383;
wire n_382;
wire n_2396;
wire n_2427;
wire n_2458;
wire n_385;
wire n_384;
wire n_2489;
wire n_2520;
wire n_2551;
wire n_387;
wire n_386;
wire n_2582;
wire n_2613;
wire n_2644;
wire n_389;
wire n_388;
wire n_2675;
wire n_2706;
wire n_2737;
wire n_391;
wire n_390;
wire n_2768;
wire n_2799;
wire n_2830;
wire n_393;
wire n_392;
wire n_2859;
wire n_395;
wire n_394;
wire n_397;
wire n_396;
wire n_399;
wire n_398;
wire n_401;
wire n_400;
wire n_403;
wire n_402;
wire n_405;
wire n_404;
wire n_407;
wire n_406;
wire n_409;
wire n_408;
wire n_411;
wire n_410;
wire n_413;
wire n_412;
wire n_415;
wire n_414;
wire n_417;
wire n_416;
wire n_419;
wire n_418;
wire n_2178;
wire n_2209;
wire n_2240;
wire n_421;
wire n_420;
wire n_2271;
wire n_2302;
wire n_2333;
wire n_423;
wire n_422;
wire n_2364;
wire n_2395;
wire n_2426;
wire n_425;
wire n_424;
wire n_2457;
wire n_2488;
wire n_2519;
wire n_427;
wire n_426;
wire n_2550;
wire n_2581;
wire n_2612;
wire n_429;
wire n_428;
wire n_2643;
wire n_2674;
wire n_2705;
wire n_431;
wire n_430;
wire n_2736;
wire n_2767;
wire n_2798;
wire n_433;
wire n_432;
wire n_2829;
wire n_2858;
wire n_435;
wire n_434;
wire n_437;
wire n_436;
wire n_439;
wire n_438;
wire n_441;
wire n_440;
wire n_443;
wire n_442;
wire n_445;
wire n_444;
wire n_447;
wire n_446;
wire n_449;
wire n_448;
wire n_451;
wire n_450;
wire n_453;
wire n_452;
wire n_455;
wire n_454;
wire n_457;
wire n_456;
wire n_459;
wire n_458;
wire n_461;
wire n_460;
wire n_2146;
wire n_2177;
wire n_2208;
wire n_463;
wire n_462;
wire n_2239;
wire n_2270;
wire n_2301;
wire n_465;
wire n_464;
wire n_2332;
wire n_2363;
wire n_2394;
wire n_467;
wire n_466;
wire n_2425;
wire n_2456;
wire n_2487;
wire n_469;
wire n_468;
wire n_2518;
wire n_2549;
wire n_2580;
wire n_471;
wire n_470;
wire n_2611;
wire n_2642;
wire n_2673;
wire n_473;
wire n_472;
wire n_2704;
wire n_2735;
wire n_2766;
wire n_475;
wire n_474;
wire n_2797;
wire n_2828;
wire n_2857;
wire n_477;
wire n_476;
wire n_479;
wire n_478;
wire n_481;
wire n_480;
wire n_483;
wire n_482;
wire n_485;
wire n_484;
wire n_487;
wire n_486;
wire n_489;
wire n_488;
wire n_491;
wire n_490;
wire n_493;
wire n_492;
wire n_495;
wire n_494;
wire n_497;
wire n_496;
wire n_499;
wire n_498;
wire n_501;
wire n_500;
wire n_503;
wire n_502;
wire n_505;
wire n_504;
wire n_2114;
wire n_2145;
wire n_2176;
wire n_507;
wire n_506;
wire n_2207;
wire n_2238;
wire n_2269;
wire n_509;
wire n_508;
wire n_2300;
wire n_2331;
wire n_2362;
wire n_511;
wire n_510;
wire n_2393;
wire n_2424;
wire n_2455;
wire n_513;
wire n_512;
wire n_2486;
wire n_2517;
wire n_2548;
wire n_515;
wire n_514;
wire n_2579;
wire n_2610;
wire n_2641;
wire n_517;
wire n_516;
wire n_2672;
wire n_2703;
wire n_2734;
wire n_519;
wire n_518;
wire n_2765;
wire n_2796;
wire n_2827;
wire n_521;
wire n_520;
wire n_2856;
wire n_523;
wire n_522;
wire n_525;
wire n_524;
wire n_527;
wire n_526;
wire n_529;
wire n_528;
wire n_531;
wire n_530;
wire n_533;
wire n_532;
wire n_535;
wire n_534;
wire n_537;
wire n_536;
wire n_539;
wire n_538;
wire n_541;
wire n_540;
wire n_543;
wire n_542;
wire n_545;
wire n_544;
wire n_547;
wire n_546;
wire n_549;
wire n_548;
wire n_551;
wire n_550;
wire n_2082;
wire n_2113;
wire n_2144;
wire n_553;
wire n_552;
wire n_2175;
wire n_2206;
wire n_2237;
wire n_555;
wire n_554;
wire n_2268;
wire n_2299;
wire n_2330;
wire n_557;
wire n_556;
wire n_2361;
wire n_2392;
wire n_2423;
wire n_559;
wire n_558;
wire n_2454;
wire n_2485;
wire n_2516;
wire n_561;
wire n_560;
wire n_2547;
wire n_2578;
wire n_2609;
wire n_563;
wire n_562;
wire n_2640;
wire n_2671;
wire n_2702;
wire n_565;
wire n_564;
wire n_2733;
wire n_2764;
wire n_2795;
wire n_567;
wire n_566;
wire n_2826;
wire n_2855;
wire n_569;
wire n_568;
wire n_571;
wire n_570;
wire n_573;
wire n_572;
wire n_575;
wire n_574;
wire n_577;
wire n_576;
wire n_579;
wire n_578;
wire n_581;
wire n_580;
wire n_583;
wire n_582;
wire n_585;
wire n_584;
wire n_587;
wire n_586;
wire n_589;
wire n_588;
wire n_591;
wire n_590;
wire n_593;
wire n_592;
wire n_595;
wire n_594;
wire n_597;
wire n_596;
wire n_599;
wire n_598;
wire n_2050;
wire n_2081;
wire n_2112;
wire n_601;
wire n_600;
wire n_2143;
wire n_2174;
wire n_2205;
wire n_603;
wire n_602;
wire n_2236;
wire n_2267;
wire n_2298;
wire n_605;
wire n_604;
wire n_2329;
wire n_2360;
wire n_2391;
wire n_607;
wire n_606;
wire n_2422;
wire n_2453;
wire n_2484;
wire n_609;
wire n_608;
wire n_2515;
wire n_2546;
wire n_2577;
wire n_611;
wire n_610;
wire n_2608;
wire n_2639;
wire n_2670;
wire n_613;
wire n_612;
wire n_2701;
wire n_2732;
wire n_2763;
wire n_615;
wire n_614;
wire n_2794;
wire n_2825;
wire n_2854;
wire n_617;
wire n_616;
wire n_619;
wire n_618;
wire n_621;
wire n_620;
wire n_623;
wire n_622;
wire n_625;
wire n_624;
wire n_627;
wire n_626;
wire n_629;
wire n_628;
wire n_631;
wire n_630;
wire n_633;
wire n_632;
wire n_635;
wire n_634;
wire n_637;
wire n_636;
wire n_639;
wire n_638;
wire n_641;
wire n_640;
wire n_643;
wire n_642;
wire n_645;
wire n_644;
wire n_647;
wire n_646;
wire n_649;
wire n_648;
wire n_2018;
wire n_2049;
wire n_2080;
wire n_651;
wire n_650;
wire n_2111;
wire n_2142;
wire n_2173;
wire n_653;
wire n_652;
wire n_2204;
wire n_2235;
wire n_2266;
wire n_655;
wire n_654;
wire n_2297;
wire n_2328;
wire n_2359;
wire n_657;
wire n_656;
wire n_2390;
wire n_2421;
wire n_2452;
wire n_659;
wire n_658;
wire n_2483;
wire n_2514;
wire n_2545;
wire n_661;
wire n_660;
wire n_2576;
wire n_2607;
wire n_2638;
wire n_663;
wire n_662;
wire n_2669;
wire n_2700;
wire n_2731;
wire n_665;
wire n_664;
wire n_2762;
wire n_2793;
wire n_2824;
wire n_667;
wire n_666;
wire n_2853;
wire n_669;
wire n_668;
wire n_671;
wire n_670;
wire n_673;
wire n_672;
wire n_675;
wire n_674;
wire n_677;
wire n_676;
wire n_679;
wire n_678;
wire n_681;
wire n_680;
wire n_683;
wire n_682;
wire n_685;
wire n_684;
wire n_687;
wire n_686;
wire n_689;
wire n_688;
wire n_691;
wire n_690;
wire n_693;
wire n_692;
wire n_695;
wire n_694;
wire n_697;
wire n_696;
wire n_699;
wire n_698;
wire n_701;
wire n_700;
wire n_1986;
wire n_2017;
wire n_2048;
wire n_703;
wire n_702;
wire n_2079;
wire n_2110;
wire n_2141;
wire n_705;
wire n_704;
wire n_2172;
wire n_2203;
wire n_2234;
wire n_707;
wire n_706;
wire n_2265;
wire n_2296;
wire n_2327;
wire n_709;
wire n_708;
wire n_2358;
wire n_2389;
wire n_2420;
wire n_711;
wire n_710;
wire n_2451;
wire n_2482;
wire n_2513;
wire n_713;
wire n_712;
wire n_2544;
wire n_2575;
wire n_2606;
wire n_715;
wire n_714;
wire n_2637;
wire n_2668;
wire n_2699;
wire n_717;
wire n_716;
wire n_2730;
wire n_2761;
wire n_2792;
wire n_719;
wire n_718;
wire n_2823;
wire n_2852;
wire n_721;
wire n_720;
wire n_723;
wire n_722;
wire n_725;
wire n_724;
wire n_727;
wire n_726;
wire n_729;
wire n_728;
wire n_731;
wire n_730;
wire n_733;
wire n_732;
wire n_735;
wire n_734;
wire n_737;
wire n_736;
wire n_739;
wire n_738;
wire n_741;
wire n_740;
wire n_743;
wire n_742;
wire n_745;
wire n_744;
wire n_747;
wire n_746;
wire n_749;
wire n_748;
wire n_751;
wire n_750;
wire n_753;
wire n_752;
wire n_755;
wire n_754;
wire n_1954;
wire n_1985;
wire n_2016;
wire n_757;
wire n_756;
wire n_2047;
wire n_2078;
wire n_2109;
wire n_759;
wire n_758;
wire n_2140;
wire n_2171;
wire n_2202;
wire n_761;
wire n_760;
wire n_2233;
wire n_2264;
wire n_2295;
wire n_763;
wire n_762;
wire n_2326;
wire n_2357;
wire n_2388;
wire n_765;
wire n_764;
wire n_2419;
wire n_2450;
wire n_2481;
wire n_767;
wire n_766;
wire n_2512;
wire n_2543;
wire n_2574;
wire n_769;
wire n_768;
wire n_2605;
wire n_2636;
wire n_2667;
wire n_771;
wire n_770;
wire n_2698;
wire n_2729;
wire n_2760;
wire n_773;
wire n_772;
wire n_2791;
wire n_2822;
wire n_2851;
wire n_775;
wire n_774;
wire n_777;
wire n_776;
wire n_779;
wire n_778;
wire n_781;
wire n_780;
wire n_783;
wire n_782;
wire n_785;
wire n_784;
wire n_787;
wire n_786;
wire n_789;
wire n_788;
wire n_791;
wire n_790;
wire n_793;
wire n_792;
wire n_795;
wire n_794;
wire n_797;
wire n_796;
wire n_799;
wire n_798;
wire n_801;
wire n_800;
wire n_803;
wire n_802;
wire n_805;
wire n_804;
wire n_807;
wire n_806;
wire n_809;
wire n_808;
wire n_811;
wire n_810;
wire n_1922;
wire n_1953;
wire n_1984;
wire n_813;
wire n_812;
wire n_2015;
wire n_2046;
wire n_2077;
wire n_815;
wire n_814;
wire n_2108;
wire n_2139;
wire n_2170;
wire n_817;
wire n_816;
wire n_2201;
wire n_2232;
wire n_2263;
wire n_819;
wire n_818;
wire n_2294;
wire n_2325;
wire n_2356;
wire n_821;
wire n_820;
wire n_2387;
wire n_2418;
wire n_2449;
wire n_823;
wire n_822;
wire n_2480;
wire n_2511;
wire n_2542;
wire n_825;
wire n_824;
wire n_2573;
wire n_2604;
wire n_2635;
wire n_827;
wire n_826;
wire n_2666;
wire n_2697;
wire n_2728;
wire n_829;
wire n_828;
wire n_2759;
wire n_2790;
wire n_2821;
wire n_831;
wire n_830;
wire n_2850;
wire n_833;
wire n_832;
wire n_835;
wire n_834;
wire n_837;
wire n_836;
wire n_839;
wire n_838;
wire n_841;
wire n_840;
wire n_843;
wire n_842;
wire n_845;
wire n_844;
wire n_847;
wire n_846;
wire n_849;
wire n_848;
wire n_851;
wire n_850;
wire n_853;
wire n_852;
wire n_855;
wire n_854;
wire n_857;
wire n_856;
wire n_859;
wire n_858;
wire n_861;
wire n_860;
wire n_863;
wire n_862;
wire n_865;
wire n_864;
wire n_867;
wire n_866;
wire n_869;
wire n_868;
wire n_1890;
wire n_1921;
wire n_1952;
wire n_871;
wire n_870;
wire n_1983;
wire n_2014;
wire n_2045;
wire n_873;
wire n_872;
wire n_2076;
wire n_2107;
wire n_2138;
wire n_875;
wire n_874;
wire n_2169;
wire n_2200;
wire n_2231;
wire n_877;
wire n_876;
wire n_2262;
wire n_2293;
wire n_2324;
wire n_879;
wire n_878;
wire n_2355;
wire n_2386;
wire n_2417;
wire n_881;
wire n_880;
wire n_2448;
wire n_2479;
wire n_2510;
wire n_883;
wire n_882;
wire n_2541;
wire n_2572;
wire n_2603;
wire n_885;
wire n_884;
wire n_2634;
wire n_2665;
wire n_2696;
wire n_887;
wire n_886;
wire n_2727;
wire n_2758;
wire n_2789;
wire n_889;
wire n_888;
wire n_2820;
wire n_2849;
wire n_891;
wire n_890;
wire n_893;
wire n_892;
wire n_895;
wire n_894;
wire n_897;
wire n_896;
wire n_899;
wire n_898;
wire n_901;
wire n_900;
wire n_903;
wire n_902;
wire n_905;
wire n_904;
wire n_907;
wire n_906;
wire n_909;
wire n_908;
wire n_911;
wire n_910;
wire n_913;
wire n_912;
wire n_915;
wire n_914;
wire n_917;
wire n_916;
wire n_919;
wire n_918;
wire n_921;
wire n_920;
wire n_923;
wire n_922;
wire n_925;
wire n_924;
wire n_927;
wire n_926;
wire n_929;
wire n_928;
wire n_1889;
wire n_1920;
wire n_1951;
wire n_931;
wire n_930;
wire n_1982;
wire n_2013;
wire n_2044;
wire n_933;
wire n_932;
wire n_2075;
wire n_2106;
wire n_2137;
wire n_935;
wire n_934;
wire n_2168;
wire n_2199;
wire n_2230;
wire n_937;
wire n_936;
wire n_2261;
wire n_2292;
wire n_2323;
wire n_939;
wire n_938;
wire n_2354;
wire n_2385;
wire n_2416;
wire n_941;
wire n_940;
wire n_2447;
wire n_2478;
wire n_2509;
wire n_943;
wire n_942;
wire n_2540;
wire n_2571;
wire n_2602;
wire n_945;
wire n_944;
wire n_2633;
wire n_2664;
wire n_2695;
wire n_947;
wire n_946;
wire n_2726;
wire n_2757;
wire n_2788;
wire n_949;
wire n_948;
wire n_2819;
wire n_951;
wire n_950;
wire n_953;
wire n_952;
wire n_955;
wire n_954;
wire n_957;
wire n_956;
wire n_959;
wire n_958;
wire n_961;
wire n_960;
wire n_963;
wire n_962;
wire n_965;
wire n_964;
wire n_967;
wire n_966;
wire n_969;
wire n_968;
wire n_971;
wire n_970;
wire n_973;
wire n_972;
wire n_975;
wire n_974;
wire n_977;
wire n_976;
wire n_979;
wire n_978;
wire n_981;
wire n_980;
wire n_983;
wire n_982;
wire n_985;
wire n_984;
wire n_987;
wire n_986;
wire n_989;
wire n_988;
wire n_1888;
wire n_1919;
wire n_1950;
wire n_991;
wire n_990;
wire n_1981;
wire n_2012;
wire n_2043;
wire n_993;
wire n_992;
wire n_2074;
wire n_2105;
wire n_2136;
wire n_995;
wire n_994;
wire n_2167;
wire n_2198;
wire n_2229;
wire n_997;
wire n_996;
wire n_2260;
wire n_2291;
wire n_2322;
wire n_999;
wire n_998;
wire n_2353;
wire n_2384;
wire n_2415;
wire n_1001;
wire n_1000;
wire n_2446;
wire n_2477;
wire n_2508;
wire n_1003;
wire n_1002;
wire n_2539;
wire n_2570;
wire n_2601;
wire n_1005;
wire n_1004;
wire n_2632;
wire n_2663;
wire n_2694;
wire n_1007;
wire n_1006;
wire n_2725;
wire n_2756;
wire n_2787;
wire n_1009;
wire n_1008;
wire n_1011;
wire n_1010;
wire n_1013;
wire n_1012;
wire n_1015;
wire n_1014;
wire n_1017;
wire n_1016;
wire n_1019;
wire n_1018;
wire n_1021;
wire n_1020;
wire n_1023;
wire n_1022;
wire n_1025;
wire n_1024;
wire n_1027;
wire n_1026;
wire n_1029;
wire n_1028;
wire n_1031;
wire n_1030;
wire n_1033;
wire n_1032;
wire n_1035;
wire n_1034;
wire n_1037;
wire n_1036;
wire n_1039;
wire n_1038;
wire n_1041;
wire n_1040;
wire n_1043;
wire n_1042;
wire n_1045;
wire n_1044;
wire n_1047;
wire n_1046;
wire n_1887;
wire n_1918;
wire n_1949;
wire n_1049;
wire n_1048;
wire n_1980;
wire n_2011;
wire n_2042;
wire n_1051;
wire n_1050;
wire n_2073;
wire n_2104;
wire n_2135;
wire n_1053;
wire n_1052;
wire n_2166;
wire n_2197;
wire n_2228;
wire n_1055;
wire n_1054;
wire n_2259;
wire n_2290;
wire n_2321;
wire n_1057;
wire n_1056;
wire n_2352;
wire n_2383;
wire n_2414;
wire n_1059;
wire n_1058;
wire n_2445;
wire n_2476;
wire n_2507;
wire n_1061;
wire n_1060;
wire n_2538;
wire n_2569;
wire n_2600;
wire n_1063;
wire n_1062;
wire n_2631;
wire n_2662;
wire n_2693;
wire n_1065;
wire n_1064;
wire n_2724;
wire n_2755;
wire n_1067;
wire n_1066;
wire n_1069;
wire n_1068;
wire n_1071;
wire n_1070;
wire n_1073;
wire n_1072;
wire n_1075;
wire n_1074;
wire n_1077;
wire n_1076;
wire n_1079;
wire n_1078;
wire n_1081;
wire n_1080;
wire n_1083;
wire n_1082;
wire n_1085;
wire n_1084;
wire n_1087;
wire n_1086;
wire n_1089;
wire n_1088;
wire n_1091;
wire n_1090;
wire n_1093;
wire n_1092;
wire n_1095;
wire n_1094;
wire n_1097;
wire n_1096;
wire n_1099;
wire n_1098;
wire n_1101;
wire n_1100;
wire n_1103;
wire n_1102;
wire n_1886;
wire n_1917;
wire n_1948;
wire n_1105;
wire n_1104;
wire n_1979;
wire n_2010;
wire n_2041;
wire n_1107;
wire n_1106;
wire n_2072;
wire n_2103;
wire n_2134;
wire n_1109;
wire n_1108;
wire n_2165;
wire n_2196;
wire n_2227;
wire n_1111;
wire n_1110;
wire n_2258;
wire n_2289;
wire n_2320;
wire n_1113;
wire n_1112;
wire n_2351;
wire n_2382;
wire n_2413;
wire n_1115;
wire n_1114;
wire n_2444;
wire n_2475;
wire n_2506;
wire n_1117;
wire n_1116;
wire n_2537;
wire n_2568;
wire n_2599;
wire n_1119;
wire n_1118;
wire n_2630;
wire n_2661;
wire n_2692;
wire n_1121;
wire n_1120;
wire n_2723;
wire n_1123;
wire n_1122;
wire n_1125;
wire n_1124;
wire n_1127;
wire n_1126;
wire n_1129;
wire n_1128;
wire n_1131;
wire n_1130;
wire n_1133;
wire n_1132;
wire n_1135;
wire n_1134;
wire n_1137;
wire n_1136;
wire n_1139;
wire n_1138;
wire n_1141;
wire n_1140;
wire n_1143;
wire n_1142;
wire n_1145;
wire n_1144;
wire n_1147;
wire n_1146;
wire n_1149;
wire n_1148;
wire n_1151;
wire n_1150;
wire n_1153;
wire n_1152;
wire n_1155;
wire n_1154;
wire n_1157;
wire n_1156;
wire n_1885;
wire n_1916;
wire n_1947;
wire n_1159;
wire n_1158;
wire n_1978;
wire n_2009;
wire n_2040;
wire n_1161;
wire n_1160;
wire n_2071;
wire n_2102;
wire n_2133;
wire n_1163;
wire n_1162;
wire n_2164;
wire n_2195;
wire n_2226;
wire n_1165;
wire n_1164;
wire n_2257;
wire n_2288;
wire n_2319;
wire n_1167;
wire n_1166;
wire n_2350;
wire n_2381;
wire n_2412;
wire n_1169;
wire n_1168;
wire n_2443;
wire n_2474;
wire n_2505;
wire n_1171;
wire n_1170;
wire n_2536;
wire n_2567;
wire n_2598;
wire n_1173;
wire n_1172;
wire n_2629;
wire n_2660;
wire n_2691;
wire n_1175;
wire n_1174;
wire n_1177;
wire n_1176;
wire n_1179;
wire n_1178;
wire n_1181;
wire n_1180;
wire n_1183;
wire n_1182;
wire n_1185;
wire n_1184;
wire n_1187;
wire n_1186;
wire n_1189;
wire n_1188;
wire n_1191;
wire n_1190;
wire n_1193;
wire n_1192;
wire n_1195;
wire n_1194;
wire n_1197;
wire n_1196;
wire n_1199;
wire n_1198;
wire n_1201;
wire n_1200;
wire n_1203;
wire n_1202;
wire n_1205;
wire n_1204;
wire n_1207;
wire n_1206;
wire n_1209;
wire n_1208;
wire n_1884;
wire n_1915;
wire n_1946;
wire n_1211;
wire n_1210;
wire n_1977;
wire n_2008;
wire n_2039;
wire n_1213;
wire n_1212;
wire n_2070;
wire n_2101;
wire n_2132;
wire n_1215;
wire n_1214;
wire n_2163;
wire n_2194;
wire n_2225;
wire n_1217;
wire n_1216;
wire n_2256;
wire n_2287;
wire n_2318;
wire n_1219;
wire n_1218;
wire n_2349;
wire n_2380;
wire n_2411;
wire n_1221;
wire n_1220;
wire n_2442;
wire n_2473;
wire n_2504;
wire n_1223;
wire n_1222;
wire n_2535;
wire n_2566;
wire n_2597;
wire n_1225;
wire n_1224;
wire n_2628;
wire n_2659;
wire n_1227;
wire n_1226;
wire n_1229;
wire n_1228;
wire n_1231;
wire n_1230;
wire n_1233;
wire n_1232;
wire n_1235;
wire n_1234;
wire n_1237;
wire n_1236;
wire n_1239;
wire n_1238;
wire n_1241;
wire n_1240;
wire n_1243;
wire n_1242;
wire n_1245;
wire n_1244;
wire n_1247;
wire n_1246;
wire n_1249;
wire n_1248;
wire n_1251;
wire n_1250;
wire n_1253;
wire n_1252;
wire n_1255;
wire n_1254;
wire n_1257;
wire n_1256;
wire n_1259;
wire n_1258;
wire n_1883;
wire n_1914;
wire n_1945;
wire n_1261;
wire n_1260;
wire n_1976;
wire n_2007;
wire n_2038;
wire n_1263;
wire n_1262;
wire n_2069;
wire n_2100;
wire n_2131;
wire n_1265;
wire n_1264;
wire n_2162;
wire n_2193;
wire n_2224;
wire n_1267;
wire n_1266;
wire n_2255;
wire n_2286;
wire n_2317;
wire n_1269;
wire n_1268;
wire n_2348;
wire n_2379;
wire n_2410;
wire n_1271;
wire n_1270;
wire n_2441;
wire n_2472;
wire n_2503;
wire n_1273;
wire n_1272;
wire n_2534;
wire n_2565;
wire n_2596;
wire n_1275;
wire n_1274;
wire n_2627;
wire n_1277;
wire n_1276;
wire n_1279;
wire n_1278;
wire n_1281;
wire n_1280;
wire n_1283;
wire n_1282;
wire n_1285;
wire n_1284;
wire n_1287;
wire n_1286;
wire n_1289;
wire n_1288;
wire n_1291;
wire n_1290;
wire n_1293;
wire n_1292;
wire n_1295;
wire n_1294;
wire n_1297;
wire n_1296;
wire n_1299;
wire n_1298;
wire n_1301;
wire n_1300;
wire n_1303;
wire n_1302;
wire n_1305;
wire n_1304;
wire n_1307;
wire n_1306;
wire n_1882;
wire n_1913;
wire n_1944;
wire n_1309;
wire n_1308;
wire n_1975;
wire n_2006;
wire n_2037;
wire n_1311;
wire n_1310;
wire n_2068;
wire n_2099;
wire n_2130;
wire n_1313;
wire n_1312;
wire n_2161;
wire n_2192;
wire n_2223;
wire n_1315;
wire n_1314;
wire n_2254;
wire n_2285;
wire n_2316;
wire n_1317;
wire n_1316;
wire n_2347;
wire n_2378;
wire n_2409;
wire n_1319;
wire n_1318;
wire n_2440;
wire n_2471;
wire n_2502;
wire n_1321;
wire n_1320;
wire n_2533;
wire n_2564;
wire n_2595;
wire n_1323;
wire n_1322;
wire n_1325;
wire n_1324;
wire n_1327;
wire n_1326;
wire n_1329;
wire n_1328;
wire n_1331;
wire n_1330;
wire n_1333;
wire n_1332;
wire n_1335;
wire n_1334;
wire n_1337;
wire n_1336;
wire n_1339;
wire n_1338;
wire n_1341;
wire n_1340;
wire n_1343;
wire n_1342;
wire n_1345;
wire n_1344;
wire n_1347;
wire n_1346;
wire n_1349;
wire n_1348;
wire n_1351;
wire n_1350;
wire n_1353;
wire n_1352;
wire n_1881;
wire n_1912;
wire n_1943;
wire n_1355;
wire n_1354;
wire n_1974;
wire n_2005;
wire n_2036;
wire n_1357;
wire n_1356;
wire n_2067;
wire n_2098;
wire n_2129;
wire n_1359;
wire n_1358;
wire n_2160;
wire n_2191;
wire n_2222;
wire n_1361;
wire n_1360;
wire n_2253;
wire n_2284;
wire n_2315;
wire n_1363;
wire n_1362;
wire n_2346;
wire n_2377;
wire n_2408;
wire n_1365;
wire n_1364;
wire n_2439;
wire n_2470;
wire n_2501;
wire n_1367;
wire n_1366;
wire n_2532;
wire n_2563;
wire n_1369;
wire n_1368;
wire n_1371;
wire n_1370;
wire n_1373;
wire n_1372;
wire n_1375;
wire n_1374;
wire n_1377;
wire n_1376;
wire n_1379;
wire n_1378;
wire n_1381;
wire n_1380;
wire n_1383;
wire n_1382;
wire n_1385;
wire n_1384;
wire n_1387;
wire n_1386;
wire n_1389;
wire n_1388;
wire n_1391;
wire n_1390;
wire n_1393;
wire n_1392;
wire n_1395;
wire n_1394;
wire n_1397;
wire n_1396;
wire n_1880;
wire n_1911;
wire n_1942;
wire n_1399;
wire n_1398;
wire n_1973;
wire n_2004;
wire n_2035;
wire n_1401;
wire n_1400;
wire n_2066;
wire n_2097;
wire n_2128;
wire n_1403;
wire n_1402;
wire n_2159;
wire n_2190;
wire n_2221;
wire n_1405;
wire n_1404;
wire n_2252;
wire n_2283;
wire n_2314;
wire n_1407;
wire n_1406;
wire n_2345;
wire n_2376;
wire n_2407;
wire n_1409;
wire n_1408;
wire n_2438;
wire n_2469;
wire n_2500;
wire n_1411;
wire n_1410;
wire n_2531;
wire n_1413;
wire n_1412;
wire n_1415;
wire n_1414;
wire n_1417;
wire n_1416;
wire n_1419;
wire n_1418;
wire n_1421;
wire n_1420;
wire n_1423;
wire n_1422;
wire n_1425;
wire n_1424;
wire n_1427;
wire n_1426;
wire n_1429;
wire n_1428;
wire n_1431;
wire n_1430;
wire n_1433;
wire n_1432;
wire n_1435;
wire n_1434;
wire n_1437;
wire n_1436;
wire n_1439;
wire n_1438;
wire n_1879;
wire n_1910;
wire n_1941;
wire n_1441;
wire n_1440;
wire n_1972;
wire n_2003;
wire n_2034;
wire n_1443;
wire n_1442;
wire n_2065;
wire n_2096;
wire n_2127;
wire n_1445;
wire n_1444;
wire n_2158;
wire n_2189;
wire n_2220;
wire n_1447;
wire n_1446;
wire n_2251;
wire n_2282;
wire n_2313;
wire n_1449;
wire n_1448;
wire n_2344;
wire n_2375;
wire n_2406;
wire n_1451;
wire n_1450;
wire n_2437;
wire n_2468;
wire n_2499;
wire n_1453;
wire n_1452;
wire n_1455;
wire n_1454;
wire n_1457;
wire n_1456;
wire n_1459;
wire n_1458;
wire n_1461;
wire n_1460;
wire n_1463;
wire n_1462;
wire n_1465;
wire n_1464;
wire n_1467;
wire n_1466;
wire n_1469;
wire n_1468;
wire n_1471;
wire n_1470;
wire n_1473;
wire n_1472;
wire n_1475;
wire n_1474;
wire n_1477;
wire n_1476;
wire n_1479;
wire n_1478;
wire n_1878;
wire n_1909;
wire n_1940;
wire n_1481;
wire n_1480;
wire n_1971;
wire n_2002;
wire n_2033;
wire n_1483;
wire n_1482;
wire n_2064;
wire n_2095;
wire n_2126;
wire n_1485;
wire n_1484;
wire n_2157;
wire n_2188;
wire n_2219;
wire n_1487;
wire n_1486;
wire n_2250;
wire n_2281;
wire n_2312;
wire n_1489;
wire n_1488;
wire n_2343;
wire n_2374;
wire n_2405;
wire n_1491;
wire n_1490;
wire n_2436;
wire n_2467;
wire n_1493;
wire n_1492;
wire n_1495;
wire n_1494;
wire n_1497;
wire n_1496;
wire n_1499;
wire n_1498;
wire n_1501;
wire n_1500;
wire n_1503;
wire n_1502;
wire n_1505;
wire n_1504;
wire n_1507;
wire n_1506;
wire n_1509;
wire n_1508;
wire n_1511;
wire n_1510;
wire n_1513;
wire n_1512;
wire n_1515;
wire n_1514;
wire n_1517;
wire n_1516;
wire n_1877;
wire n_1908;
wire n_1939;
wire n_1519;
wire n_1518;
wire n_1970;
wire n_2001;
wire n_2032;
wire n_1521;
wire n_1520;
wire n_2063;
wire n_2094;
wire n_2125;
wire n_1523;
wire n_1522;
wire n_2156;
wire n_2187;
wire n_2218;
wire n_1525;
wire n_1524;
wire n_2249;
wire n_2280;
wire n_2311;
wire n_1527;
wire n_1526;
wire n_2342;
wire n_2373;
wire n_2404;
wire n_1529;
wire n_1528;
wire n_2435;
wire n_1531;
wire n_1530;
wire n_1533;
wire n_1532;
wire n_1535;
wire n_1534;
wire n_1537;
wire n_1536;
wire n_1539;
wire n_1538;
wire n_1541;
wire n_1540;
wire n_1543;
wire n_1542;
wire n_1545;
wire n_1544;
wire n_1547;
wire n_1546;
wire n_1549;
wire n_1548;
wire n_1551;
wire n_1550;
wire n_1553;
wire n_1552;
wire n_1876;
wire n_1907;
wire n_1938;
wire n_1555;
wire n_1554;
wire n_1969;
wire n_2000;
wire n_2031;
wire n_1557;
wire n_1556;
wire n_2062;
wire n_2093;
wire n_2124;
wire n_1559;
wire n_1558;
wire n_2155;
wire n_2186;
wire n_2217;
wire n_1561;
wire n_1560;
wire n_2248;
wire n_2279;
wire n_2310;
wire n_1563;
wire n_1562;
wire n_2341;
wire n_2372;
wire n_2403;
wire n_1565;
wire n_1564;
wire n_1567;
wire n_1566;
wire n_1569;
wire n_1568;
wire n_1571;
wire n_1570;
wire n_1573;
wire n_1572;
wire n_1575;
wire n_1574;
wire n_1577;
wire n_1576;
wire n_1579;
wire n_1578;
wire n_1581;
wire n_1580;
wire n_1583;
wire n_1582;
wire n_1585;
wire n_1584;
wire n_1587;
wire n_1586;
wire n_1875;
wire n_1906;
wire n_1937;
wire n_1589;
wire n_1588;
wire n_1968;
wire n_1999;
wire n_2030;
wire n_1591;
wire n_1590;
wire n_2061;
wire n_2092;
wire n_2123;
wire n_1593;
wire n_1592;
wire n_2154;
wire n_2185;
wire n_2216;
wire n_1595;
wire n_1594;
wire n_2247;
wire n_2278;
wire n_2309;
wire n_1597;
wire n_1596;
wire n_2340;
wire n_2371;
wire n_1599;
wire n_1598;
wire n_1601;
wire n_1600;
wire n_1603;
wire n_1602;
wire n_1605;
wire n_1604;
wire n_1607;
wire n_1606;
wire n_1609;
wire n_1608;
wire n_1611;
wire n_1610;
wire n_1613;
wire n_1612;
wire n_1615;
wire n_1614;
wire n_1617;
wire n_1616;
wire n_1619;
wire n_1618;
wire n_1874;
wire n_1905;
wire n_1936;
wire n_1621;
wire n_1620;
wire n_1967;
wire n_1998;
wire n_2029;
wire n_1623;
wire n_1622;
wire n_2060;
wire n_2091;
wire n_2122;
wire n_1625;
wire n_1624;
wire n_2153;
wire n_2184;
wire n_2215;
wire n_1627;
wire n_1626;
wire n_2246;
wire n_2277;
wire n_2308;
wire n_1629;
wire n_1628;
wire n_2339;
wire n_1631;
wire n_1630;
wire n_1633;
wire n_1632;
wire n_1635;
wire n_1634;
wire n_1637;
wire n_1636;
wire n_1639;
wire n_1638;
wire n_1641;
wire n_1640;
wire n_1643;
wire n_1642;
wire n_1645;
wire n_1644;
wire n_1647;
wire n_1646;
wire n_1649;
wire n_1648;
wire n_1873;
wire n_1904;
wire n_1935;
wire n_1651;
wire n_1650;
wire n_1966;
wire n_1997;
wire n_2028;
wire n_1653;
wire n_1652;
wire n_2059;
wire n_2090;
wire n_2121;
wire n_1655;
wire n_1654;
wire n_2152;
wire n_2183;
wire n_2214;
wire n_1657;
wire n_1656;
wire n_2245;
wire n_2276;
wire n_2307;
wire n_1659;
wire n_1658;
wire n_1661;
wire n_1660;
wire n_1663;
wire n_1662;
wire n_1665;
wire n_1664;
wire n_1667;
wire n_1666;
wire n_1669;
wire n_1668;
wire n_1671;
wire n_1670;
wire n_1673;
wire n_1672;
wire n_1675;
wire n_1674;
wire n_1677;
wire n_1676;
wire n_1872;
wire n_1903;
wire n_1934;
wire n_1679;
wire n_1678;
wire n_1965;
wire n_1996;
wire n_2027;
wire n_1681;
wire n_1680;
wire n_2058;
wire n_2089;
wire n_2120;
wire n_1683;
wire n_1682;
wire n_2151;
wire n_2182;
wire n_2213;
wire n_1685;
wire n_1684;
wire n_2244;
wire n_2275;
wire n_1687;
wire n_1686;
wire n_1689;
wire n_1688;
wire n_1691;
wire n_1690;
wire n_1693;
wire n_1692;
wire n_1695;
wire n_1694;
wire n_1697;
wire n_1696;
wire n_1699;
wire n_1698;
wire n_1701;
wire n_1700;
wire n_1703;
wire n_1702;
wire n_1871;
wire n_1902;
wire n_1933;
wire n_1705;
wire n_1704;
wire n_1964;
wire n_1995;
wire n_2026;
wire n_1707;
wire n_1706;
wire n_2057;
wire n_2088;
wire n_2119;
wire n_1709;
wire n_1708;
wire n_2150;
wire n_2181;
wire n_2212;
wire n_1711;
wire n_1710;
wire n_2243;
wire n_1713;
wire n_1712;
wire n_1715;
wire n_1714;
wire n_1717;
wire n_1716;
wire n_1719;
wire n_1718;
wire n_1721;
wire n_1720;
wire n_1723;
wire n_1722;
wire n_1725;
wire n_1724;
wire n_1727;
wire n_1726;
wire n_1870;
wire n_1901;
wire n_1932;
wire n_1729;
wire n_1728;
wire n_1963;
wire n_1994;
wire n_2025;
wire n_1731;
wire n_1730;
wire n_2056;
wire n_2087;
wire n_2118;
wire n_1733;
wire n_1732;
wire n_2149;
wire n_2180;
wire n_2211;
wire n_1735;
wire n_1734;
wire n_1737;
wire n_1736;
wire n_1739;
wire n_1738;
wire n_1741;
wire n_1740;
wire n_1743;
wire n_1742;
wire n_1745;
wire n_1744;
wire n_1747;
wire n_1746;
wire n_1749;
wire n_1748;
wire n_1869;
wire n_1900;
wire n_1931;
wire n_1751;
wire n_1750;
wire n_1962;
wire n_1993;
wire n_2024;
wire n_1753;
wire n_1752;
wire n_2055;
wire n_2086;
wire n_2117;
wire n_1755;
wire n_1754;
wire n_2148;
wire n_2179;
wire n_1757;
wire n_1756;
wire n_1759;
wire n_1758;
wire n_1761;
wire n_1760;
wire n_1763;
wire n_1762;
wire n_1765;
wire n_1764;
wire n_1767;
wire n_1766;
wire n_1769;
wire n_1768;
wire n_1868;
wire n_1899;
wire n_1930;
wire n_1771;
wire n_1770;
wire n_1961;
wire n_1992;
wire n_2023;
wire n_1773;
wire n_1772;
wire n_2054;
wire n_2085;
wire n_2116;
wire n_1775;
wire n_1774;
wire n_2147;
wire n_1777;
wire n_1776;
wire n_1779;
wire n_1778;
wire n_1781;
wire n_1780;
wire n_1783;
wire n_1782;
wire n_1785;
wire n_1784;
wire n_1787;
wire n_1786;
wire n_1867;
wire n_1898;
wire n_1929;
wire n_1789;
wire n_1788;
wire n_1960;
wire n_1991;
wire n_2022;
wire n_1791;
wire n_1790;
wire n_2053;
wire n_2084;
wire n_2115;
wire n_1793;
wire n_1792;
wire n_1795;
wire n_1794;
wire n_1797;
wire n_1796;
wire n_1799;
wire n_1798;
wire n_1801;
wire n_1800;
wire n_1803;
wire n_1802;
wire n_1866;
wire n_1897;
wire n_1928;
wire n_1805;
wire n_1804;
wire n_1959;
wire n_1990;
wire n_2021;
wire n_1807;
wire n_1806;
wire n_2052;
wire n_2083;
wire n_1809;
wire n_1808;
wire n_1811;
wire n_1810;
wire n_1813;
wire n_1812;
wire n_1815;
wire n_1814;
wire n_1817;
wire n_1816;
wire n_1865;
wire n_1896;
wire n_1927;
wire n_1819;
wire n_1818;
wire n_1958;
wire n_1989;
wire n_2020;
wire n_1821;
wire n_1820;
wire n_2051;
wire n_1823;
wire n_1822;
wire n_1825;
wire n_1824;
wire n_1827;
wire n_1826;
wire n_1829;
wire n_1828;
wire n_1864;
wire n_1895;
wire n_1926;
wire n_1831;
wire n_1830;
wire n_1957;
wire n_1988;
wire n_2019;
wire n_1833;
wire n_1832;
wire n_1835;
wire n_1834;
wire n_1837;
wire n_1836;
wire n_1839;
wire n_1838;
wire n_1863;
wire n_1894;
wire n_1925;
wire n_1841;
wire n_1840;
wire n_1956;
wire n_1987;
wire n_1843;
wire n_1842;
wire n_1845;
wire n_1844;
wire n_1847;
wire n_1846;
wire n_1862;
wire n_1893;
wire n_1924;
wire n_1849;
wire n_1848;
wire n_1955;
wire n_1851;
wire n_1850;
wire n_1853;
wire n_1852;
wire n_1861;
wire n_1892;
wire n_1923;
wire n_1855;
wire n_1854;
wire n_1857;
wire n_1856;
wire n_1860;
wire n_1891;
wire n_1859;
wire n_1858;
wire n_3309;
wire n_3276;
wire n_3275;
wire n_3274;
wire n_3273;
wire n_3272;
wire n_3271;
wire n_3270;
wire n_3269;
wire n_3268;
wire n_3267;
wire n_3266;
wire n_3265;
wire n_3264;
wire n_3263;
wire n_3262;
wire n_3261;
wire n_3260;
wire n_3259;
wire n_3258;
wire n_3257;
wire n_3256;
wire n_3255;
wire n_3254;
wire n_3253;
wire n_3252;
wire n_3251;
wire n_3250;
wire n_3249;
wire n_3248;
wire n_3247;
wire n_3246;
wire n_3308;
wire n_3277;
wire n_3307;
wire n_3306;
wire n_3305;
wire n_3304;
wire n_3303;
wire n_3302;
wire n_3301;
wire n_3300;
wire n_3299;
wire n_3298;
wire n_3297;
wire n_3296;
wire n_3295;
wire n_3294;
wire n_3293;
wire n_3292;
wire n_3291;
wire n_3290;
wire n_3289;
wire n_3288;
wire n_3287;
wire n_3286;
wire n_3285;
wire n_3284;
wire n_3283;
wire n_3282;
wire n_3281;
wire n_3280;
wire n_3279;
wire n_3278;
wire n_2878;
wire n_3230;
wire n_3233;
wire n_3232;
wire n_2879;
wire n_3229;
wire n_3235;
wire n_3228;
wire n_2880;
wire n_3236;
wire n_3226;
wire n_2881;
wire n_3225;
wire n_2888;
wire n_2887;
wire n_2884;
wire n_2885;
wire n_2882;
wire n_3222;
wire n_3213;
wire n_2889;
wire n_2883;
wire n_3223;
wire n_3217;
wire n_2886;
wire n_3220;
wire n_3218;
wire n_3224;
wire n_3215;
wire n_3211;
wire n_2896;
wire n_2895;
wire n_2892;
wire n_2893;
wire n_2890;
wire n_3208;
wire n_3199;
wire n_2897;
wire n_2891;
wire n_3209;
wire n_3203;
wire n_2894;
wire n_3206;
wire n_3204;
wire n_3210;
wire n_3201;
wire n_3197;
wire n_2904;
wire n_2903;
wire n_2900;
wire n_2901;
wire n_2898;
wire n_3194;
wire n_3185;
wire n_2905;
wire n_2899;
wire n_3195;
wire n_3189;
wire n_2902;
wire n_3192;
wire n_3190;
wire n_3196;
wire n_3187;
wire n_3183;
wire n_2912;
wire n_2911;
wire n_2908;
wire n_2909;
wire n_2906;
wire n_3149;
wire n_3139;
wire n_2913;
wire n_2907;
wire n_3148;
wire n_3151;
wire n_3141;
wire n_2910;
wire n_3150;
wire n_3146;
wire n_3143;
wire n_3153;
wire n_2941;
wire n_2920;
wire n_2919;
wire n_2916;
wire n_2917;
wire n_2914;
wire n_3177;
wire n_3121;
wire n_2921;
wire n_2915;
wire n_3176;
wire n_3179;
wire n_3123;
wire n_2918;
wire n_3178;
wire n_3182;
wire n_3125;
wire n_3181;
wire n_2939;
wire n_2928;
wire n_2927;
wire n_2924;
wire n_2925;
wire n_2922;
wire n_3160;
wire n_3133;
wire n_2929;
wire n_2923;
wire n_3159;
wire n_3162;
wire n_3135;
wire n_2926;
wire n_3161;
wire n_3157;
wire n_3137;
wire n_3164;
wire n_2937;
wire n_2936;
wire n_2935;
wire n_2932;
wire n_2933;
wire n_2930;
wire n_3169;
wire n_3127;
wire n_2943;
wire n_2931;
wire n_3168;
wire n_3171;
wire n_3130;
wire n_2934;
wire n_3170;
wire n_3166;
wire n_3131;
wire n_2938;
wire n_3132;
wire n_3156;
wire n_2940;
wire n_3120;
wire n_3174;
wire n_2942;
wire n_3138;
wire n_3145;
wire n_3172;
wire n_3245;
wire n_3244;
wire n_3118;
wire n_2950;
wire n_2949;
wire n_2946;
wire n_2947;
wire n_2944;
wire n_3087;
wire n_3077;
wire n_2951;
wire n_2945;
wire n_3086;
wire n_3089;
wire n_3079;
wire n_2948;
wire n_3088;
wire n_3084;
wire n_3081;
wire n_3091;
wire n_2979;
wire n_2958;
wire n_2957;
wire n_2954;
wire n_2955;
wire n_2952;
wire n_3112;
wire n_3070;
wire n_2959;
wire n_2953;
wire n_3111;
wire n_3114;
wire n_3072;
wire n_2956;
wire n_3113;
wire n_3117;
wire n_3074;
wire n_3116;
wire n_2977;
wire n_2966;
wire n_2965;
wire n_2962;
wire n_2963;
wire n_2960;
wire n_3098;
wire n_3056;
wire n_2967;
wire n_2961;
wire n_3097;
wire n_3100;
wire n_3058;
wire n_2964;
wire n_3099;
wire n_3095;
wire n_3060;
wire n_3102;
wire n_2976;
wire n_2975;
wire n_2973;
wire n_2972;
wire n_2969;
wire n_2968;
wire n_3066;
wire n_3106;
wire n_3063;
wire n_2981;
wire n_2970;
wire n_2971;
wire n_3105;
wire n_3064;
wire n_2974;
wire n_3107;
wire n_3067;
wire n_3068;
wire n_3055;
wire n_3094;
wire n_2978;
wire n_3069;
wire n_3109;
wire n_2980;
wire n_3076;
wire n_3083;
wire n_3108;
wire n_3053;
wire n_2988;
wire n_2987;
wire n_2984;
wire n_2985;
wire n_2982;
wire n_3050;
wire n_3041;
wire n_2989;
wire n_2983;
wire n_3051;
wire n_3045;
wire n_2986;
wire n_3048;
wire n_3046;
wire n_3052;
wire n_3043;
wire n_2996;
wire n_2995;
wire n_2992;
wire n_2993;
wire n_2990;
wire n_3036;
wire n_3027;
wire n_2997;
wire n_2991;
wire n_3037;
wire n_3031;
wire n_2994;
wire n_3034;
wire n_3032;
wire n_3038;
wire n_3029;
wire n_3025;
wire n_3004;
wire n_3003;
wire n_3002;
wire n_2999;
wire n_2998;
wire n_3015;
wire n_3022;
wire n_3011;
wire n_3005;
wire n_3000;
wire n_3001;
wire n_3021;
wire n_3012;
wire n_3023;
wire n_3019;
wire n_3017;
wire n_3024;
wire n_3013;
wire n_3009;
wire n_3006;
wire n_3238;
wire n_3243;
wire n_3242;
wire n_3008;
wire n_3007;
wire n_3240;
wire n_3241;
wire n_3239;
wire n_3010;
wire n_3014;
wire n_3018;
wire n_3020;
wire n_3016;
wire n_3026;
wire n_3030;
wire n_3033;
wire n_3028;
wire n_3035;
wire n_3040;
wire n_3044;
wire n_3047;
wire n_3042;
wire n_3049;
wire n_3075;
wire n_3054;
wire n_3082;
wire n_3061;
wire n_3103;
wire n_3093;
wire n_3057;
wire n_3101;
wire n_3096;
wire n_3059;
wire n_3062;
wire n_3065;
wire n_3104;
wire n_3071;
wire n_3115;
wire n_3110;
wire n_3073;
wire n_3092;
wire n_3078;
wire n_3090;
wire n_3085;
wire n_3080;
wire n_3126;
wire n_3144;
wire n_3154;
wire n_3155;
wire n_3165;
wire n_3122;
wire n_3180;
wire n_3175;
wire n_3124;
wire n_3167;
wire n_3129;
wire n_3173;
wire n_3128;
wire n_3134;
wire n_3163;
wire n_3158;
wire n_3136;
wire n_3140;
wire n_3152;
wire n_3147;
wire n_3142;
wire n_3184;
wire n_3188;
wire n_3191;
wire n_3186;
wire n_3193;
wire n_3198;
wire n_3202;
wire n_3205;
wire n_3200;
wire n_3207;
wire n_3212;
wire n_3216;
wire n_3219;
wire n_3214;
wire n_3221;
wire n_3237;
wire n_3227;
wire n_3234;
wire sgo__n3;
wire sgo__n5;
wire sgo__n208;
wire sgo__n10;
wire sgo__sro_n216;
wire sgo__n19;
wire sgo__sro_n217;
wire sgo__sro_n224;
wire sgo__sro_n225;
wire sgo__sro_n226;
wire sgo__sro_n227;
wire sgo__n43;
wire sgo__n78;
wire sgo__n98;
wire sgo__n99;
wire sgo__n109;
wire sgo__n122;
wire CLOCK_sgo__n358;
wire sgo__n134;
wire sgo__n141;
wire sgo__n147;
wire sgo__n148;
wire sgo__n150;
wire sgo__n162;
wire sgo__n164;
wire sgo__n168;
wire sgo__n170;
wire sgo__n172;
wire sgo__n174;
wire CLOCK_sgo__n359;
wire sgo__n176;
wire sgo__n177;
wire sgo__n178;
wire sgo__n180;
wire sgo__n182;
wire CLOCK_opt_ipo_n357;
wire sgo__n195;
wire sgo__n201;
wire sgo__n203;


INV_X4 i_2443 (.ZN (n_3309), .A (b[31]));
INV_X4 i_2442 (.ZN (n_3308), .A (b[30]));
INV_X8 i_2441 (.ZN (n_3307), .A (b[29]));
INV_X8 i_2440 (.ZN (n_3306), .A (b[28]));
INV_X4 i_2439 (.ZN (n_3305), .A (b[27]));
INV_X4 i_2438 (.ZN (n_3304), .A (b[26]));
INV_X4 i_2437 (.ZN (n_3303), .A (b[25]));
INV_X8 i_2436 (.ZN (n_3302), .A (b[24]));
INV_X4 i_2435 (.ZN (n_3301), .A (b[23]));
INV_X4 i_2434 (.ZN (n_3300), .A (b[22]));
INV_X4 i_2433 (.ZN (n_3299), .A (b[21]));
INV_X2 i_2432 (.ZN (n_3298), .A (b[20]));
INV_X2 i_2431 (.ZN (n_3297), .A (b[19]));
INV_X2 i_2430 (.ZN (n_3296), .A (b[18]));
INV_X2 i_2429 (.ZN (n_3295), .A (b[17]));
INV_X4 i_2428 (.ZN (n_3294), .A (b[16]));
INV_X4 i_2427 (.ZN (n_3293), .A (b[15]));
INV_X2 i_2426 (.ZN (n_3292), .A (b[14]));
INV_X4 i_2425 (.ZN (n_3291), .A (b[13]));
INV_X2 i_2424 (.ZN (n_3290), .A (b[12]));
INV_X4 i_2423 (.ZN (n_3289), .A (b[11]));
INV_X2 i_2422 (.ZN (n_3288), .A (b[10]));
INV_X2 i_2421 (.ZN (n_3287), .A (b[9]));
INV_X4 i_2420 (.ZN (n_3286), .A (b[8]));
INV_X4 i_2419 (.ZN (n_3285), .A (b[7]));
INV_X2 i_2418 (.ZN (n_3284), .A (b[6]));
INV_X4 i_2417 (.ZN (n_3283), .A (b[5]));
INV_X4 i_2416 (.ZN (n_3282), .A (b[4]));
INV_X4 i_2415 (.ZN (n_3281), .A (b[3]));
INV_X4 i_2414 (.ZN (n_3280), .A (b[2]));
INV_X4 i_2413 (.ZN (n_3279), .A (b[1]));
INV_X4 i_2412 (.ZN (n_3278), .A (b[0]));
INV_X2 i_2411 (.ZN (n_3277), .A (a[31]));
INV_X2 i_2410 (.ZN (n_3276), .A (a[30]));
INV_X2 i_2409 (.ZN (n_3275), .A (a[29]));
INV_X4 i_2408 (.ZN (n_3274), .A (a[28]));
INV_X4 i_2407 (.ZN (n_3273), .A (a[27]));
INV_X2 i_2406 (.ZN (n_3272), .A (a[26]));
INV_X4 i_2405 (.ZN (n_3271), .A (a[25]));
INV_X2 i_2404 (.ZN (n_3270), .A (a[24]));
INV_X4 i_2403 (.ZN (n_3269), .A (a[23]));
INV_X4 i_2402 (.ZN (n_3268), .A (a[22]));
INV_X4 i_2401 (.ZN (n_3267), .A (a[21]));
INV_X4 i_2400 (.ZN (n_3266), .A (a[20]));
INV_X4 i_2399 (.ZN (n_3265), .A (a[19]));
INV_X2 i_2398 (.ZN (n_3264), .A (a[18]));
INV_X2 i_2397 (.ZN (n_3263), .A (a[17]));
INV_X4 i_2396 (.ZN (n_3262), .A (a[16]));
INV_X4 i_2395 (.ZN (n_3261), .A (a[15]));
INV_X2 i_2394 (.ZN (n_3260), .A (a[14]));
INV_X4 i_2393 (.ZN (n_3259), .A (a[13]));
INV_X4 i_2392 (.ZN (n_3258), .A (a[12]));
INV_X2 i_2391 (.ZN (n_3257), .A (a[11]));
INV_X4 i_2390 (.ZN (n_3256), .A (a[10]));
INV_X4 i_2389 (.ZN (n_3255), .A (a[9]));
INV_X4 i_2388 (.ZN (n_3254), .A (a[8]));
INV_X2 i_2387 (.ZN (n_3253), .A (a[7]));
INV_X2 i_2386 (.ZN (n_3252), .A (a[6]));
INV_X2 i_2385 (.ZN (n_3251), .A (a[5]));
INV_X2 i_2384 (.ZN (n_3250), .A (a[4]));
INV_X2 i_2383 (.ZN (n_3249), .A (a[3]));
INV_X2 i_2382 (.ZN (n_3248), .A (a[2]));
INV_X2 i_2381 (.ZN (n_3247), .A (a[1]));
INV_X2 i_2380 (.ZN (n_3246), .A (a[0]));
INV_X1 i_2379 (.ZN (n_3245), .A (n_929));
INV_X1 i_2378 (.ZN (n_3244), .A (n_988));
INV_X1 i_2377 (.ZN (n_3243), .A (n_1857));
INV_X1 i_2376 (.ZN (n_3242), .A (n_1858));
NOR2_X1 i_2375 (.ZN (n_3241), .A1 (n_3309), .A2 (n_3277));
NOR2_X1 i_2374 (.ZN (n_3240), .A1 (n_1859), .A2 (n_3241));
NAND2_X1 i_2373 (.ZN (n_3239), .A1 (n_1859), .A2 (n_3241));
NOR2_X1 i_2372 (.ZN (n_3238), .A1 (n_3243), .A2 (n_3242));
AND2_X1 i_2371 (.ZN (n_3237), .A1 (n_6), .A2 (n_10));
NAND2_X1 i_2370 (.ZN (n_3236), .A1 (n_2), .A2 (n_4));
NOR2_X1 i_2369 (.ZN (n_3235), .A1 (n_3278), .A2 (n_3248));
NOR2_X1 i_2368 (.ZN (n_3234), .A1 (n_0), .A2 (n_3235));
NOR2_X1 i_2367 (.ZN (n_3233), .A1 (n_3279), .A2 (n_3246));
NOR2_X1 i_2366 (.ZN (n_3232), .A1 (n_3278), .A2 (n_3247));
NOR2_X1 i_2365 (.ZN (p_0[0]), .A1 (n_3278), .A2 (n_3246));
NOR2_X1 i_2364 (.ZN (n_3231), .A1 (n_3279), .A2 (n_3247));
NAND2_X1 i_2363 (.ZN (n_3230), .A1 (p_0[0]), .A2 (n_3231));
NAND2_X1 i_2362 (.ZN (n_3229), .A1 (n_0), .A2 (n_3235));
AOI21_X1 i_2361 (.ZN (n_3228), .A (n_3234), .B1 (n_3230), .B2 (n_3229));
OAI21_X1 i_2360 (.ZN (n_3227), .A (n_3228), .B1 (n_2), .B2 (n_4));
NAND2_X1 i_2359 (.ZN (n_3226), .A1 (n_3236), .A2 (n_3227));
OAI22_X1 i_2358 (.ZN (n_3225), .A1 (n_6), .A2 (n_10), .B1 (n_3237), .B2 (n_3226));
NOR2_X1 i_2357 (.ZN (n_3224), .A1 (n_52), .A2 (n_54));
NOR2_X1 i_2356 (.ZN (n_3223), .A1 (n_26), .A2 (n_28));
NOR2_X1 i_2355 (.ZN (n_3222), .A1 (n_38), .A2 (n_40));
OR3_X1 i_2354 (.ZN (n_3221), .A1 (n_3224), .A2 (n_3222), .A3 (n_3223));
NOR2_X1 i_2353 (.ZN (n_3220), .A1 (n_16), .A2 (n_18));
NOR3_X1 i_2352 (.ZN (n_3219), .A1 (n_3221), .A2 (n_3220), .A3 (n_3225));
NAND2_X1 i_2351 (.ZN (n_3218), .A1 (n_16), .A2 (n_18));
NAND2_X1 i_2350 (.ZN (n_3217), .A1 (n_26), .A2 (n_28));
AOI21_X1 i_2349 (.ZN (n_3216), .A (n_3221), .B1 (n_3218), .B2 (n_3217));
AND2_X1 i_2348 (.ZN (n_3215), .A1 (n_52), .A2 (n_54));
NAND2_X1 i_2347 (.ZN (n_3214), .A1 (n_38), .A2 (n_40));
INV_X1 i_2346 (.ZN (n_3213), .A (n_3214));
NOR2_X1 i_2345 (.ZN (n_3212), .A1 (n_3224), .A2 (n_3214));
NOR4_X1 i_2344 (.ZN (n_3211), .A1 (n_3215), .A2 (n_3212), .A3 (n_3216), .A4 (n_3219));
NOR2_X1 i_2343 (.ZN (n_3210), .A1 (n_128), .A2 (n_130));
NOR2_X1 i_2342 (.ZN (n_3209), .A1 (n_86), .A2 (n_88));
NOR2_X1 i_2341 (.ZN (n_3208), .A1 (n_106), .A2 (n_108));
OR3_X1 i_2340 (.ZN (n_3207), .A1 (n_3210), .A2 (n_3208), .A3 (n_3209));
NOR2_X1 i_2339 (.ZN (n_3206), .A1 (n_68), .A2 (n_70));
NOR3_X1 i_2338 (.ZN (n_3205), .A1 (n_3207), .A2 (n_3206), .A3 (n_3211));
NAND2_X1 i_2337 (.ZN (n_3204), .A1 (n_68), .A2 (n_70));
NAND2_X1 i_2336 (.ZN (n_3203), .A1 (n_86), .A2 (n_88));
AOI21_X1 i_2335 (.ZN (n_3202), .A (n_3207), .B1 (n_3204), .B2 (n_3203));
AND2_X1 i_2334 (.ZN (n_3201), .A1 (n_128), .A2 (n_130));
NAND2_X1 i_2333 (.ZN (n_3200), .A1 (n_106), .A2 (n_108));
INV_X1 i_2332 (.ZN (n_3199), .A (n_3200));
NOR2_X1 i_2331 (.ZN (n_3198), .A1 (n_3210), .A2 (n_3200));
NOR4_X1 i_2330 (.ZN (n_3197), .A1 (n_3201), .A2 (n_3198), .A3 (n_3202), .A4 (n_3205));
NOR2_X1 i_2329 (.ZN (n_3196), .A1 (n_236), .A2 (n_238));
NOR2_X1 i_2328 (.ZN (n_3195), .A1 (n_178), .A2 (n_180));
NOR2_X1 i_2327 (.ZN (n_3194), .A1 (n_206), .A2 (n_208));
OR3_X1 i_2326 (.ZN (n_3193), .A1 (n_3196), .A2 (n_3194), .A3 (n_3195));
NOR2_X1 i_2325 (.ZN (n_3192), .A1 (n_152), .A2 (n_154));
NOR3_X1 i_2324 (.ZN (n_3191), .A1 (n_3193), .A2 (n_3192), .A3 (n_3197));
NAND2_X1 i_2323 (.ZN (n_3190), .A1 (n_152), .A2 (n_154));
NAND2_X1 i_2322 (.ZN (n_3189), .A1 (n_178), .A2 (n_180));
AOI21_X1 i_2321 (.ZN (n_3188), .A (n_3193), .B1 (n_3190), .B2 (n_3189));
AND2_X1 i_2320 (.ZN (n_3187), .A1 (n_236), .A2 (n_238));
NAND2_X1 i_2319 (.ZN (n_3186), .A1 (n_206), .A2 (n_208));
INV_X1 i_2318 (.ZN (n_3185), .A (n_3186));
NOR2_X1 i_2317 (.ZN (n_3184), .A1 (n_3196), .A2 (n_3186));
NOR4_X4 i_2316 (.ZN (n_3183), .A1 (n_3187), .A2 (n_3184), .A3 (n_3188), .A4 (n_3191));
NOR2_X1 i_2315 (.ZN (n_3182), .A1 (n_379), .A2 (n_418));
NOR2_X1 i_2314 (.ZN (n_3181), .A1 (n_505), .A2 (n_550));
INV_X1 i_2313 (.ZN (n_3180), .A (n_3181));
NOR2_X1 i_2312 (.ZN (n_3179), .A1 (n_419), .A2 (n_460));
INV_X1 i_2311 (.ZN (n_3178), .A (n_3179));
NOR2_X1 i_2310 (.ZN (n_3177), .A1 (n_461), .A2 (n_504));
INV_X1 i_2309 (.ZN (n_3176), .A (n_3177));
NAND3_X1 i_2308 (.ZN (n_3175), .A1 (n_3180), .A2 (n_3176), .A3 (n_3178));
OR2_X2 i_2307 (.ZN (n_3174), .A1 (n_3182), .A2 (n_3175));
NOR2_X2 i_2306 (.ZN (n_3173), .A1 (n_929), .A2 (n_988));
INV_X1 i_2305 (.ZN (n_3172), .A (n_3173));
NOR2_X1 i_2304 (.ZN (n_3171), .A1 (n_811), .A2 (n_868));
INV_X1 i_2303 (.ZN (n_3170), .A (n_3171));
NOR2_X1 i_2302 (.ZN (n_3169), .A1 (n_869), .A2 (n_928));
INV_X1 i_2301 (.ZN (n_3168), .A (n_3169));
NAND3_X1 i_2300 (.ZN (n_3167), .A1 (n_3172), .A2 (n_3168), .A3 (n_3170));
NOR2_X1 i_2299 (.ZN (n_3166), .A1 (n_755), .A2 (n_810));
OR2_X2 i_2298 (.ZN (n_3165), .A1 (n_3167), .A2 (n_3166));
NOR2_X1 i_2297 (.ZN (n_3164), .A1 (n_701), .A2 (n_754));
INV_X1 i_2296 (.ZN (n_3163), .A (n_3164));
NOR2_X1 i_2295 (.ZN (n_3162), .A1 (n_599), .A2 (n_648));
INV_X1 i_2294 (.ZN (n_3161), .A (n_3162));
NOR2_X1 i_2293 (.ZN (n_3160), .A1 (n_649), .A2 (n_700));
INV_X1 i_2292 (.ZN (n_3159), .A (n_3160));
NAND3_X1 i_2291 (.ZN (n_3158), .A1 (n_3163), .A2 (n_3159), .A3 (n_3161));
NOR2_X1 i_2290 (.ZN (n_3157), .A1 (n_596), .A2 (n_598));
OR2_X1 i_2289 (.ZN (n_3156), .A1 (n_3158), .A2 (n_3157));
OR2_X2 i_2288 (.ZN (n_3155), .A1 (n_3165), .A2 (n_3156));
OR2_X1 i_2287 (.ZN (n_3154), .A1 (n_3174), .A2 (n_3155));
NOR2_X1 i_2286 (.ZN (n_3153), .A1 (n_376), .A2 (n_378));
INV_X1 i_2285 (.ZN (n_3152), .A (n_3153));
NOR2_X1 i_2284 (.ZN (n_3151), .A1 (n_271), .A2 (n_304));
INV_X1 i_2283 (.ZN (n_3150), .A (n_3151));
NOR2_X1 i_2282 (.ZN (n_3149), .A1 (n_305), .A2 (n_340));
INV_X1 i_2281 (.ZN (n_3148), .A (n_3149));
NAND3_X1 i_2280 (.ZN (n_3147), .A1 (n_3152), .A2 (n_3148), .A3 (n_3150));
NOR2_X1 i_2279 (.ZN (n_3146), .A1 (n_268), .A2 (n_270));
OR2_X1 i_2278 (.ZN (n_3145), .A1 (n_3147), .A2 (n_3146));
NOR3_X1 i_2277 (.ZN (n_3144), .A1 (n_3154), .A2 (n_3145), .A3 (n_3183));
NAND2_X1 i_2276 (.ZN (n_3143), .A1 (n_268), .A2 (n_270));
NAND2_X1 i_2275 (.ZN (n_3142), .A1 (n_271), .A2 (n_304));
INV_X1 i_2274 (.ZN (n_3141), .A (n_3142));
AOI21_X1 i_2273 (.ZN (n_3140), .A (n_3147), .B1 (n_3143), .B2 (n_3142));
AND2_X1 i_2272 (.ZN (n_3139), .A1 (n_305), .A2 (n_340));
AOI221_X2 i_2271 (.ZN (n_3138), .A (n_3140), .B1 (n_376), .B2 (n_378), .C1 (n_3152), .C2 (n_3139));
NAND2_X1 i_2270 (.ZN (n_3137), .A1 (n_596), .A2 (n_598));
NAND2_X1 i_2269 (.ZN (n_3136), .A1 (n_599), .A2 (n_648));
INV_X1 i_2268 (.ZN (n_3135), .A (n_3136));
AOI21_X1 i_2267 (.ZN (n_3134), .A (n_3158), .B1 (n_3137), .B2 (n_3136));
AND2_X1 i_2266 (.ZN (n_3133), .A1 (n_649), .A2 (n_700));
AOI221_X1 i_2265 (.ZN (n_3132), .A (n_3134), .B1 (n_701), .B2 (n_754), .C1 (n_3163), .C2 (n_3133));
NAND2_X1 i_2264 (.ZN (n_3131), .A1 (n_755), .A2 (n_810));
AND2_X1 i_2263 (.ZN (n_3130), .A1 (n_811), .A2 (n_868));
AOI21_X1 i_2262 (.ZN (n_3129), .A (n_3130), .B1 (n_755), .B2 (n_810));
NAND2_X1 i_2261 (.ZN (n_3128), .A1 (n_869), .A2 (n_928));
INV_X1 i_2260 (.ZN (n_3127), .A (n_3128));
OAI222_X1 i_2259 (.ZN (n_3126), .A1 (n_3167), .A2 (n_3129), .B1 (n_3173), .B2 (n_3128)
    , .C1 (n_3245), .C2 (n_3244));
NAND2_X1 i_2258 (.ZN (n_3125), .A1 (n_379), .A2 (n_418));
NAND2_X1 i_2257 (.ZN (n_3124), .A1 (n_419), .A2 (n_460));
INV_X1 i_2256 (.ZN (n_3123), .A (n_3124));
AOI21_X1 i_2255 (.ZN (n_3122), .A (n_3175), .B1 (n_3125), .B2 (n_3124));
AND2_X1 i_2254 (.ZN (n_3121), .A1 (n_461), .A2 (n_504));
AOI221_X2 i_2253 (.ZN (n_3120), .A (n_3122), .B1 (n_505), .B2 (n_550), .C1 (n_3180), .C2 (n_3121));
NOR3_X2 i_2251 (.ZN (n_3118), .A1 (n_3126), .A2 (sgo__sro_n216), .A3 (n_3144));
NOR2_X1 i_2250 (.ZN (n_3117), .A1 (n_1209), .A2 (n_1258));
NOR2_X1 i_2249 (.ZN (n_3116), .A1 (n_1353), .A2 (n_1396));
INV_X1 i_2248 (.ZN (n_3115), .A (n_3116));
NOR2_X1 i_2247 (.ZN (n_3114), .A1 (n_1259), .A2 (n_1306));
INV_X1 i_2246 (.ZN (n_3113), .A (n_3114));
NOR2_X1 i_2245 (.ZN (n_3112), .A1 (n_1307), .A2 (n_1352));
INV_X1 i_2244 (.ZN (n_3111), .A (n_3112));
NAND3_X1 i_2243 (.ZN (n_3110), .A1 (n_3115), .A2 (n_3111), .A3 (n_3113));
OR2_X1 i_2242 (.ZN (n_3109), .A1 (n_3117), .A2 (n_3110));
NOR2_X1 i_2241 (.ZN (n_3108), .A1 (n_1649), .A2 (n_1676));
NOR2_X1 i_2240 (.ZN (n_3107), .A1 (n_1587), .A2 (n_1618));
NOR2_X1 i_2239 (.ZN (n_3106), .A1 (n_1619), .A2 (n_1648));
NOR2_X1 i_2238 (.ZN (n_3105), .A1 (n_3107), .A2 (n_3106));
NOR3_X1 i_2237 (.ZN (n_3104), .A1 (n_3108), .A2 (n_3106), .A3 (n_3107));
OAI21_X1 i_2236 (.ZN (n_3103), .A (n_3104), .B1 (n_1553), .B2 (n_1586));
NOR2_X1 i_2235 (.ZN (n_3102), .A1 (n_1517), .A2 (n_1552));
INV_X1 i_2234 (.ZN (n_3101), .A (n_3102));
NOR2_X1 i_2233 (.ZN (n_3100), .A1 (n_1439), .A2 (n_1478));
INV_X1 i_2232 (.ZN (n_3099), .A (n_3100));
NOR2_X1 i_2231 (.ZN (n_3098), .A1 (n_1479), .A2 (n_1516));
INV_X1 i_2230 (.ZN (n_3097), .A (n_3098));
NAND3_X1 i_2229 (.ZN (n_3096), .A1 (n_3101), .A2 (n_3097), .A3 (n_3099));
NOR2_X1 i_2228 (.ZN (n_3095), .A1 (n_1397), .A2 (n_1438));
OR2_X1 i_2227 (.ZN (n_3094), .A1 (n_3096), .A2 (n_3095));
OR2_X1 i_2226 (.ZN (n_3093), .A1 (n_3103), .A2 (n_3094));
OR2_X4 i_2225 (.ZN (n_3092), .A1 (n_3109), .A2 (n_3093));
NOR2_X1 i_2224 (.ZN (n_3091), .A1 (n_1157), .A2 (n_1208));
INV_X1 i_2223 (.ZN (n_3090), .A (n_3091));
NOR2_X1 i_2222 (.ZN (n_3089), .A1 (n_1047), .A2 (n_1102));
INV_X1 i_2221 (.ZN (n_3088), .A (n_3089));
NOR2_X1 i_2220 (.ZN (n_3087), .A1 (n_1103), .A2 (n_1156));
INV_X1 i_2219 (.ZN (n_3086), .A (n_3087));
NAND3_X1 i_2218 (.ZN (n_3085), .A1 (n_3090), .A2 (n_3086), .A3 (n_3088));
NOR2_X1 i_2217 (.ZN (n_3084), .A1 (n_989), .A2 (n_1046));
OR2_X2 i_2216 (.ZN (n_3083), .A1 (n_3085), .A2 (n_3084));
NOR3_X2 i_2215 (.ZN (n_3082), .A1 (n_3092), .A2 (n_3083), .A3 (sgo__n208));
NAND2_X1 i_2214 (.ZN (n_3081), .A1 (n_989), .A2 (n_1046));
NAND2_X1 i_2213 (.ZN (n_3080), .A1 (n_1047), .A2 (n_1102));
INV_X1 i_2212 (.ZN (n_3079), .A (n_3080));
AOI21_X1 i_2211 (.ZN (n_3078), .A (n_3085), .B1 (n_3081), .B2 (n_3080));
AND2_X1 i_2210 (.ZN (n_3077), .A1 (n_1103), .A2 (n_1156));
AOI221_X1 i_2209 (.ZN (n_3076), .A (n_3078), .B1 (n_1157), .B2 (n_1208), .C1 (n_3090), .C2 (n_3077));
NOR2_X4 i_2208 (.ZN (n_3075), .A1 (n_3092), .A2 (n_3076));
NAND2_X1 i_2207 (.ZN (n_3074), .A1 (n_1209), .A2 (n_1258));
NAND2_X1 i_2206 (.ZN (n_3073), .A1 (n_1259), .A2 (n_1306));
INV_X1 i_2205 (.ZN (n_3072), .A (n_3073));
AOI21_X1 i_2204 (.ZN (n_3071), .A (n_3110), .B1 (n_3074), .B2 (n_3073));
AND2_X1 i_2203 (.ZN (n_3070), .A1 (n_1307), .A2 (n_1352));
AOI221_X1 i_2202 (.ZN (n_3069), .A (n_3071), .B1 (n_1353), .B2 (n_1396), .C1 (n_3115), .C2 (n_3070));
NAND2_X1 i_2201 (.ZN (n_3068), .A1 (n_1553), .A2 (n_1586));
INV_X1 i_2200 (.ZN (n_3067), .A (n_3068));
AND2_X1 i_2199 (.ZN (n_3066), .A1 (n_1587), .A2 (n_1618));
OAI21_X1 i_2198 (.ZN (n_3065), .A (n_3104), .B1 (n_3067), .B2 (n_3066));
NAND2_X1 i_2197 (.ZN (n_3064), .A1 (n_1619), .A2 (n_1648));
INV_X1 i_2196 (.ZN (n_3063), .A (n_3064));
OAI21_X1 i_2195 (.ZN (n_3062), .A (n_3065), .B1 (n_3108), .B2 (n_3064));
AOI21_X1 i_2194 (.ZN (n_3061), .A (n_3062), .B1 (n_1649), .B2 (n_1676));
NAND2_X1 i_2193 (.ZN (n_3060), .A1 (n_1397), .A2 (n_1438));
NAND2_X1 i_2192 (.ZN (n_3059), .A1 (n_1439), .A2 (n_1478));
INV_X1 i_2191 (.ZN (n_3058), .A (n_3059));
AOI21_X1 i_2190 (.ZN (n_3057), .A (n_3096), .B1 (n_3060), .B2 (n_3059));
AND2_X1 i_2189 (.ZN (n_3056), .A1 (n_1479), .A2 (n_1516));
AOI221_X1 i_2188 (.ZN (n_3055), .A (n_3057), .B1 (n_1517), .B2 (n_1552), .C1 (n_3101), .C2 (n_3056));
OAI221_X1 i_2187 (.ZN (n_3054), .A (n_3061), .B1 (n_3103), .B2 (n_3055), .C1 (n_3093), .C2 (n_3069));
NOR3_X4 i_2186 (.ZN (n_3053), .A1 (n_3075), .A2 (CLOCK_opt_ipo_n357), .A3 (n_3082));
NOR2_X1 i_2185 (.ZN (n_3052), .A1 (n_1749), .A2 (n_1768));
NOR2_X1 i_2184 (.ZN (n_3051), .A1 (n_1703), .A2 (n_1726));
NOR2_X1 i_2183 (.ZN (n_3050), .A1 (n_1727), .A2 (n_1748));
OR3_X1 i_2182 (.ZN (n_3049), .A1 (n_3052), .A2 (n_3050), .A3 (n_3051));
NOR2_X1 i_2181 (.ZN (n_3048), .A1 (n_1677), .A2 (n_1702));
NOR3_X1 i_2180 (.ZN (n_3047), .A1 (n_3049), .A2 (n_3048), .A3 (n_3053));
NAND2_X1 i_2179 (.ZN (n_3046), .A1 (n_1677), .A2 (n_1702));
NAND2_X1 i_2178 (.ZN (n_3045), .A1 (n_1703), .A2 (n_1726));
AOI21_X1 i_2177 (.ZN (n_3044), .A (n_3049), .B1 (n_3046), .B2 (n_3045));
AND2_X1 i_2176 (.ZN (n_3043), .A1 (n_1749), .A2 (n_1768));
NAND2_X1 i_2175 (.ZN (n_3042), .A1 (n_1727), .A2 (n_1748));
INV_X1 i_2174 (.ZN (n_3041), .A (n_3042));
NOR2_X1 i_2173 (.ZN (n_3040), .A1 (n_3052), .A2 (n_3042));
NOR2_X1 i_2171 (.ZN (n_3038), .A1 (n_1817), .A2 (n_1828));
NOR2_X1 i_2170 (.ZN (n_3037), .A1 (n_1787), .A2 (n_1802));
NOR2_X1 i_2169 (.ZN (n_3036), .A1 (n_1803), .A2 (n_1816));
OR3_X1 i_2168 (.ZN (n_3035), .A1 (n_3038), .A2 (n_3036), .A3 (n_3037));
NOR2_X1 i_2167 (.ZN (n_3034), .A1 (n_1769), .A2 (n_1786));
NOR3_X1 i_2166 (.ZN (n_3033), .A1 (n_3035), .A2 (n_3034), .A3 (sgo__sro_n224));
NAND2_X1 i_2165 (.ZN (n_3032), .A1 (n_1769), .A2 (n_1786));
NAND2_X1 i_2164 (.ZN (n_3031), .A1 (n_1787), .A2 (n_1802));
AOI21_X1 i_2163 (.ZN (n_3030), .A (n_3035), .B1 (n_3032), .B2 (n_3031));
AND2_X1 i_2162 (.ZN (n_3029), .A1 (n_1817), .A2 (n_1828));
NAND2_X1 i_2161 (.ZN (n_3028), .A1 (n_1803), .A2 (n_1816));
INV_X1 i_2160 (.ZN (n_3027), .A (n_3028));
NOR2_X1 i_2159 (.ZN (n_3026), .A1 (n_3038), .A2 (n_3028));
NOR4_X2 i_2158 (.ZN (n_3025), .A1 (n_3029), .A2 (n_3026), .A3 (n_3030), .A4 (n_3033));
NOR2_X1 i_2157 (.ZN (n_3024), .A1 (n_1853), .A2 (n_1856));
NOR2_X1 i_2156 (.ZN (n_3023), .A1 (n_1839), .A2 (n_1846));
NOR2_X1 i_2155 (.ZN (n_3022), .A1 (n_1847), .A2 (n_1852));
NOR2_X1 i_2154 (.ZN (n_3021), .A1 (n_3023), .A2 (n_3022));
OAI21_X1 i_2153 (.ZN (n_3020), .A (n_3021), .B1 (n_1853), .B2 (n_1856));
NOR2_X1 i_2152 (.ZN (n_3019), .A1 (n_1829), .A2 (n_1838));
NOR3_X1 i_2151 (.ZN (n_3018), .A1 (n_3020), .A2 (n_3019), .A3 (n_3025));
NAND2_X1 i_2150 (.ZN (n_3017), .A1 (n_1829), .A2 (n_1838));
NAND2_X1 i_2149 (.ZN (n_3016), .A1 (n_1839), .A2 (n_1846));
INV_X1 i_2148 (.ZN (n_3015), .A (n_3016));
AOI21_X1 i_2147 (.ZN (n_3014), .A (n_3020), .B1 (n_3017), .B2 (n_3016));
AND2_X1 i_2146 (.ZN (n_3013), .A1 (n_1853), .A2 (n_1856));
NAND2_X1 i_2145 (.ZN (n_3012), .A1 (n_1847), .A2 (n_1852));
INV_X1 i_2144 (.ZN (n_3011), .A (n_3012));
NOR2_X1 i_2143 (.ZN (n_3010), .A1 (n_3024), .A2 (n_3012));
OR4_X2 i_2142 (.ZN (n_3009), .A1 (n_3013), .A2 (n_3010), .A3 (n_3014), .A4 (n_3018));
OAI22_X2 i_2141 (.ZN (n_3008), .A1 (n_1857), .A2 (n_1858), .B1 (n_3238), .B2 (n_3009));
AOI21_X1 i_2140 (.ZN (p_0[63]), .A (n_3240), .B1 (n_3239), .B2 (n_3008));
AOI21_X1 i_2139 (.ZN (n_3007), .A (n_3240), .B1 (n_1859), .B2 (n_3241));
XNOR2_X1 i_2138 (.ZN (p_0[62]), .A (n_3008), .B (n_3007));
AOI21_X1 i_2137 (.ZN (n_3006), .A (n_3238), .B1 (n_3243), .B2 (n_3242));
XOR2_X1 i_2136 (.Z (p_0[61]), .A (n_3009), .B (n_3006));
NOR2_X1 i_2135 (.ZN (n_3005), .A1 (n_3024), .A2 (n_3013));
OAI21_X1 i_2134 (.ZN (n_3004), .A (n_3017), .B1 (n_1829), .B2 (n_1838));
AOI21_X1 i_2133 (.ZN (n_3003), .A (n_3019), .B1 (n_3025), .B2 (n_3017));
NOR2_X1 i_2132 (.ZN (n_3002), .A1 (n_3023), .A2 (n_3015));
NAND2_X1 i_2131 (.ZN (n_3001), .A1 (n_3012), .A2 (n_3002));
OAI22_X1 i_2130 (.ZN (n_3000), .A1 (n_3003), .A2 (n_3001), .B1 (n_3021), .B2 (n_3011));
XNOR2_X1 i_2129 (.ZN (p_0[60]), .A (n_3005), .B (n_3000));
NOR2_X1 i_2128 (.ZN (n_2999), .A1 (n_3022), .A2 (n_3011));
OAI22_X1 i_2127 (.ZN (n_2998), .A1 (n_1839), .A2 (n_1846), .B1 (n_3015), .B2 (n_3003));
XNOR2_X1 i_2126 (.ZN (p_0[59]), .A (n_2999), .B (n_2998));
XOR2_X1 i_2125 (.Z (p_0[58]), .A (n_3003), .B (n_3002));
XOR2_X1 i_2124 (.Z (p_0[57]), .A (n_3025), .B (n_3004));
NOR2_X1 i_2123 (.ZN (n_2997), .A1 (n_3038), .A2 (n_3029));
OAI21_X1 i_2122 (.ZN (n_2996), .A (n_3032), .B1 (n_1769), .B2 (n_1786));
AOI21_X1 i_2121 (.ZN (n_2995), .A (n_3034), .B1 (sgo__sro_n224), .B2 (n_3032));
INV_X1 i_2120 (.ZN (n_2994), .A (n_2995));
AOI21_X1 i_2119 (.ZN (n_2993), .A (n_3037), .B1 (n_3031), .B2 (n_2994));
AOI21_X1 i_2118 (.ZN (n_2992), .A (n_3037), .B1 (n_1787), .B2 (n_1802));
OAI22_X1 i_2117 (.ZN (n_2991), .A1 (n_1803), .A2 (n_1816), .B1 (n_3027), .B2 (n_2993));
XNOR2_X1 i_2116 (.ZN (p_0[56]), .A (n_2997), .B (n_2991));
NOR2_X1 i_2115 (.ZN (n_2990), .A1 (n_3036), .A2 (n_3027));
XOR2_X1 i_2114 (.Z (p_0[55]), .A (n_2993), .B (n_2990));
XOR2_X1 i_2113 (.Z (p_0[54]), .A (n_2995), .B (n_2992));
XOR2_X1 i_2112 (.Z (p_0[53]), .A (sgo__sro_n224), .B (n_2996));
NOR2_X1 i_2111 (.ZN (n_2989), .A1 (n_3052), .A2 (n_3043));
OAI21_X1 i_2110 (.ZN (n_2988), .A (n_3046), .B1 (n_1677), .B2 (n_1702));
AOI21_X1 i_2109 (.ZN (n_2987), .A (n_3048), .B1 (n_3053), .B2 (n_3046));
INV_X1 i_2108 (.ZN (n_2986), .A (n_2987));
AOI21_X1 i_2107 (.ZN (n_2985), .A (n_3051), .B1 (n_3045), .B2 (n_2986));
AOI21_X1 i_2106 (.ZN (n_2984), .A (n_3051), .B1 (n_1703), .B2 (n_1726));
OAI22_X1 i_2105 (.ZN (n_2983), .A1 (n_1727), .A2 (n_1748), .B1 (n_3041), .B2 (n_2985));
XNOR2_X1 i_2104 (.ZN (p_0[52]), .A (n_2989), .B (n_2983));
NOR2_X1 i_2103 (.ZN (n_2982), .A1 (n_3050), .A2 (n_3041));
XOR2_X1 i_2102 (.Z (p_0[51]), .A (n_2985), .B (n_2982));
XOR2_X1 i_2101 (.Z (p_0[50]), .A (n_2987), .B (n_2984));
XOR2_X1 i_2100 (.Z (p_0[49]), .A (n_3053), .B (n_2988));
AOI21_X1 i_2099 (.ZN (n_2981), .A (n_3108), .B1 (n_1649), .B2 (n_1676));
OAI21_X1 i_2098 (.ZN (n_2980), .A (n_3076), .B1 (sgo__n208), .B2 (n_3083));
INV_X4 i_2097 (.ZN (n_2979), .A (n_2980));
OAI21_X1 i_2096 (.ZN (n_2978), .A (n_3069), .B1 (n_3109), .B2 (n_2979));
INV_X1 i_2095 (.ZN (n_2977), .A (n_2978));
OAI21_X1 i_2094 (.ZN (n_2976), .A (n_3055), .B1 (n_3094), .B2 (n_2977));
OAI21_X1 i_2093 (.ZN (n_2975), .A (n_3068), .B1 (n_1553), .B2 (n_1586));
OAI22_X1 i_2092 (.ZN (n_2974), .A1 (n_1553), .A2 (n_1586), .B1 (n_3067), .B2 (n_2976));
INV_X1 i_2091 (.ZN (n_2973), .A (n_2974));
NOR2_X1 i_2090 (.ZN (n_2972), .A1 (n_3107), .A2 (n_3066));
NAND3_X1 i_2089 (.ZN (n_2971), .A1 (n_3064), .A2 (n_2972), .A3 (n_2974));
OAI21_X1 i_2088 (.ZN (n_2970), .A (n_2971), .B1 (n_3105), .B2 (n_3063));
XNOR2_X1 i_2087 (.ZN (p_0[48]), .A (n_2981), .B (n_2970));
NOR2_X1 i_2086 (.ZN (n_2969), .A1 (n_3106), .A2 (n_3063));
OAI22_X1 i_2085 (.ZN (n_2968), .A1 (n_1587), .A2 (n_1618), .B1 (n_3066), .B2 (n_2973));
XNOR2_X1 i_2084 (.ZN (p_0[47]), .A (n_2969), .B (n_2968));
XOR2_X1 i_2083 (.Z (p_0[46]), .A (n_2973), .B (n_2972));
XNOR2_X1 i_2082 (.ZN (p_0[45]), .A (n_2976), .B (n_2975));
AOI21_X1 i_2081 (.ZN (n_2967), .A (n_3102), .B1 (n_1517), .B2 (n_1552));
OAI21_X1 i_2080 (.ZN (n_2966), .A (n_3060), .B1 (n_1397), .B2 (n_1438));
AOI21_X1 i_2079 (.ZN (n_2965), .A (n_3095), .B1 (n_3060), .B2 (n_2977));
OAI21_X1 i_2078 (.ZN (n_2964), .A (n_3099), .B1 (n_3058), .B2 (n_2965));
INV_X1 i_2077 (.ZN (n_2963), .A (n_2964));
NOR2_X1 i_2076 (.ZN (n_2962), .A1 (n_3100), .A2 (n_3058));
OAI21_X1 i_2075 (.ZN (n_2961), .A (n_3097), .B1 (n_3056), .B2 (n_2963));
XNOR2_X1 i_2074 (.ZN (p_0[44]), .A (n_2967), .B (n_2961));
NOR2_X1 i_2073 (.ZN (n_2960), .A1 (n_3098), .A2 (n_3056));
XOR2_X1 i_2072 (.Z (p_0[43]), .A (n_2963), .B (n_2960));
XOR2_X1 i_2071 (.Z (p_0[42]), .A (n_2965), .B (n_2962));
XOR2_X1 i_2070 (.Z (p_0[41]), .A (n_2977), .B (n_2966));
AOI21_X1 i_2069 (.ZN (n_2959), .A (n_3116), .B1 (n_1353), .B2 (n_1396));
OAI21_X1 i_2068 (.ZN (n_2958), .A (n_3074), .B1 (n_1209), .B2 (n_1258));
AOI21_X1 i_2067 (.ZN (n_2957), .A (n_3117), .B1 (n_3074), .B2 (n_2979));
OAI21_X1 i_2066 (.ZN (n_2956), .A (n_3113), .B1 (n_3072), .B2 (n_2957));
INV_X1 i_2065 (.ZN (n_2955), .A (n_2956));
NOR2_X1 i_2064 (.ZN (n_2954), .A1 (n_3114), .A2 (n_3072));
OAI21_X1 i_2063 (.ZN (n_2953), .A (n_3111), .B1 (n_3070), .B2 (n_2955));
XNOR2_X1 i_2062 (.ZN (p_0[40]), .A (n_2959), .B (n_2953));
NOR2_X1 i_2061 (.ZN (n_2952), .A1 (n_3112), .A2 (n_3070));
XOR2_X1 i_2060 (.Z (p_0[39]), .A (n_2955), .B (n_2952));
XOR2_X1 i_2059 (.Z (p_0[38]), .A (n_2957), .B (n_2954));
XOR2_X1 i_2058 (.Z (p_0[37]), .A (n_2979), .B (n_2958));
AOI21_X1 i_2057 (.ZN (n_2951), .A (n_3091), .B1 (n_1157), .B2 (n_1208));
OAI21_X1 i_2056 (.ZN (n_2950), .A (n_3081), .B1 (n_989), .B2 (n_1046));
AOI21_X1 i_2055 (.ZN (n_2949), .A (n_3084), .B1 (sgo__n208), .B2 (n_3081));
OAI21_X1 i_2054 (.ZN (n_2948), .A (n_3088), .B1 (n_3079), .B2 (n_2949));
INV_X1 i_2053 (.ZN (n_2947), .A (n_2948));
NOR2_X1 i_2052 (.ZN (n_2946), .A1 (n_3089), .A2 (n_3079));
OAI21_X1 i_2051 (.ZN (n_2945), .A (n_3086), .B1 (n_3077), .B2 (n_2947));
XNOR2_X2 i_2050 (.ZN (p_0[36]), .A (n_2951), .B (n_2945));
NOR2_X1 i_2049 (.ZN (n_2944), .A1 (n_3087), .A2 (n_3077));
XOR2_X2 i_2048 (.Z (p_0[35]), .A (n_2947), .B (n_2944));
XOR2_X1 i_2047 (.Z (p_0[34]), .A (n_2949), .B (n_2946));
XOR2_X1 i_2046 (.Z (p_0[33]), .A (sgo__n208), .B (n_2950));
OAI21_X1 i_2045 (.ZN (n_2943), .A (n_3172), .B1 (n_3245), .B2 (n_3244));
OAI21_X1 i_2044 (.ZN (n_2942), .A (n_3138), .B1 (n_3183), .B2 (n_3145));
INV_X1 i_2043 (.ZN (n_2941), .A (n_2942));
OAI21_X1 i_2042 (.ZN (n_2940), .A (n_3120), .B1 (n_3174), .B2 (n_2941));
INV_X1 i_2041 (.ZN (n_2939), .A (n_2940));
OAI21_X1 i_2040 (.ZN (n_2938), .A (n_3132), .B1 (n_3156), .B2 (n_2939));
INV_X1 i_2039 (.ZN (n_2937), .A (n_2938));
OAI21_X1 i_2038 (.ZN (n_2936), .A (n_3131), .B1 (n_755), .B2 (n_810));
AOI21_X1 i_2037 (.ZN (n_2935), .A (n_3166), .B1 (n_3131), .B2 (n_2937));
OAI21_X1 i_2036 (.ZN (n_2934), .A (n_3170), .B1 (n_3130), .B2 (n_2935));
INV_X1 i_2035 (.ZN (n_2933), .A (n_2934));
NOR2_X1 i_2034 (.ZN (n_2932), .A1 (n_3171), .A2 (n_3130));
OAI21_X1 i_2033 (.ZN (n_2931), .A (n_3168), .B1 (n_3127), .B2 (n_2933));
XOR2_X1 i_2032 (.Z (p_0[32]), .A (n_2943), .B (n_2931));
NOR2_X1 i_2031 (.ZN (n_2930), .A1 (n_3169), .A2 (n_3127));
XOR2_X1 i_2030 (.Z (p_0[31]), .A (n_2933), .B (n_2930));
XOR2_X1 i_2029 (.Z (p_0[30]), .A (n_2935), .B (n_2932));
XOR2_X1 i_2028 (.Z (p_0[29]), .A (n_2937), .B (n_2936));
AOI21_X1 i_2027 (.ZN (n_2929), .A (n_3164), .B1 (n_701), .B2 (n_754));
OAI21_X1 i_2026 (.ZN (n_2928), .A (n_3137), .B1 (n_596), .B2 (n_598));
AOI21_X1 i_2025 (.ZN (n_2927), .A (n_3157), .B1 (n_3137), .B2 (n_2939));
OAI21_X1 i_2024 (.ZN (n_2926), .A (n_3161), .B1 (n_3135), .B2 (n_2927));
INV_X1 i_2023 (.ZN (n_2925), .A (n_2926));
NOR2_X1 i_2022 (.ZN (n_2924), .A1 (n_3162), .A2 (n_3135));
OAI21_X1 i_2021 (.ZN (n_2923), .A (n_3159), .B1 (n_3133), .B2 (n_2925));
XNOR2_X1 i_2020 (.ZN (p_0[28]), .A (n_2929), .B (n_2923));
NOR2_X1 i_2019 (.ZN (n_2922), .A1 (n_3160), .A2 (n_3133));
XOR2_X1 i_2018 (.Z (p_0[27]), .A (n_2925), .B (n_2922));
XOR2_X1 i_2017 (.Z (p_0[26]), .A (n_2927), .B (n_2924));
XOR2_X1 i_2016 (.Z (p_0[25]), .A (n_2939), .B (n_2928));
AOI21_X1 i_2015 (.ZN (n_2921), .A (n_3181), .B1 (n_505), .B2 (n_550));
OAI21_X1 i_2014 (.ZN (n_2920), .A (n_3125), .B1 (n_379), .B2 (n_418));
AOI21_X1 i_2013 (.ZN (n_2919), .A (n_3182), .B1 (n_3125), .B2 (n_2941));
OAI21_X1 i_2012 (.ZN (n_2918), .A (n_3178), .B1 (n_3123), .B2 (n_2919));
INV_X1 i_2011 (.ZN (n_2917), .A (n_2918));
NOR2_X1 i_2010 (.ZN (n_2916), .A1 (n_3179), .A2 (n_3123));
OAI21_X1 i_2009 (.ZN (n_2915), .A (n_3176), .B1 (n_3121), .B2 (n_2917));
XNOR2_X1 i_2008 (.ZN (p_0[24]), .A (n_2921), .B (n_2915));
NOR2_X1 i_2007 (.ZN (n_2914), .A1 (n_3177), .A2 (n_3121));
XOR2_X1 i_2006 (.Z (p_0[23]), .A (n_2917), .B (n_2914));
XOR2_X1 i_2005 (.Z (p_0[22]), .A (n_2919), .B (n_2916));
XOR2_X1 i_2004 (.Z (p_0[21]), .A (n_2941), .B (n_2920));
AOI21_X1 i_2003 (.ZN (n_2913), .A (n_3153), .B1 (n_376), .B2 (n_378));
OAI21_X1 i_2002 (.ZN (n_2912), .A (n_3143), .B1 (n_268), .B2 (n_270));
AOI21_X1 i_2001 (.ZN (n_2911), .A (n_3146), .B1 (n_3183), .B2 (n_3143));
OAI21_X1 i_2000 (.ZN (n_2910), .A (n_3150), .B1 (n_3141), .B2 (n_2911));
INV_X1 i_1999 (.ZN (n_2909), .A (n_2910));
NOR2_X1 i_1998 (.ZN (n_2908), .A1 (n_3151), .A2 (n_3141));
OAI21_X1 i_1997 (.ZN (n_2907), .A (n_3148), .B1 (n_3139), .B2 (n_2909));
XNOR2_X1 i_1996 (.ZN (p_0[20]), .A (n_2913), .B (n_2907));
NOR2_X1 i_1995 (.ZN (n_2906), .A1 (n_3149), .A2 (n_3139));
XOR2_X1 i_1994 (.Z (p_0[19]), .A (n_2909), .B (n_2906));
XOR2_X1 i_1993 (.Z (p_0[18]), .A (n_2911), .B (n_2908));
XOR2_X1 i_1992 (.Z (p_0[17]), .A (n_3183), .B (n_2912));
NOR2_X1 i_1991 (.ZN (n_2905), .A1 (n_3196), .A2 (n_3187));
OAI21_X1 i_1990 (.ZN (n_2904), .A (n_3190), .B1 (n_152), .B2 (n_154));
AOI21_X1 i_1989 (.ZN (n_2903), .A (n_3192), .B1 (n_3197), .B2 (n_3190));
INV_X1 i_1988 (.ZN (n_2902), .A (n_2903));
AOI21_X1 i_1987 (.ZN (n_2901), .A (n_3195), .B1 (n_3189), .B2 (n_2902));
AOI21_X1 i_1986 (.ZN (n_2900), .A (n_3195), .B1 (n_178), .B2 (n_180));
OAI22_X1 i_1985 (.ZN (n_2899), .A1 (n_206), .A2 (n_208), .B1 (n_3185), .B2 (n_2901));
XNOR2_X1 i_1984 (.ZN (p_0[16]), .A (n_2905), .B (n_2899));
NOR2_X1 i_1983 (.ZN (n_2898), .A1 (n_3194), .A2 (n_3185));
XOR2_X1 i_1982 (.Z (p_0[15]), .A (n_2901), .B (n_2898));
XOR2_X1 i_1981 (.Z (p_0[14]), .A (n_2903), .B (n_2900));
XOR2_X1 i_1980 (.Z (p_0[13]), .A (n_3197), .B (n_2904));
NOR2_X1 i_1979 (.ZN (n_2897), .A1 (n_3210), .A2 (n_3201));
OAI21_X1 i_1978 (.ZN (n_2896), .A (n_3204), .B1 (n_68), .B2 (n_70));
AOI21_X1 i_1977 (.ZN (n_2895), .A (n_3206), .B1 (n_3211), .B2 (n_3204));
INV_X1 i_1976 (.ZN (n_2894), .A (n_2895));
AOI21_X1 i_1975 (.ZN (n_2893), .A (n_3209), .B1 (n_3203), .B2 (n_2894));
AOI21_X1 i_1974 (.ZN (n_2892), .A (n_3209), .B1 (n_86), .B2 (n_88));
OAI22_X1 i_1973 (.ZN (n_2891), .A1 (n_106), .A2 (n_108), .B1 (n_3199), .B2 (n_2893));
XNOR2_X1 i_1972 (.ZN (p_0[12]), .A (n_2897), .B (n_2891));
NOR2_X1 i_1971 (.ZN (n_2890), .A1 (n_3208), .A2 (n_3199));
XOR2_X1 i_1970 (.Z (p_0[11]), .A (n_2893), .B (n_2890));
XOR2_X1 i_1969 (.Z (p_0[10]), .A (n_2895), .B (n_2892));
XOR2_X1 i_1968 (.Z (p_0[9]), .A (n_3211), .B (n_2896));
NOR2_X1 i_1967 (.ZN (n_2889), .A1 (n_3224), .A2 (n_3215));
OAI21_X1 i_1966 (.ZN (n_2888), .A (n_3218), .B1 (n_16), .B2 (n_18));
AOI21_X1 i_1965 (.ZN (n_2887), .A (n_3220), .B1 (n_3225), .B2 (n_3218));
INV_X1 i_1964 (.ZN (n_2886), .A (n_2887));
AOI21_X1 i_1963 (.ZN (n_2885), .A (n_3223), .B1 (n_3217), .B2 (n_2886));
AOI21_X1 i_1962 (.ZN (n_2884), .A (n_3223), .B1 (n_26), .B2 (n_28));
OAI22_X1 i_1961 (.ZN (n_2883), .A1 (n_38), .A2 (n_40), .B1 (n_3213), .B2 (n_2885));
XNOR2_X1 i_1960 (.ZN (p_0[8]), .A (n_2889), .B (n_2883));
NOR2_X1 i_1959 (.ZN (n_2882), .A1 (n_3222), .A2 (n_3213));
XOR2_X1 i_1958 (.Z (p_0[7]), .A (n_2885), .B (n_2882));
XOR2_X1 i_1957 (.Z (p_0[6]), .A (n_2887), .B (n_2884));
XOR2_X1 i_1956 (.Z (p_0[5]), .A (n_3225), .B (n_2888));
XOR2_X1 i_1955 (.Z (n_2881), .A (n_6), .B (n_10));
XOR2_X1 i_1954 (.Z (p_0[4]), .A (n_3226), .B (n_2881));
OAI21_X1 i_1953 (.ZN (n_2880), .A (n_3236), .B1 (n_2), .B2 (n_4));
XNOR2_X1 i_1952 (.ZN (p_0[3]), .A (n_3228), .B (n_2880));
OAI21_X1 i_1951 (.ZN (n_2879), .A (n_3229), .B1 (n_0), .B2 (n_3235));
XOR2_X1 i_1950 (.Z (p_0[2]), .A (n_3230), .B (n_2879));
OAI21_X1 i_1949 (.ZN (n_2878), .A (n_3230), .B1 (n_3233), .B2 (n_3232));
INV_X1 i_1948 (.ZN (p_0[1]), .A (n_2878));
NOR2_X1 i_1947 (.ZN (n_2877), .A1 (n_3278), .A2 (sgo__n10));
NOR2_X1 i_1946 (.ZN (n_2876), .A1 (n_3278), .A2 (n_3250));
NOR2_X1 i_1945 (.ZN (n_2875), .A1 (n_3278), .A2 (n_3251));
NOR2_X1 i_1944 (.ZN (n_2874), .A1 (n_3278), .A2 (n_3252));
NOR2_X1 i_1943 (.ZN (n_2873), .A1 (n_3278), .A2 (n_3253));
NOR2_X1 i_1942 (.ZN (n_2872), .A1 (n_3278), .A2 (n_3254));
NOR2_X1 i_1941 (.ZN (n_2871), .A1 (n_3278), .A2 (n_3255));
NOR2_X1 i_1940 (.ZN (n_2870), .A1 (n_3278), .A2 (sgo__n182));
NOR2_X1 i_1939 (.ZN (n_2869), .A1 (n_3278), .A2 (n_3257));
NOR2_X1 i_1938 (.ZN (n_2868), .A1 (n_3278), .A2 (n_3258));
NOR2_X1 i_1937 (.ZN (n_2867), .A1 (n_3278), .A2 (n_3259));
NOR2_X1 i_1936 (.ZN (n_2866), .A1 (n_3278), .A2 (n_3260));
NOR2_X1 i_1935 (.ZN (n_2865), .A1 (n_3278), .A2 (sgo__n148));
NOR2_X1 i_1934 (.ZN (n_2864), .A1 (n_3278), .A2 (n_3262));
NOR2_X1 i_1933 (.ZN (n_2863), .A1 (n_3278), .A2 (n_3263));
NOR2_X1 i_1932 (.ZN (n_2862), .A1 (n_3278), .A2 (n_3264));
NOR2_X1 i_1931 (.ZN (n_2861), .A1 (n_3278), .A2 (n_3265));
NOR2_X1 i_1930 (.ZN (n_2860), .A1 (n_3278), .A2 (n_3266));
NOR2_X1 i_1929 (.ZN (n_2859), .A1 (n_3278), .A2 (n_3267));
NOR2_X1 i_1928 (.ZN (n_2858), .A1 (n_3278), .A2 (n_3268));
NOR2_X1 i_1927 (.ZN (n_2857), .A1 (n_3278), .A2 (n_3269));
NOR2_X1 i_1926 (.ZN (n_2856), .A1 (n_3278), .A2 (n_3270));
NOR2_X1 i_1925 (.ZN (n_2855), .A1 (n_3278), .A2 (n_3271));
NOR2_X1 i_1924 (.ZN (n_2854), .A1 (n_3278), .A2 (n_3272));
NOR2_X1 i_1923 (.ZN (n_2853), .A1 (n_3278), .A2 (n_3273));
NOR2_X1 i_1922 (.ZN (n_2852), .A1 (n_3278), .A2 (n_3274));
NOR2_X1 i_1921 (.ZN (n_2851), .A1 (n_3278), .A2 (n_3275));
NOR2_X1 i_1920 (.ZN (n_2850), .A1 (n_3278), .A2 (n_3276));
NOR2_X1 i_1919 (.ZN (n_2849), .A1 (n_3278), .A2 (n_3277));
NOR2_X1 i_1918 (.ZN (n_2848), .A1 (n_3279), .A2 (n_3248));
NOR2_X1 i_1917 (.ZN (n_2847), .A1 (n_3279), .A2 (sgo__n10));
NOR2_X1 i_1916 (.ZN (n_2846), .A1 (n_3279), .A2 (n_3250));
NOR2_X2 i_1915 (.ZN (n_2845), .A1 (n_3279), .A2 (n_3251));
NOR2_X1 i_1914 (.ZN (n_2844), .A1 (n_3279), .A2 (n_3252));
NOR2_X1 i_1913 (.ZN (n_2843), .A1 (n_3279), .A2 (n_3253));
NOR2_X1 i_1912 (.ZN (n_2842), .A1 (n_3279), .A2 (n_3254));
NOR2_X1 i_1911 (.ZN (n_2841), .A1 (n_3279), .A2 (n_3255));
NOR2_X1 i_1910 (.ZN (n_2840), .A1 (n_3279), .A2 (sgo__n182));
NOR2_X1 i_1909 (.ZN (n_2839), .A1 (n_3279), .A2 (n_3257));
NOR2_X1 i_1908 (.ZN (n_2838), .A1 (n_3279), .A2 (n_3258));
NOR2_X1 i_1907 (.ZN (n_2837), .A1 (n_3279), .A2 (n_3259));
NOR2_X1 i_1906 (.ZN (n_2836), .A1 (n_3279), .A2 (n_3260));
NOR2_X1 i_1905 (.ZN (n_2835), .A1 (n_3279), .A2 (sgo__n148));
NOR2_X1 i_1904 (.ZN (n_2834), .A1 (n_3279), .A2 (n_3262));
NOR2_X4 i_1903 (.ZN (n_2833), .A1 (n_3279), .A2 (n_3263));
NOR2_X1 i_1902 (.ZN (n_2832), .A1 (n_3279), .A2 (n_3264));
NOR2_X1 i_1901 (.ZN (n_2831), .A1 (n_3279), .A2 (n_3265));
NOR2_X1 i_1900 (.ZN (n_2830), .A1 (n_3279), .A2 (n_3266));
NOR2_X1 i_1899 (.ZN (n_2829), .A1 (n_3279), .A2 (n_3267));
NOR2_X1 i_1898 (.ZN (n_2828), .A1 (n_3279), .A2 (n_3268));
NOR2_X1 i_1897 (.ZN (n_2827), .A1 (n_3279), .A2 (n_3269));
NOR2_X1 i_1896 (.ZN (n_2826), .A1 (n_3279), .A2 (n_3270));
NOR2_X1 i_1895 (.ZN (n_2825), .A1 (n_3279), .A2 (n_3271));
NOR2_X1 i_1894 (.ZN (n_2824), .A1 (n_3279), .A2 (n_3272));
NOR2_X1 i_1893 (.ZN (n_2823), .A1 (n_3279), .A2 (n_3273));
NOR2_X1 i_1892 (.ZN (n_2822), .A1 (n_3279), .A2 (n_3274));
NOR2_X1 i_1891 (.ZN (n_2821), .A1 (n_3279), .A2 (n_3275));
NOR2_X1 i_1890 (.ZN (n_2820), .A1 (n_3279), .A2 (n_3276));
NOR2_X1 i_1889 (.ZN (n_2819), .A1 (n_3279), .A2 (n_3277));
NOR2_X1 i_1888 (.ZN (n_2818), .A1 (n_3280), .A2 (n_3246));
NOR2_X1 i_1887 (.ZN (n_2817), .A1 (n_3280), .A2 (n_3247));
NOR2_X1 i_1886 (.ZN (n_2816), .A1 (n_3280), .A2 (n_3248));
NOR2_X1 i_1885 (.ZN (n_2815), .A1 (n_3280), .A2 (sgo__n10));
NOR2_X1 i_1884 (.ZN (n_2814), .A1 (n_3280), .A2 (n_3250));
NOR2_X1 i_1883 (.ZN (n_2813), .A1 (n_3280), .A2 (n_3251));
NOR2_X1 i_1882 (.ZN (n_2812), .A1 (n_3280), .A2 (n_3252));
NOR2_X1 i_1881 (.ZN (n_2811), .A1 (n_3280), .A2 (n_3253));
NOR2_X1 i_1880 (.ZN (n_2810), .A1 (n_3280), .A2 (n_3254));
NOR2_X1 i_1879 (.ZN (n_2809), .A1 (n_3280), .A2 (n_3255));
NOR2_X1 i_1878 (.ZN (n_2808), .A1 (n_3280), .A2 (sgo__n182));
NOR2_X1 i_1877 (.ZN (n_2807), .A1 (n_3280), .A2 (n_3257));
NOR2_X1 i_1876 (.ZN (n_2806), .A1 (n_3280), .A2 (n_3258));
NOR2_X1 i_1875 (.ZN (n_2805), .A1 (n_3280), .A2 (n_3259));
NOR2_X1 i_1874 (.ZN (n_2804), .A1 (n_3280), .A2 (n_3260));
NOR2_X1 i_1873 (.ZN (n_2803), .A1 (n_3280), .A2 (sgo__n148));
NOR2_X4 i_1872 (.ZN (n_2802), .A1 (n_3280), .A2 (n_3262));
NOR2_X1 i_1871 (.ZN (n_2801), .A1 (n_3280), .A2 (n_3263));
NOR2_X1 i_1870 (.ZN (n_2800), .A1 (n_3280), .A2 (n_3264));
NOR2_X1 i_1869 (.ZN (n_2799), .A1 (n_3280), .A2 (n_3265));
NOR2_X1 i_1868 (.ZN (n_2798), .A1 (n_3280), .A2 (n_3266));
NOR2_X1 i_1867 (.ZN (n_2797), .A1 (n_3280), .A2 (n_3267));
NOR2_X1 i_1866 (.ZN (n_2796), .A1 (n_3280), .A2 (n_3268));
NOR2_X1 i_1865 (.ZN (n_2795), .A1 (n_3280), .A2 (n_3269));
NOR2_X1 i_1864 (.ZN (n_2794), .A1 (n_3280), .A2 (sgo__n203));
NOR2_X1 i_1863 (.ZN (n_2793), .A1 (n_3280), .A2 (n_3271));
NOR2_X1 i_1862 (.ZN (n_2792), .A1 (n_3280), .A2 (n_3272));
NOR2_X1 i_1861 (.ZN (n_2791), .A1 (n_3280), .A2 (n_3273));
NOR2_X1 i_1860 (.ZN (n_2790), .A1 (n_3280), .A2 (n_3274));
NOR2_X1 i_1859 (.ZN (n_2789), .A1 (n_3280), .A2 (n_3275));
NOR2_X1 i_1858 (.ZN (n_2788), .A1 (n_3280), .A2 (n_3276));
NOR2_X1 i_1857 (.ZN (n_2787), .A1 (n_3280), .A2 (n_3277));
NOR2_X1 i_1856 (.ZN (n_2786), .A1 (n_3281), .A2 (n_3246));
NOR2_X1 i_1855 (.ZN (n_2785), .A1 (n_3281), .A2 (n_3247));
NOR2_X1 i_1854 (.ZN (n_2784), .A1 (n_3281), .A2 (n_3248));
NOR2_X1 i_1853 (.ZN (n_2783), .A1 (n_3281), .A2 (sgo__n10));
NOR2_X1 i_1852 (.ZN (n_2782), .A1 (n_3281), .A2 (n_3250));
NOR2_X1 i_1851 (.ZN (n_2781), .A1 (n_3281), .A2 (n_3251));
NOR2_X1 i_1850 (.ZN (n_2780), .A1 (n_3281), .A2 (n_3252));
NOR2_X1 i_1849 (.ZN (n_2779), .A1 (n_3281), .A2 (n_3253));
NOR2_X1 i_1848 (.ZN (n_2778), .A1 (n_3281), .A2 (n_3254));
NOR2_X1 i_1847 (.ZN (n_2777), .A1 (n_3281), .A2 (n_3255));
NOR2_X1 i_1846 (.ZN (n_2776), .A1 (n_3281), .A2 (sgo__n182));
NOR2_X1 i_1845 (.ZN (n_2775), .A1 (n_3281), .A2 (n_3257));
NOR2_X1 i_1844 (.ZN (n_2774), .A1 (n_3281), .A2 (n_3258));
NOR2_X1 i_1843 (.ZN (n_2773), .A1 (n_3281), .A2 (n_3259));
NOR2_X1 i_1842 (.ZN (n_2772), .A1 (n_3281), .A2 (n_3260));
NOR2_X1 i_1841 (.ZN (n_2771), .A1 (n_3281), .A2 (sgo__n148));
NOR2_X1 i_1840 (.ZN (n_2770), .A1 (n_3281), .A2 (n_3262));
NOR2_X1 i_1839 (.ZN (n_2769), .A1 (n_3281), .A2 (n_3263));
NOR2_X1 i_1838 (.ZN (n_2768), .A1 (n_3281), .A2 (n_3264));
NOR2_X1 i_1837 (.ZN (n_2767), .A1 (n_3281), .A2 (n_3265));
NOR2_X1 i_1836 (.ZN (n_2766), .A1 (n_3281), .A2 (n_3266));
NOR2_X1 i_1835 (.ZN (n_2765), .A1 (n_3281), .A2 (n_3267));
NOR2_X1 i_1834 (.ZN (n_2764), .A1 (n_3281), .A2 (n_3268));
NOR2_X1 i_1833 (.ZN (n_2763), .A1 (n_3281), .A2 (n_3269));
NOR2_X1 i_1832 (.ZN (n_2762), .A1 (n_3281), .A2 (n_3270));
NOR2_X1 i_1831 (.ZN (n_2761), .A1 (n_3281), .A2 (n_3271));
NOR2_X1 i_1830 (.ZN (n_2760), .A1 (n_3281), .A2 (n_3272));
NOR2_X1 i_1829 (.ZN (n_2759), .A1 (n_3281), .A2 (n_3273));
NOR2_X1 i_1828 (.ZN (n_2758), .A1 (n_3281), .A2 (n_3274));
NOR2_X1 i_1827 (.ZN (n_2757), .A1 (n_3281), .A2 (n_3275));
NOR2_X1 i_1826 (.ZN (n_2756), .A1 (n_3281), .A2 (n_3276));
NOR2_X1 i_1825 (.ZN (n_2755), .A1 (n_3281), .A2 (n_3277));
NOR2_X1 i_1824 (.ZN (n_2754), .A1 (n_3282), .A2 (n_3246));
NOR2_X1 i_1823 (.ZN (n_2753), .A1 (n_3282), .A2 (n_3247));
NOR2_X1 i_1822 (.ZN (n_2752), .A1 (n_3282), .A2 (n_3248));
NOR2_X1 i_1821 (.ZN (n_2751), .A1 (n_3282), .A2 (sgo__n10));
NOR2_X1 i_1820 (.ZN (n_2750), .A1 (n_3282), .A2 (n_3250));
NOR2_X1 i_1819 (.ZN (n_2749), .A1 (n_3282), .A2 (n_3251));
NOR2_X1 i_1818 (.ZN (n_2748), .A1 (n_3282), .A2 (n_3252));
NOR2_X1 i_1817 (.ZN (n_2747), .A1 (n_3282), .A2 (n_3253));
NOR2_X1 i_1816 (.ZN (n_2746), .A1 (n_3282), .A2 (n_3254));
NOR2_X1 i_1815 (.ZN (n_2745), .A1 (n_3282), .A2 (n_3255));
NOR2_X1 i_1814 (.ZN (n_2744), .A1 (n_3282), .A2 (sgo__n182));
NOR2_X1 i_1813 (.ZN (n_2743), .A1 (n_3282), .A2 (n_3257));
NOR2_X1 i_1812 (.ZN (n_2742), .A1 (n_3282), .A2 (n_3258));
NOR2_X1 i_1811 (.ZN (n_2741), .A1 (n_3282), .A2 (n_3259));
NOR2_X1 i_1810 (.ZN (n_2740), .A1 (n_3282), .A2 (n_3260));
NOR2_X1 i_1809 (.ZN (n_2739), .A1 (n_3282), .A2 (n_3261));
NOR2_X1 i_1808 (.ZN (n_2738), .A1 (n_3282), .A2 (n_3262));
NOR2_X1 i_1807 (.ZN (n_2737), .A1 (n_3282), .A2 (n_3263));
NOR2_X1 i_1806 (.ZN (n_2736), .A1 (n_3282), .A2 (n_3264));
NOR2_X1 i_1805 (.ZN (n_2735), .A1 (n_3282), .A2 (n_3265));
NOR2_X1 i_1804 (.ZN (n_2734), .A1 (n_3282), .A2 (n_3266));
NOR2_X1 i_1803 (.ZN (n_2733), .A1 (n_3282), .A2 (n_3267));
NOR2_X1 i_1802 (.ZN (n_2732), .A1 (n_3282), .A2 (sgo__n170));
NOR2_X1 i_1801 (.ZN (n_2731), .A1 (n_3282), .A2 (n_3269));
NOR2_X1 i_1800 (.ZN (n_2730), .A1 (n_3282), .A2 (n_3270));
NOR2_X1 i_1799 (.ZN (n_2729), .A1 (n_3282), .A2 (n_3271));
NOR2_X1 i_1798 (.ZN (n_2728), .A1 (n_3282), .A2 (n_3272));
NOR2_X1 i_1797 (.ZN (n_2727), .A1 (n_3282), .A2 (n_3273));
NOR2_X1 i_1796 (.ZN (n_2726), .A1 (n_3282), .A2 (n_3274));
NOR2_X1 i_1795 (.ZN (n_2725), .A1 (n_3282), .A2 (n_3275));
NOR2_X1 i_1794 (.ZN (n_2724), .A1 (n_3282), .A2 (n_3276));
NOR2_X1 i_1793 (.ZN (n_2723), .A1 (n_3282), .A2 (n_3277));
NOR2_X1 i_1792 (.ZN (n_2722), .A1 (n_3283), .A2 (n_3246));
NOR2_X1 i_1791 (.ZN (n_2721), .A1 (n_3283), .A2 (n_3247));
NOR2_X1 i_1790 (.ZN (n_2720), .A1 (n_3283), .A2 (n_3248));
NOR2_X1 i_1789 (.ZN (n_2719), .A1 (n_3283), .A2 (sgo__n10));
NOR2_X1 i_1788 (.ZN (n_2718), .A1 (n_3283), .A2 (n_3250));
NOR2_X1 i_1787 (.ZN (n_2717), .A1 (n_3283), .A2 (n_3251));
NOR2_X1 i_1786 (.ZN (n_2716), .A1 (n_3283), .A2 (n_3252));
NOR2_X1 i_1785 (.ZN (n_2715), .A1 (n_3283), .A2 (n_3253));
NOR2_X1 i_1784 (.ZN (n_2714), .A1 (n_3283), .A2 (n_3254));
NOR2_X1 i_1783 (.ZN (n_2713), .A1 (n_3283), .A2 (n_3255));
NOR2_X1 i_1782 (.ZN (n_2712), .A1 (n_3283), .A2 (n_3256));
NOR2_X1 i_1781 (.ZN (n_2711), .A1 (n_3283), .A2 (n_3257));
NOR2_X1 i_1780 (.ZN (n_2710), .A1 (n_3283), .A2 (n_3258));
NOR2_X1 i_1779 (.ZN (n_2709), .A1 (n_3283), .A2 (n_3259));
NOR2_X1 i_1778 (.ZN (n_2708), .A1 (n_3283), .A2 (n_3260));
NOR2_X1 i_1777 (.ZN (n_2707), .A1 (n_3283), .A2 (n_3261));
NOR2_X1 i_1776 (.ZN (n_2706), .A1 (n_3283), .A2 (n_3262));
NOR2_X1 i_1775 (.ZN (n_2705), .A1 (n_3283), .A2 (n_3263));
NOR2_X1 i_1774 (.ZN (n_2704), .A1 (n_3283), .A2 (n_3264));
NOR2_X1 i_1773 (.ZN (n_2703), .A1 (n_3283), .A2 (n_3265));
NOR2_X1 i_1772 (.ZN (n_2702), .A1 (n_3283), .A2 (n_3266));
NOR2_X1 i_1771 (.ZN (n_2701), .A1 (n_3283), .A2 (n_3267));
NOR2_X1 i_1770 (.ZN (n_2700), .A1 (n_3283), .A2 (n_3268));
NOR2_X1 i_1769 (.ZN (n_2699), .A1 (n_3283), .A2 (n_3269));
NOR2_X1 i_1768 (.ZN (n_2698), .A1 (n_3283), .A2 (n_3270));
NOR2_X1 i_1767 (.ZN (n_2697), .A1 (n_3283), .A2 (n_3271));
NOR2_X4 i_1766 (.ZN (n_2696), .A1 (n_3283), .A2 (n_3272));
NOR2_X1 i_1765 (.ZN (n_2695), .A1 (n_3283), .A2 (n_3273));
NOR2_X1 i_1764 (.ZN (n_2694), .A1 (n_3283), .A2 (n_3274));
NOR2_X1 i_1763 (.ZN (n_2693), .A1 (n_3283), .A2 (n_3275));
NOR2_X1 i_1762 (.ZN (n_2692), .A1 (n_3283), .A2 (n_3276));
NOR2_X1 i_1761 (.ZN (n_2691), .A1 (n_3283), .A2 (n_3277));
NOR2_X1 i_1760 (.ZN (n_2690), .A1 (n_3284), .A2 (n_3246));
NOR2_X1 i_1759 (.ZN (n_2689), .A1 (n_3284), .A2 (n_3247));
NOR2_X1 i_1758 (.ZN (n_2688), .A1 (n_3284), .A2 (n_3248));
NOR2_X1 i_1757 (.ZN (n_2687), .A1 (n_3284), .A2 (sgo__n10));
NOR2_X1 i_1756 (.ZN (n_2686), .A1 (n_3284), .A2 (n_3250));
NOR2_X1 i_1755 (.ZN (n_2685), .A1 (n_3284), .A2 (n_3251));
NOR2_X1 i_1754 (.ZN (n_2684), .A1 (n_3284), .A2 (n_3252));
NOR2_X1 i_1753 (.ZN (n_2683), .A1 (n_3284), .A2 (n_3253));
NOR2_X1 i_1752 (.ZN (n_2682), .A1 (n_3284), .A2 (n_3254));
NOR2_X1 i_1751 (.ZN (n_2681), .A1 (n_3284), .A2 (sgo__n177));
NOR2_X1 i_1750 (.ZN (n_2680), .A1 (n_3284), .A2 (n_3256));
NOR2_X1 i_1749 (.ZN (n_2679), .A1 (n_3284), .A2 (n_3257));
NOR2_X1 i_1748 (.ZN (n_2678), .A1 (n_3284), .A2 (n_3258));
NOR2_X1 i_1747 (.ZN (n_2677), .A1 (n_3284), .A2 (n_3259));
NOR2_X1 i_1746 (.ZN (n_2676), .A1 (n_3284), .A2 (n_3260));
NOR2_X1 i_1745 (.ZN (n_2675), .A1 (n_3284), .A2 (n_3261));
NOR2_X1 i_1744 (.ZN (n_2674), .A1 (n_3284), .A2 (n_3262));
NOR2_X1 i_1743 (.ZN (n_2673), .A1 (n_3284), .A2 (n_3263));
NOR2_X1 i_1742 (.ZN (n_2672), .A1 (n_3284), .A2 (n_3264));
NOR2_X1 i_1741 (.ZN (n_2671), .A1 (n_3284), .A2 (n_3265));
NOR2_X1 i_1740 (.ZN (n_2670), .A1 (n_3284), .A2 (n_3266));
NOR2_X1 i_1739 (.ZN (n_2669), .A1 (n_3284), .A2 (n_3267));
NOR2_X1 i_1738 (.ZN (n_2668), .A1 (n_3284), .A2 (n_3268));
NOR2_X4 i_1737 (.ZN (n_2667), .A1 (n_3284), .A2 (n_3269));
NOR2_X1 i_1736 (.ZN (n_2666), .A1 (n_3284), .A2 (sgo__n203));
NOR2_X1 i_1735 (.ZN (n_2665), .A1 (n_3284), .A2 (n_3271));
NOR2_X1 i_1734 (.ZN (n_2664), .A1 (n_3284), .A2 (n_3272));
NOR2_X1 i_1733 (.ZN (n_2663), .A1 (n_3284), .A2 (n_3273));
NOR2_X1 i_1732 (.ZN (n_2662), .A1 (n_3284), .A2 (n_3274));
NOR2_X1 i_1731 (.ZN (n_2661), .A1 (n_3284), .A2 (n_3275));
NOR2_X1 i_1730 (.ZN (n_2660), .A1 (n_3284), .A2 (n_3276));
NOR2_X1 i_1729 (.ZN (n_2659), .A1 (n_3284), .A2 (n_3277));
NOR2_X1 i_1728 (.ZN (n_2658), .A1 (n_3285), .A2 (n_3246));
NOR2_X1 i_1727 (.ZN (n_2657), .A1 (n_3285), .A2 (n_3247));
NOR2_X1 i_1726 (.ZN (n_2656), .A1 (n_3285), .A2 (n_3248));
NOR2_X1 i_1725 (.ZN (n_2655), .A1 (n_3285), .A2 (sgo__n10));
NOR2_X1 i_1724 (.ZN (n_2654), .A1 (n_3285), .A2 (n_3250));
NOR2_X1 i_1723 (.ZN (n_2653), .A1 (n_3285), .A2 (n_3251));
NOR2_X1 i_1722 (.ZN (n_2652), .A1 (n_3285), .A2 (n_3252));
NOR2_X1 i_1721 (.ZN (n_2651), .A1 (n_3285), .A2 (n_3253));
NOR2_X1 i_1720 (.ZN (n_2650), .A1 (n_3285), .A2 (n_3254));
NOR2_X1 i_1719 (.ZN (n_2649), .A1 (n_3285), .A2 (sgo__n177));
NOR2_X1 i_1718 (.ZN (n_2648), .A1 (n_3285), .A2 (n_3256));
NOR2_X1 i_1717 (.ZN (n_2647), .A1 (n_3285), .A2 (sgo__n134));
NOR2_X1 i_1716 (.ZN (n_2646), .A1 (n_3285), .A2 (n_3258));
NOR2_X1 i_1715 (.ZN (n_2645), .A1 (n_3285), .A2 (n_3259));
NOR2_X1 i_1714 (.ZN (n_2644), .A1 (n_3285), .A2 (n_3260));
NOR2_X1 i_1713 (.ZN (n_2643), .A1 (n_3285), .A2 (n_3261));
NOR2_X1 i_1712 (.ZN (n_2642), .A1 (n_3285), .A2 (n_3262));
NOR2_X1 i_1711 (.ZN (n_2641), .A1 (n_3285), .A2 (n_3263));
NOR2_X1 i_1710 (.ZN (n_2640), .A1 (n_3285), .A2 (n_3264));
NOR2_X1 i_1709 (.ZN (n_2639), .A1 (n_3285), .A2 (n_3265));
NOR2_X1 i_1708 (.ZN (n_2638), .A1 (n_3285), .A2 (n_3266));
NOR2_X1 i_1707 (.ZN (n_2637), .A1 (n_3285), .A2 (n_3267));
NOR2_X1 i_1706 (.ZN (n_2636), .A1 (n_3285), .A2 (n_3268));
NOR2_X1 i_1705 (.ZN (n_2635), .A1 (n_3285), .A2 (n_3269));
NOR2_X1 i_1704 (.ZN (n_2634), .A1 (n_3285), .A2 (n_3270));
NOR2_X1 i_1703 (.ZN (n_2633), .A1 (n_3285), .A2 (n_3271));
NOR2_X1 i_1702 (.ZN (n_2632), .A1 (n_3285), .A2 (n_3272));
NOR2_X1 i_1701 (.ZN (n_2631), .A1 (n_3285), .A2 (n_3273));
NOR2_X1 i_1700 (.ZN (n_2630), .A1 (n_3285), .A2 (n_3274));
NOR2_X1 i_1699 (.ZN (n_2629), .A1 (n_3285), .A2 (n_3275));
NOR2_X1 i_1698 (.ZN (n_2628), .A1 (n_3285), .A2 (n_3276));
NOR2_X1 i_1697 (.ZN (n_2627), .A1 (n_3285), .A2 (n_3277));
NOR2_X1 i_1696 (.ZN (n_2626), .A1 (n_3286), .A2 (n_3246));
NOR2_X1 i_1695 (.ZN (n_2625), .A1 (n_3286), .A2 (n_3247));
NOR2_X1 i_1694 (.ZN (n_2624), .A1 (n_3286), .A2 (n_3248));
NOR2_X1 i_1693 (.ZN (n_2623), .A1 (n_3286), .A2 (sgo__n10));
NOR2_X1 i_1692 (.ZN (n_2622), .A1 (n_3286), .A2 (n_3250));
NOR2_X1 i_1691 (.ZN (n_2621), .A1 (n_3286), .A2 (n_3251));
NOR2_X1 i_1690 (.ZN (n_2620), .A1 (n_3286), .A2 (n_3252));
NOR2_X1 i_1689 (.ZN (n_2619), .A1 (n_3286), .A2 (n_3253));
NOR2_X1 i_1688 (.ZN (n_2618), .A1 (n_3286), .A2 (n_3254));
NOR2_X1 i_1687 (.ZN (n_2617), .A1 (n_3286), .A2 (sgo__n177));
NOR2_X1 i_1686 (.ZN (n_2616), .A1 (sgo__n164), .A2 (n_3256));
NOR2_X1 i_1685 (.ZN (n_2615), .A1 (sgo__n164), .A2 (sgo__n134));
NOR2_X1 i_1684 (.ZN (n_2614), .A1 (sgo__n164), .A2 (n_3258));
NOR2_X1 i_1683 (.ZN (n_2613), .A1 (sgo__n164), .A2 (n_3259));
NOR2_X1 i_1682 (.ZN (n_2612), .A1 (sgo__n164), .A2 (n_3260));
NOR2_X1 i_1681 (.ZN (n_2611), .A1 (sgo__n164), .A2 (n_3261));
NOR2_X1 i_1680 (.ZN (n_2610), .A1 (n_3286), .A2 (n_3262));
NOR2_X1 i_1679 (.ZN (n_2609), .A1 (n_3286), .A2 (n_3263));
NOR2_X1 i_1678 (.ZN (n_2608), .A1 (n_3286), .A2 (n_3264));
NOR2_X1 i_1677 (.ZN (n_2607), .A1 (n_3286), .A2 (n_3265));
NOR2_X1 i_1676 (.ZN (n_2606), .A1 (n_3286), .A2 (n_3266));
NOR2_X1 i_1675 (.ZN (n_2605), .A1 (n_3286), .A2 (sgo__n99));
NOR2_X1 i_1674 (.ZN (n_2604), .A1 (n_3286), .A2 (sgo__n170));
NOR2_X1 i_1673 (.ZN (n_2603), .A1 (n_3286), .A2 (sgo__n168));
NOR2_X1 i_1672 (.ZN (n_2602), .A1 (n_3286), .A2 (n_3270));
NOR2_X1 i_1671 (.ZN (n_2601), .A1 (n_3286), .A2 (n_3271));
NOR2_X1 i_1670 (.ZN (n_2600), .A1 (n_3286), .A2 (n_3272));
NOR2_X1 i_1669 (.ZN (n_2599), .A1 (n_3286), .A2 (n_3273));
NOR2_X1 i_1668 (.ZN (n_2598), .A1 (n_3286), .A2 (n_3274));
NOR2_X1 i_1667 (.ZN (n_2597), .A1 (n_3286), .A2 (n_3275));
NOR2_X1 i_1666 (.ZN (n_2596), .A1 (n_3286), .A2 (n_3276));
NOR2_X1 i_1665 (.ZN (n_2595), .A1 (n_3286), .A2 (n_3277));
NOR2_X1 i_1664 (.ZN (n_2594), .A1 (n_3287), .A2 (n_3246));
NOR2_X1 i_1663 (.ZN (n_2593), .A1 (n_3287), .A2 (n_3247));
NOR2_X1 i_1662 (.ZN (n_2592), .A1 (n_3287), .A2 (n_3248));
NOR2_X1 i_1661 (.ZN (n_2591), .A1 (n_3287), .A2 (sgo__n10));
NOR2_X1 i_1660 (.ZN (n_2590), .A1 (n_3287), .A2 (n_3250));
NOR2_X1 i_1659 (.ZN (n_2589), .A1 (n_3287), .A2 (n_3251));
NOR2_X1 i_1658 (.ZN (n_2588), .A1 (n_3287), .A2 (n_3252));
NOR2_X1 i_1657 (.ZN (n_2587), .A1 (n_3287), .A2 (n_3253));
NOR2_X1 i_1656 (.ZN (n_2586), .A1 (n_3287), .A2 (n_3254));
NOR2_X1 i_1655 (.ZN (n_2585), .A1 (n_3287), .A2 (sgo__n178));
NOR2_X1 i_1654 (.ZN (n_2584), .A1 (n_3287), .A2 (n_3256));
NOR2_X1 i_1653 (.ZN (n_2583), .A1 (n_3287), .A2 (sgo__n134));
NOR2_X1 i_1652 (.ZN (n_2582), .A1 (n_3287), .A2 (n_3258));
NOR2_X1 i_1651 (.ZN (n_2581), .A1 (n_3287), .A2 (n_3259));
NOR2_X1 i_1650 (.ZN (n_2580), .A1 (n_3287), .A2 (n_3260));
NOR2_X1 i_1649 (.ZN (n_2579), .A1 (n_3287), .A2 (n_3261));
NOR2_X1 i_1648 (.ZN (n_2578), .A1 (n_3287), .A2 (n_3262));
NOR2_X1 i_1647 (.ZN (n_2577), .A1 (n_3287), .A2 (n_3263));
NOR2_X1 i_1646 (.ZN (n_2576), .A1 (n_3287), .A2 (n_3264));
NOR2_X1 i_1645 (.ZN (n_2575), .A1 (n_3287), .A2 (n_3265));
NOR2_X1 i_1644 (.ZN (n_2574), .A1 (n_3287), .A2 (n_3266));
NOR2_X1 i_1643 (.ZN (n_2573), .A1 (n_3287), .A2 (sgo__n99));
NOR2_X1 i_1642 (.ZN (n_2572), .A1 (n_3287), .A2 (sgo__n172));
NOR2_X1 i_1641 (.ZN (n_2571), .A1 (n_3287), .A2 (sgo__n168));
NOR2_X1 i_1640 (.ZN (n_2570), .A1 (n_3287), .A2 (n_3270));
NOR2_X1 i_1639 (.ZN (n_2569), .A1 (n_3287), .A2 (n_3271));
NOR2_X1 i_1638 (.ZN (n_2568), .A1 (n_3287), .A2 (n_3272));
NOR2_X1 i_1637 (.ZN (n_2567), .A1 (n_3287), .A2 (n_3273));
NOR2_X1 i_1636 (.ZN (n_2566), .A1 (n_3287), .A2 (n_3274));
NOR2_X1 i_1635 (.ZN (n_2565), .A1 (n_3287), .A2 (n_3275));
NOR2_X1 i_1634 (.ZN (n_2564), .A1 (n_3287), .A2 (n_3276));
NOR2_X1 i_1633 (.ZN (n_2563), .A1 (n_3287), .A2 (n_3277));
NOR2_X1 i_1632 (.ZN (n_2562), .A1 (n_3288), .A2 (n_3246));
NOR2_X1 i_1631 (.ZN (n_2561), .A1 (n_3288), .A2 (n_3247));
NOR2_X1 i_1630 (.ZN (n_2560), .A1 (n_3288), .A2 (n_3248));
NOR2_X1 i_1629 (.ZN (n_2559), .A1 (n_3288), .A2 (sgo__n10));
NOR2_X1 i_1628 (.ZN (n_2558), .A1 (n_3288), .A2 (n_3250));
NOR2_X1 i_1627 (.ZN (n_2557), .A1 (n_3288), .A2 (n_3251));
NOR2_X1 i_1626 (.ZN (n_2556), .A1 (n_3288), .A2 (n_3252));
NOR2_X1 i_1625 (.ZN (n_2555), .A1 (n_3288), .A2 (n_3253));
NOR2_X1 i_1624 (.ZN (n_2554), .A1 (n_3288), .A2 (n_3254));
NOR2_X1 i_1623 (.ZN (n_2553), .A1 (n_3288), .A2 (sgo__n178));
NOR2_X1 i_1622 (.ZN (n_2552), .A1 (n_3288), .A2 (n_3256));
NOR2_X1 i_1621 (.ZN (n_2551), .A1 (n_3288), .A2 (sgo__n134));
NOR2_X1 i_1620 (.ZN (n_2550), .A1 (n_3288), .A2 (n_3258));
NOR2_X1 i_1619 (.ZN (n_2549), .A1 (n_3288), .A2 (n_3259));
NOR2_X1 i_1618 (.ZN (n_2548), .A1 (n_3288), .A2 (n_3260));
NOR2_X1 i_1617 (.ZN (n_2547), .A1 (n_3288), .A2 (n_3261));
NOR2_X1 i_1616 (.ZN (n_2546), .A1 (n_3288), .A2 (n_3262));
NOR2_X1 i_1615 (.ZN (n_2545), .A1 (n_3288), .A2 (n_3263));
NOR2_X1 i_1614 (.ZN (n_2544), .A1 (n_3288), .A2 (n_3264));
NOR2_X1 i_1613 (.ZN (n_2543), .A1 (n_3288), .A2 (n_3265));
NOR2_X1 i_1612 (.ZN (n_2542), .A1 (n_3288), .A2 (n_3266));
NOR2_X1 i_1611 (.ZN (n_2541), .A1 (n_3288), .A2 (sgo__n99));
NOR2_X1 i_1610 (.ZN (n_2540), .A1 (n_3288), .A2 (sgo__n172));
NOR2_X1 i_1609 (.ZN (n_2539), .A1 (n_3288), .A2 (sgo__n168));
NOR2_X1 i_1608 (.ZN (n_2538), .A1 (n_3288), .A2 (n_3270));
NOR2_X1 i_1607 (.ZN (n_2537), .A1 (n_3288), .A2 (n_3271));
NOR2_X1 i_1606 (.ZN (n_2536), .A1 (n_3288), .A2 (n_3272));
NOR2_X1 i_1605 (.ZN (n_2535), .A1 (n_3288), .A2 (n_3273));
NOR2_X1 i_1604 (.ZN (n_2534), .A1 (n_3288), .A2 (n_3274));
NOR2_X1 i_1603 (.ZN (n_2533), .A1 (n_3288), .A2 (n_3275));
NOR2_X1 i_1602 (.ZN (n_2532), .A1 (n_3288), .A2 (n_3276));
NOR2_X1 i_1601 (.ZN (n_2531), .A1 (n_3288), .A2 (n_3277));
NOR2_X1 i_1600 (.ZN (n_2530), .A1 (sgo__n141), .A2 (n_3246));
NOR2_X1 i_1599 (.ZN (n_2529), .A1 (sgo__n141), .A2 (n_3247));
NOR2_X1 i_1598 (.ZN (n_2528), .A1 (sgo__n141), .A2 (n_3248));
NOR2_X1 i_1597 (.ZN (n_2527), .A1 (sgo__n141), .A2 (sgo__n10));
NOR2_X1 i_1596 (.ZN (n_2526), .A1 (sgo__n141), .A2 (n_3250));
NOR2_X1 i_1595 (.ZN (n_2525), .A1 (sgo__n141), .A2 (n_3251));
NOR2_X1 i_1594 (.ZN (n_2524), .A1 (n_3289), .A2 (n_3252));
NOR2_X1 i_1593 (.ZN (n_2523), .A1 (n_3289), .A2 (n_3253));
NOR2_X1 i_1592 (.ZN (n_2522), .A1 (n_3289), .A2 (n_3254));
NOR2_X1 i_1591 (.ZN (n_2521), .A1 (n_3289), .A2 (sgo__n178));
NOR2_X1 i_1590 (.ZN (n_2520), .A1 (n_3289), .A2 (n_3256));
NOR2_X1 i_1589 (.ZN (n_2519), .A1 (n_3289), .A2 (n_3257));
NOR2_X1 i_1588 (.ZN (n_2518), .A1 (n_3289), .A2 (n_3258));
NOR2_X1 i_1587 (.ZN (n_2517), .A1 (n_3289), .A2 (n_3259));
NOR2_X1 i_1586 (.ZN (n_2516), .A1 (n_3289), .A2 (n_3260));
NOR2_X1 i_1585 (.ZN (n_2515), .A1 (n_3289), .A2 (n_3261));
NOR2_X1 i_1584 (.ZN (n_2514), .A1 (n_3289), .A2 (n_3262));
NOR2_X1 i_1583 (.ZN (n_2513), .A1 (n_3289), .A2 (n_3263));
NOR2_X1 i_1582 (.ZN (n_2512), .A1 (n_3289), .A2 (n_3264));
NOR2_X1 i_1581 (.ZN (n_2511), .A1 (n_3289), .A2 (n_3265));
NOR2_X1 i_1580 (.ZN (n_2510), .A1 (sgo__n141), .A2 (n_3266));
NOR2_X1 i_1579 (.ZN (n_2509), .A1 (sgo__n141), .A2 (sgo__n99));
NOR2_X1 i_1578 (.ZN (n_2508), .A1 (sgo__n141), .A2 (sgo__n172));
NOR2_X1 i_1577 (.ZN (n_2507), .A1 (sgo__n141), .A2 (sgo__n168));
NOR2_X1 i_1576 (.ZN (n_2506), .A1 (n_3289), .A2 (n_3270));
NOR2_X1 i_1575 (.ZN (n_2505), .A1 (n_3289), .A2 (n_3271));
NOR2_X1 i_1574 (.ZN (n_2504), .A1 (n_3289), .A2 (n_3272));
NOR2_X1 i_1573 (.ZN (n_2503), .A1 (n_3289), .A2 (n_3273));
NOR2_X1 i_1572 (.ZN (n_2502), .A1 (n_3289), .A2 (n_3274));
NOR2_X1 i_1571 (.ZN (n_2501), .A1 (n_3289), .A2 (n_3275));
NOR2_X1 i_1570 (.ZN (n_2500), .A1 (n_3289), .A2 (n_3276));
NOR2_X1 i_1569 (.ZN (n_2499), .A1 (n_3289), .A2 (n_3277));
NOR2_X1 i_1568 (.ZN (n_2498), .A1 (n_3290), .A2 (n_3246));
NOR2_X1 i_1567 (.ZN (n_2497), .A1 (n_3290), .A2 (n_3247));
NOR2_X1 i_1566 (.ZN (n_2496), .A1 (n_3290), .A2 (n_3248));
NOR2_X1 i_1565 (.ZN (n_2495), .A1 (n_3290), .A2 (n_3249));
NOR2_X1 i_1564 (.ZN (n_2494), .A1 (n_3290), .A2 (n_3250));
NOR2_X1 i_1563 (.ZN (n_2493), .A1 (n_3290), .A2 (n_3251));
NOR2_X1 i_1562 (.ZN (n_2492), .A1 (n_3290), .A2 (n_3252));
NOR2_X1 i_1561 (.ZN (n_2491), .A1 (n_3290), .A2 (n_3253));
NOR2_X1 i_1560 (.ZN (n_2490), .A1 (n_3290), .A2 (n_3254));
NOR2_X1 i_1559 (.ZN (n_2489), .A1 (n_3290), .A2 (sgo__n178));
NOR2_X1 i_1558 (.ZN (n_2488), .A1 (n_3290), .A2 (n_3256));
NOR2_X1 i_1557 (.ZN (n_2487), .A1 (n_3290), .A2 (sgo__n134));
NOR2_X1 i_1556 (.ZN (n_2486), .A1 (n_3290), .A2 (n_3258));
NOR2_X1 i_1555 (.ZN (n_2485), .A1 (n_3290), .A2 (n_3259));
NOR2_X1 i_1554 (.ZN (n_2484), .A1 (n_3290), .A2 (n_3260));
NOR2_X1 i_1553 (.ZN (n_2483), .A1 (n_3290), .A2 (n_3261));
NOR2_X1 i_1552 (.ZN (n_2482), .A1 (n_3290), .A2 (n_3262));
NOR2_X1 i_1551 (.ZN (n_2481), .A1 (n_3290), .A2 (n_3263));
NOR2_X1 i_1550 (.ZN (n_2480), .A1 (n_3290), .A2 (n_3264));
NOR2_X1 i_1549 (.ZN (n_2479), .A1 (n_3290), .A2 (n_3265));
NOR2_X1 i_1548 (.ZN (n_2478), .A1 (n_3290), .A2 (n_3266));
NOR2_X1 i_1547 (.ZN (n_2477), .A1 (n_3290), .A2 (sgo__n99));
NOR2_X1 i_1546 (.ZN (n_2476), .A1 (n_3290), .A2 (sgo__n172));
NOR2_X1 i_1545 (.ZN (n_2475), .A1 (n_3290), .A2 (sgo__n168));
NOR2_X1 i_1544 (.ZN (n_2474), .A1 (n_3290), .A2 (n_3270));
NOR2_X1 i_1543 (.ZN (n_2473), .A1 (n_3290), .A2 (n_3271));
NOR2_X1 i_1542 (.ZN (n_2472), .A1 (n_3290), .A2 (n_3272));
NOR2_X1 i_1541 (.ZN (n_2471), .A1 (n_3290), .A2 (n_3273));
NOR2_X1 i_1540 (.ZN (n_2470), .A1 (n_3290), .A2 (n_3274));
NOR2_X1 i_1539 (.ZN (n_2469), .A1 (n_3290), .A2 (n_3275));
NOR2_X1 i_1538 (.ZN (n_2468), .A1 (n_3290), .A2 (n_3276));
NOR2_X1 i_1537 (.ZN (n_2467), .A1 (n_3290), .A2 (n_3277));
NOR2_X1 i_1536 (.ZN (n_2466), .A1 (n_3291), .A2 (n_3246));
NOR2_X1 i_1535 (.ZN (n_2465), .A1 (n_3291), .A2 (n_3247));
NOR2_X1 i_1534 (.ZN (n_2464), .A1 (n_3291), .A2 (n_3248));
NOR2_X1 i_1533 (.ZN (n_2463), .A1 (n_3291), .A2 (n_3249));
NOR2_X1 i_1532 (.ZN (n_2462), .A1 (n_3291), .A2 (n_3250));
NOR2_X1 i_1531 (.ZN (n_2461), .A1 (n_3291), .A2 (n_3251));
NOR2_X1 i_1530 (.ZN (n_2460), .A1 (n_3291), .A2 (n_3252));
NOR2_X1 i_1529 (.ZN (n_2459), .A1 (n_3291), .A2 (n_3253));
NOR2_X1 i_1528 (.ZN (n_2458), .A1 (n_3291), .A2 (n_3254));
NOR2_X1 i_1527 (.ZN (n_2457), .A1 (n_3291), .A2 (sgo__n178));
NOR2_X1 i_1526 (.ZN (n_2456), .A1 (n_3291), .A2 (n_3256));
NOR2_X1 i_1525 (.ZN (n_2455), .A1 (n_3291), .A2 (n_3257));
NOR2_X1 i_1524 (.ZN (n_2454), .A1 (n_3291), .A2 (n_3258));
NOR2_X1 i_1523 (.ZN (n_2453), .A1 (n_3291), .A2 (n_3259));
NOR2_X1 i_1522 (.ZN (n_2452), .A1 (n_3291), .A2 (n_3260));
NOR2_X1 i_1521 (.ZN (n_2451), .A1 (n_3291), .A2 (n_3261));
NOR2_X1 i_1520 (.ZN (n_2450), .A1 (n_3291), .A2 (n_3262));
NOR2_X1 i_1519 (.ZN (n_2449), .A1 (n_3291), .A2 (n_3263));
NOR2_X1 i_1518 (.ZN (n_2448), .A1 (n_3291), .A2 (n_3264));
NOR2_X1 i_1517 (.ZN (n_2447), .A1 (n_3291), .A2 (sgo__n122));
NOR2_X1 i_1516 (.ZN (n_2446), .A1 (n_3291), .A2 (n_3266));
NOR2_X1 i_1515 (.ZN (n_2445), .A1 (n_3291), .A2 (sgo__n99));
NOR2_X1 i_1514 (.ZN (n_2444), .A1 (n_3291), .A2 (sgo__n172));
NOR2_X1 i_1513 (.ZN (n_2443), .A1 (n_3291), .A2 (sgo__n168));
NOR2_X1 i_1512 (.ZN (n_2442), .A1 (n_3291), .A2 (n_3270));
NOR2_X1 i_1511 (.ZN (n_2441), .A1 (n_3291), .A2 (n_3271));
NOR2_X1 i_1510 (.ZN (n_2440), .A1 (n_3291), .A2 (n_3272));
NOR2_X1 i_1509 (.ZN (n_2439), .A1 (n_3291), .A2 (n_3273));
NOR2_X1 i_1508 (.ZN (n_2438), .A1 (n_3291), .A2 (n_3274));
NOR2_X1 i_1507 (.ZN (n_2437), .A1 (n_3291), .A2 (n_3275));
NOR2_X1 i_1506 (.ZN (n_2436), .A1 (n_3291), .A2 (n_3276));
NOR2_X1 i_1505 (.ZN (n_2435), .A1 (n_3291), .A2 (n_3277));
NOR2_X1 i_1504 (.ZN (n_2434), .A1 (n_3292), .A2 (n_3246));
NOR2_X1 i_1503 (.ZN (n_2433), .A1 (n_3292), .A2 (n_3247));
NOR2_X1 i_1502 (.ZN (n_2432), .A1 (n_3292), .A2 (n_3248));
NOR2_X1 i_1501 (.ZN (n_2431), .A1 (n_3292), .A2 (n_3249));
NOR2_X1 i_1500 (.ZN (n_2430), .A1 (n_3292), .A2 (n_3250));
NOR2_X1 i_1499 (.ZN (n_2429), .A1 (n_3292), .A2 (n_3251));
NOR2_X1 i_1498 (.ZN (n_2428), .A1 (n_3292), .A2 (n_3252));
NOR2_X1 i_1497 (.ZN (n_2427), .A1 (n_3292), .A2 (n_3253));
NOR2_X1 i_1496 (.ZN (n_2426), .A1 (n_3292), .A2 (n_3254));
NOR2_X1 i_1495 (.ZN (n_2425), .A1 (n_3292), .A2 (sgo__n178));
NOR2_X1 i_1494 (.ZN (n_2424), .A1 (n_3292), .A2 (n_3256));
NOR2_X1 i_1493 (.ZN (n_2423), .A1 (n_3292), .A2 (n_3257));
NOR2_X1 i_1492 (.ZN (n_2422), .A1 (n_3292), .A2 (n_3258));
NOR2_X1 i_1491 (.ZN (n_2421), .A1 (n_3292), .A2 (n_3259));
NOR2_X1 i_1490 (.ZN (n_2420), .A1 (n_3292), .A2 (n_3260));
NOR2_X1 i_1489 (.ZN (n_2419), .A1 (n_3292), .A2 (n_3261));
NOR2_X1 i_1488 (.ZN (n_2418), .A1 (n_3292), .A2 (n_3262));
NOR2_X1 i_1487 (.ZN (n_2417), .A1 (n_3292), .A2 (n_3263));
NOR2_X1 i_1486 (.ZN (n_2416), .A1 (n_3292), .A2 (n_3264));
NOR2_X1 i_1485 (.ZN (n_2415), .A1 (n_3292), .A2 (sgo__n122));
NOR2_X1 i_1484 (.ZN (n_2414), .A1 (n_3292), .A2 (n_3266));
NOR2_X1 i_1483 (.ZN (n_2413), .A1 (n_3292), .A2 (sgo__n99));
NOR2_X1 i_1482 (.ZN (n_2412), .A1 (n_3292), .A2 (sgo__n172));
NOR2_X1 i_1481 (.ZN (n_2411), .A1 (n_3292), .A2 (sgo__n168));
NOR2_X1 i_1480 (.ZN (n_2410), .A1 (n_3292), .A2 (n_3270));
NOR2_X1 i_1479 (.ZN (n_2409), .A1 (n_3292), .A2 (n_3271));
NOR2_X1 i_1478 (.ZN (n_2408), .A1 (n_3292), .A2 (n_3272));
NOR2_X1 i_1477 (.ZN (n_2407), .A1 (n_3292), .A2 (n_3273));
NOR2_X1 i_1476 (.ZN (n_2406), .A1 (n_3292), .A2 (n_3274));
NOR2_X1 i_1475 (.ZN (n_2405), .A1 (n_3292), .A2 (n_3275));
NOR2_X1 i_1474 (.ZN (n_2404), .A1 (n_3292), .A2 (n_3276));
NOR2_X1 i_1473 (.ZN (n_2403), .A1 (n_3292), .A2 (n_3277));
NOR2_X1 i_1472 (.ZN (n_2402), .A1 (n_3293), .A2 (n_3246));
NOR2_X1 i_1471 (.ZN (n_2401), .A1 (n_3293), .A2 (n_3247));
NOR2_X1 i_1470 (.ZN (n_2400), .A1 (n_3293), .A2 (n_3248));
NOR2_X1 i_1469 (.ZN (n_2399), .A1 (n_3293), .A2 (n_3249));
NOR2_X1 i_1468 (.ZN (n_2398), .A1 (n_3293), .A2 (n_3250));
NOR2_X1 i_1467 (.ZN (n_2397), .A1 (n_3293), .A2 (n_3251));
NOR2_X1 i_1466 (.ZN (n_2396), .A1 (n_3293), .A2 (n_3252));
NOR2_X1 i_1465 (.ZN (n_2395), .A1 (n_3293), .A2 (n_3253));
NOR2_X1 i_1464 (.ZN (n_2394), .A1 (n_3293), .A2 (n_3254));
NOR2_X1 i_1463 (.ZN (n_2393), .A1 (n_3293), .A2 (sgo__n178));
NOR2_X1 i_1462 (.ZN (n_2392), .A1 (n_3293), .A2 (n_3256));
NOR2_X1 i_1461 (.ZN (n_2391), .A1 (n_3293), .A2 (n_3257));
NOR2_X1 i_1460 (.ZN (n_2390), .A1 (n_3293), .A2 (n_3258));
NOR2_X1 i_1459 (.ZN (n_2389), .A1 (n_3293), .A2 (n_3259));
NOR2_X1 i_1458 (.ZN (n_2388), .A1 (n_3293), .A2 (n_3260));
NOR2_X1 i_1457 (.ZN (n_2387), .A1 (n_3293), .A2 (sgo__n148));
NOR2_X1 i_1456 (.ZN (n_2386), .A1 (n_3293), .A2 (n_3262));
NOR2_X1 i_1455 (.ZN (n_2385), .A1 (n_3293), .A2 (n_3263));
NOR2_X1 i_1454 (.ZN (n_2384), .A1 (n_3293), .A2 (sgo__n195));
NOR2_X1 i_1453 (.ZN (n_2383), .A1 (n_3293), .A2 (sgo__n122));
NOR2_X1 i_1452 (.ZN (n_2382), .A1 (n_3293), .A2 (n_3266));
NOR2_X1 i_1451 (.ZN (n_2381), .A1 (n_3293), .A2 (sgo__n99));
NOR2_X1 i_1450 (.ZN (n_2380), .A1 (n_3293), .A2 (sgo__n172));
NOR2_X1 i_1449 (.ZN (n_2379), .A1 (n_3293), .A2 (sgo__n168));
NOR2_X1 i_1448 (.ZN (n_2378), .A1 (n_3293), .A2 (n_3270));
NOR2_X1 i_1447 (.ZN (n_2377), .A1 (n_3293), .A2 (n_3271));
NOR2_X1 i_1446 (.ZN (n_2376), .A1 (n_3293), .A2 (n_3272));
NOR2_X1 i_1445 (.ZN (n_2375), .A1 (n_3293), .A2 (n_3273));
NOR2_X1 i_1444 (.ZN (n_2374), .A1 (n_3293), .A2 (n_3274));
NOR2_X1 i_1443 (.ZN (n_2373), .A1 (n_3293), .A2 (n_3275));
NOR2_X1 i_1442 (.ZN (n_2372), .A1 (n_3293), .A2 (n_3276));
NOR2_X1 i_1441 (.ZN (n_2371), .A1 (n_3293), .A2 (n_3277));
NOR2_X1 i_1440 (.ZN (n_2370), .A1 (n_3294), .A2 (n_3246));
NOR2_X1 i_1439 (.ZN (n_2369), .A1 (n_3294), .A2 (n_3247));
NOR2_X1 i_1438 (.ZN (n_2368), .A1 (n_3294), .A2 (n_3248));
NOR2_X1 i_1437 (.ZN (n_2367), .A1 (n_3294), .A2 (n_3249));
NOR2_X1 i_1436 (.ZN (n_2366), .A1 (n_3294), .A2 (n_3250));
NOR2_X1 i_1435 (.ZN (n_2365), .A1 (n_3294), .A2 (n_3251));
NOR2_X1 i_1434 (.ZN (n_2364), .A1 (n_3294), .A2 (n_3252));
NOR2_X1 i_1433 (.ZN (n_2363), .A1 (n_3294), .A2 (n_3253));
NOR2_X1 i_1432 (.ZN (n_2362), .A1 (n_3294), .A2 (n_3254));
NOR2_X1 i_1431 (.ZN (n_2361), .A1 (n_3294), .A2 (n_3255));
NOR2_X1 i_1430 (.ZN (n_2360), .A1 (n_3294), .A2 (n_3256));
NOR2_X1 i_1429 (.ZN (n_2359), .A1 (n_3294), .A2 (n_3257));
NOR2_X1 i_1428 (.ZN (n_2358), .A1 (n_3294), .A2 (n_3258));
NOR2_X1 i_1427 (.ZN (n_2357), .A1 (n_3294), .A2 (n_3259));
NOR2_X1 i_1426 (.ZN (n_2356), .A1 (n_3294), .A2 (n_3260));
NOR2_X1 i_1425 (.ZN (n_2355), .A1 (n_3294), .A2 (sgo__n150));
NOR2_X1 i_1424 (.ZN (n_2354), .A1 (n_3294), .A2 (n_3262));
NOR2_X1 i_1423 (.ZN (n_2353), .A1 (n_3294), .A2 (n_3263));
NOR2_X1 i_1422 (.ZN (n_2352), .A1 (n_3294), .A2 (sgo__n195));
NOR2_X1 i_1421 (.ZN (n_2351), .A1 (n_3294), .A2 (sgo__n122));
NOR2_X1 i_1420 (.ZN (n_2350), .A1 (n_3294), .A2 (n_3266));
NOR2_X1 i_1419 (.ZN (n_2349), .A1 (n_3294), .A2 (sgo__n99));
NOR2_X1 i_1418 (.ZN (n_2348), .A1 (n_3294), .A2 (sgo__n172));
NOR2_X1 i_1417 (.ZN (n_2347), .A1 (n_3294), .A2 (n_3269));
NOR2_X1 i_1416 (.ZN (n_2346), .A1 (n_3294), .A2 (n_3270));
NOR2_X1 i_1415 (.ZN (n_2345), .A1 (n_3294), .A2 (n_3271));
NOR2_X1 i_1414 (.ZN (n_2344), .A1 (n_3294), .A2 (n_3272));
NOR2_X1 i_1413 (.ZN (n_2343), .A1 (n_3294), .A2 (n_3273));
NOR2_X1 i_1412 (.ZN (n_2342), .A1 (n_3294), .A2 (n_3274));
NOR2_X1 i_1411 (.ZN (n_2341), .A1 (n_3294), .A2 (n_3275));
NOR2_X1 i_1410 (.ZN (n_2340), .A1 (n_3294), .A2 (n_3276));
NOR2_X1 i_1409 (.ZN (n_2339), .A1 (n_3294), .A2 (n_3277));
NOR2_X1 i_1408 (.ZN (n_2338), .A1 (n_3295), .A2 (n_3246));
NOR2_X1 i_1407 (.ZN (n_2337), .A1 (n_3295), .A2 (n_3247));
NOR2_X1 i_1406 (.ZN (n_2336), .A1 (n_3295), .A2 (n_3248));
NOR2_X1 i_1405 (.ZN (n_2335), .A1 (n_3295), .A2 (n_3249));
NOR2_X1 i_1404 (.ZN (n_2334), .A1 (n_3295), .A2 (n_3250));
NOR2_X1 i_1403 (.ZN (n_2333), .A1 (n_3295), .A2 (n_3251));
NOR2_X1 i_1402 (.ZN (n_2332), .A1 (n_3295), .A2 (n_3252));
NOR2_X1 i_1401 (.ZN (n_2331), .A1 (n_3295), .A2 (n_3253));
NOR2_X1 i_1400 (.ZN (n_2330), .A1 (n_3295), .A2 (n_3254));
NOR2_X1 i_1399 (.ZN (n_2329), .A1 (n_3295), .A2 (n_3255));
NOR2_X1 i_1398 (.ZN (n_2328), .A1 (n_3295), .A2 (n_3256));
NOR2_X1 i_1397 (.ZN (n_2327), .A1 (n_3295), .A2 (n_3257));
NOR2_X1 i_1396 (.ZN (n_2326), .A1 (n_3295), .A2 (n_3258));
NOR2_X1 i_1395 (.ZN (n_2325), .A1 (n_3295), .A2 (n_3259));
NOR2_X1 i_1394 (.ZN (n_2324), .A1 (sgo__n78), .A2 (n_3260));
NOR2_X1 i_1393 (.ZN (n_2323), .A1 (sgo__n78), .A2 (sgo__n150));
NOR2_X1 i_1392 (.ZN (n_2322), .A1 (sgo__n78), .A2 (sgo__n176));
NOR2_X1 i_1391 (.ZN (n_2321), .A1 (sgo__n78), .A2 (sgo__n162));
NOR2_X1 i_1390 (.ZN (n_2320), .A1 (sgo__n78), .A2 (sgo__n195));
NOR2_X1 i_1389 (.ZN (n_2319), .A1 (sgo__n78), .A2 (sgo__n122));
NOR2_X1 i_1388 (.ZN (n_2318), .A1 (sgo__n78), .A2 (n_3266));
NOR2_X1 i_1387 (.ZN (n_2317), .A1 (sgo__n78), .A2 (sgo__n99));
NOR2_X1 i_1386 (.ZN (n_2316), .A1 (sgo__n78), .A2 (sgo__n172));
NOR2_X1 i_1385 (.ZN (n_2315), .A1 (sgo__n78), .A2 (n_3269));
NOR2_X1 i_1384 (.ZN (n_2314), .A1 (sgo__n78), .A2 (n_3270));
NOR2_X1 i_1383 (.ZN (n_2313), .A1 (sgo__n78), .A2 (n_3271));
NOR2_X1 i_1382 (.ZN (n_2312), .A1 (n_3295), .A2 (n_3272));
NOR2_X1 i_1381 (.ZN (n_2311), .A1 (n_3295), .A2 (n_3273));
NOR2_X1 i_1380 (.ZN (n_2310), .A1 (n_3295), .A2 (n_3274));
NOR2_X1 i_1379 (.ZN (n_2309), .A1 (n_3295), .A2 (n_3275));
NOR2_X1 i_1378 (.ZN (n_2308), .A1 (n_3295), .A2 (n_3276));
NOR2_X1 i_1377 (.ZN (n_2307), .A1 (n_3295), .A2 (n_3277));
NOR2_X1 i_1376 (.ZN (n_2306), .A1 (n_3296), .A2 (n_3246));
NOR2_X1 i_1375 (.ZN (n_2305), .A1 (n_3296), .A2 (n_3247));
NOR2_X1 i_1374 (.ZN (n_2304), .A1 (n_3296), .A2 (n_3248));
NOR2_X1 i_1373 (.ZN (n_2303), .A1 (n_3296), .A2 (n_3249));
NOR2_X1 i_1372 (.ZN (n_2302), .A1 (n_3296), .A2 (n_3250));
NOR2_X1 i_1371 (.ZN (n_2301), .A1 (n_3296), .A2 (n_3251));
NOR2_X1 i_1370 (.ZN (n_2300), .A1 (n_3296), .A2 (n_3252));
NOR2_X1 i_1369 (.ZN (n_2299), .A1 (n_3296), .A2 (n_3253));
NOR2_X1 i_1368 (.ZN (n_2298), .A1 (n_3296), .A2 (n_3254));
NOR2_X1 i_1367 (.ZN (n_2297), .A1 (n_3296), .A2 (n_3255));
NOR2_X1 i_1366 (.ZN (n_2296), .A1 (n_3296), .A2 (n_3256));
NOR2_X1 i_1365 (.ZN (n_2295), .A1 (n_3296), .A2 (n_3257));
NOR2_X1 i_1364 (.ZN (n_2294), .A1 (n_3296), .A2 (n_3258));
NOR2_X1 i_1363 (.ZN (n_2293), .A1 (n_3296), .A2 (n_3259));
NOR2_X1 i_1362 (.ZN (n_2292), .A1 (sgo__n98), .A2 (n_3260));
NOR2_X1 i_1361 (.ZN (n_2291), .A1 (sgo__n98), .A2 (sgo__n147));
NOR2_X1 i_1360 (.ZN (n_2290), .A1 (sgo__n98), .A2 (sgo__n176));
NOR2_X1 i_1359 (.ZN (n_2289), .A1 (sgo__n98), .A2 (sgo__n162));
NOR2_X1 i_1358 (.ZN (n_2288), .A1 (sgo__n98), .A2 (sgo__n195));
NOR2_X1 i_1357 (.ZN (n_2287), .A1 (sgo__n98), .A2 (sgo__n122));
NOR2_X1 i_1356 (.ZN (n_2286), .A1 (sgo__n98), .A2 (n_3266));
NOR2_X1 i_1355 (.ZN (n_2285), .A1 (sgo__n98), .A2 (sgo__n99));
NOR2_X1 i_1354 (.ZN (n_2284), .A1 (sgo__n98), .A2 (sgo__n172));
NOR2_X1 i_1353 (.ZN (n_2283), .A1 (sgo__n98), .A2 (n_3269));
NOR2_X1 i_1352 (.ZN (n_2282), .A1 (sgo__n98), .A2 (n_3270));
NOR2_X1 i_1351 (.ZN (n_2281), .A1 (sgo__n98), .A2 (n_3271));
NOR2_X1 i_1350 (.ZN (n_2280), .A1 (sgo__n98), .A2 (n_3272));
NOR2_X1 i_1349 (.ZN (n_2279), .A1 (n_3296), .A2 (n_3273));
NOR2_X1 i_1348 (.ZN (n_2278), .A1 (sgo__n98), .A2 (n_3274));
NOR2_X1 i_1347 (.ZN (n_2277), .A1 (n_3296), .A2 (n_3275));
NOR2_X1 i_1346 (.ZN (n_2276), .A1 (n_3296), .A2 (n_3276));
NOR2_X1 i_1345 (.ZN (n_2275), .A1 (n_3296), .A2 (n_3277));
NOR2_X1 i_1344 (.ZN (n_2274), .A1 (n_3297), .A2 (n_3246));
NOR2_X1 i_1343 (.ZN (n_2273), .A1 (n_3297), .A2 (n_3247));
NOR2_X1 i_1342 (.ZN (n_2272), .A1 (n_3297), .A2 (n_3248));
NOR2_X1 i_1341 (.ZN (n_2271), .A1 (n_3297), .A2 (n_3249));
NOR2_X1 i_1340 (.ZN (n_2270), .A1 (n_3297), .A2 (n_3250));
NOR2_X1 i_1339 (.ZN (n_2269), .A1 (n_3297), .A2 (n_3251));
NOR2_X1 i_1338 (.ZN (n_2268), .A1 (n_3297), .A2 (n_3252));
NOR2_X1 i_1337 (.ZN (n_2267), .A1 (n_3297), .A2 (n_3253));
NOR2_X1 i_1336 (.ZN (n_2266), .A1 (n_3297), .A2 (n_3254));
NOR2_X1 i_1335 (.ZN (n_2265), .A1 (n_3297), .A2 (n_3255));
NOR2_X1 i_1334 (.ZN (n_2264), .A1 (n_3297), .A2 (n_3256));
NOR2_X1 i_1333 (.ZN (n_2263), .A1 (n_3297), .A2 (n_3257));
NOR2_X1 i_1332 (.ZN (n_2262), .A1 (n_3297), .A2 (n_3258));
NOR2_X1 i_1331 (.ZN (n_2261), .A1 (n_3297), .A2 (n_3259));
NOR2_X1 i_1330 (.ZN (n_2260), .A1 (sgo__n43), .A2 (sgo__n201));
NOR2_X1 i_1329 (.ZN (n_2259), .A1 (sgo__n43), .A2 (sgo__n147));
NOR2_X1 i_1328 (.ZN (n_2258), .A1 (sgo__n43), .A2 (sgo__n176));
NOR2_X1 i_1327 (.ZN (n_2257), .A1 (sgo__n43), .A2 (sgo__n162));
NOR2_X1 i_1326 (.ZN (n_2256), .A1 (sgo__n43), .A2 (sgo__n195));
NOR2_X1 i_1325 (.ZN (n_2255), .A1 (sgo__n43), .A2 (sgo__n122));
NOR2_X1 i_1324 (.ZN (n_2254), .A1 (sgo__n43), .A2 (n_3266));
NOR2_X1 i_1323 (.ZN (n_2253), .A1 (sgo__n43), .A2 (sgo__n99));
NOR2_X1 i_1322 (.ZN (n_2252), .A1 (sgo__n43), .A2 (sgo__n172));
NOR2_X1 i_1321 (.ZN (n_2251), .A1 (sgo__n43), .A2 (n_3269));
NOR2_X1 i_1320 (.ZN (n_2250), .A1 (sgo__n43), .A2 (n_3270));
NOR2_X1 i_1319 (.ZN (n_2249), .A1 (sgo__n43), .A2 (n_3271));
NOR2_X1 i_1318 (.ZN (n_2248), .A1 (n_3297), .A2 (n_3272));
NOR2_X1 i_1317 (.ZN (n_2247), .A1 (sgo__n43), .A2 (n_3273));
NOR2_X1 i_1316 (.ZN (n_2246), .A1 (n_3297), .A2 (n_3274));
NOR2_X1 i_1315 (.ZN (n_2245), .A1 (n_3297), .A2 (n_3275));
NOR2_X1 i_1314 (.ZN (n_2244), .A1 (n_3297), .A2 (n_3276));
NOR2_X1 i_1313 (.ZN (n_2243), .A1 (n_3297), .A2 (n_3277));
NOR2_X1 i_1312 (.ZN (n_2242), .A1 (sgo__n5), .A2 (n_3246));
NOR2_X1 i_1311 (.ZN (n_2241), .A1 (sgo__n5), .A2 (n_3247));
NOR2_X1 i_1310 (.ZN (n_2240), .A1 (sgo__n5), .A2 (n_3248));
NOR2_X1 i_1309 (.ZN (n_2239), .A1 (sgo__n5), .A2 (n_3249));
NOR2_X1 i_1308 (.ZN (n_2238), .A1 (sgo__n5), .A2 (n_3250));
NOR2_X1 i_1307 (.ZN (n_2237), .A1 (n_3298), .A2 (n_3251));
NOR2_X1 i_1306 (.ZN (n_2236), .A1 (n_3298), .A2 (n_3252));
NOR2_X1 i_1305 (.ZN (n_2235), .A1 (n_3298), .A2 (n_3253));
NOR2_X1 i_1304 (.ZN (n_2234), .A1 (n_3298), .A2 (n_3254));
NOR2_X1 i_1303 (.ZN (n_2233), .A1 (n_3298), .A2 (sgo__n180));
NOR2_X1 i_1302 (.ZN (n_2232), .A1 (sgo__n3), .A2 (sgo__n182));
NOR2_X1 i_1301 (.ZN (n_2231), .A1 (sgo__n3), .A2 (n_3257));
NOR2_X1 i_1300 (.ZN (n_2230), .A1 (sgo__n3), .A2 (n_3258));
NOR2_X1 i_1299 (.ZN (n_2229), .A1 (sgo__n3), .A2 (sgo__n174));
NOR2_X1 i_1298 (.ZN (n_2228), .A1 (sgo__n3), .A2 (sgo__n201));
NOR2_X1 i_1297 (.ZN (n_2227), .A1 (sgo__n3), .A2 (sgo__n147));
NOR2_X1 i_1296 (.ZN (n_2226), .A1 (sgo__n3), .A2 (sgo__n176));
NOR2_X1 i_1295 (.ZN (n_2225), .A1 (sgo__n3), .A2 (sgo__n162));
NOR2_X1 i_1294 (.ZN (n_2224), .A1 (sgo__n3), .A2 (sgo__n195));
NOR2_X1 i_1293 (.ZN (n_2223), .A1 (sgo__n3), .A2 (sgo__n122));
NOR2_X1 i_1292 (.ZN (n_2222), .A1 (sgo__n3), .A2 (n_3266));
NOR2_X1 i_1291 (.ZN (n_2221), .A1 (sgo__n3), .A2 (sgo__n99));
NOR2_X1 i_1290 (.ZN (n_2220), .A1 (sgo__n3), .A2 (sgo__n172));
NOR2_X1 i_1289 (.ZN (n_2219), .A1 (sgo__n3), .A2 (n_3269));
NOR2_X1 i_1288 (.ZN (n_2218), .A1 (sgo__n3), .A2 (n_3270));
NOR2_X1 i_1287 (.ZN (n_2217), .A1 (n_3298), .A2 (n_3271));
NOR2_X1 i_1286 (.ZN (n_2216), .A1 (n_3298), .A2 (n_3272));
NOR2_X1 i_1285 (.ZN (n_2215), .A1 (n_3298), .A2 (n_3273));
NOR2_X1 i_1284 (.ZN (n_2214), .A1 (n_3298), .A2 (n_3274));
NOR2_X1 i_1283 (.ZN (n_2213), .A1 (n_3298), .A2 (n_3275));
NOR2_X1 i_1282 (.ZN (n_2212), .A1 (n_3298), .A2 (n_3276));
NOR2_X1 i_1281 (.ZN (n_2211), .A1 (n_3298), .A2 (n_3277));
NOR2_X1 i_1280 (.ZN (n_2210), .A1 (n_3299), .A2 (n_3246));
NOR2_X1 i_1279 (.ZN (n_2209), .A1 (n_3299), .A2 (n_3247));
NOR2_X1 i_1278 (.ZN (n_2208), .A1 (n_3299), .A2 (n_3248));
NOR2_X1 i_1277 (.ZN (n_2207), .A1 (n_3299), .A2 (n_3249));
NOR2_X1 i_1276 (.ZN (n_2206), .A1 (n_3299), .A2 (n_3250));
NOR2_X1 i_1275 (.ZN (n_2205), .A1 (n_3299), .A2 (n_3251));
NOR2_X1 i_1274 (.ZN (n_2204), .A1 (n_3299), .A2 (n_3252));
NOR2_X1 i_1273 (.ZN (n_2203), .A1 (n_3299), .A2 (n_3253));
NOR2_X1 i_1272 (.ZN (n_2202), .A1 (n_3299), .A2 (n_3254));
NOR2_X1 i_1271 (.ZN (n_2201), .A1 (n_3299), .A2 (n_3255));
NOR2_X1 i_1270 (.ZN (n_2200), .A1 (n_3299), .A2 (sgo__n182));
NOR2_X1 i_1269 (.ZN (n_2199), .A1 (n_3299), .A2 (n_3257));
NOR2_X1 i_1268 (.ZN (n_2198), .A1 (n_3299), .A2 (n_3258));
NOR2_X1 i_1267 (.ZN (n_2197), .A1 (n_3299), .A2 (sgo__n174));
NOR2_X1 i_1266 (.ZN (n_2196), .A1 (n_3299), .A2 (sgo__n201));
NOR2_X1 i_1265 (.ZN (n_2195), .A1 (n_3299), .A2 (sgo__n147));
NOR2_X1 i_1264 (.ZN (n_2194), .A1 (n_3299), .A2 (sgo__n176));
NOR2_X1 i_1263 (.ZN (n_2193), .A1 (n_3299), .A2 (sgo__n162));
NOR2_X1 i_1262 (.ZN (n_2192), .A1 (n_3299), .A2 (sgo__n195));
NOR2_X1 i_1261 (.ZN (n_2191), .A1 (n_3299), .A2 (sgo__n122));
NOR2_X1 i_1260 (.ZN (n_2190), .A1 (n_3299), .A2 (n_3266));
NOR2_X1 i_1259 (.ZN (n_2189), .A1 (n_3299), .A2 (sgo__n99));
NOR2_X1 i_1258 (.ZN (n_2188), .A1 (n_3299), .A2 (n_3268));
NOR2_X1 i_1257 (.ZN (n_2187), .A1 (n_3299), .A2 (n_3269));
NOR2_X1 i_1256 (.ZN (n_2186), .A1 (n_3299), .A2 (n_3270));
NOR2_X1 i_1255 (.ZN (n_2185), .A1 (n_3299), .A2 (n_3271));
NOR2_X1 i_1254 (.ZN (n_2184), .A1 (n_3299), .A2 (n_3272));
NOR2_X1 i_1253 (.ZN (n_2183), .A1 (n_3299), .A2 (n_3273));
NOR2_X1 i_1252 (.ZN (n_2182), .A1 (n_3299), .A2 (n_3274));
NOR2_X1 i_1251 (.ZN (n_2181), .A1 (n_3299), .A2 (n_3275));
NOR2_X1 i_1250 (.ZN (n_2180), .A1 (n_3299), .A2 (n_3276));
NOR2_X1 i_1249 (.ZN (n_2179), .A1 (n_3299), .A2 (n_3277));
NOR2_X1 i_1248 (.ZN (n_2178), .A1 (n_3300), .A2 (n_3246));
NOR2_X1 i_1247 (.ZN (n_2177), .A1 (n_3300), .A2 (n_3247));
NOR2_X1 i_1246 (.ZN (n_2176), .A1 (n_3300), .A2 (n_3248));
NOR2_X1 i_1245 (.ZN (n_2175), .A1 (n_3300), .A2 (n_3249));
NOR2_X1 i_1244 (.ZN (n_2174), .A1 (n_3300), .A2 (n_3250));
NOR2_X1 i_1243 (.ZN (n_2173), .A1 (n_3300), .A2 (n_3251));
NOR2_X1 i_1242 (.ZN (n_2172), .A1 (n_3300), .A2 (n_3252));
NOR2_X1 i_1241 (.ZN (n_2171), .A1 (n_3300), .A2 (n_3253));
NOR2_X1 i_1240 (.ZN (n_2170), .A1 (n_3300), .A2 (n_3254));
NOR2_X1 i_1239 (.ZN (n_2169), .A1 (n_3300), .A2 (n_3255));
NOR2_X1 i_1238 (.ZN (n_2168), .A1 (n_3300), .A2 (sgo__n182));
NOR2_X1 i_1237 (.ZN (n_2167), .A1 (n_3300), .A2 (n_3257));
NOR2_X1 i_1236 (.ZN (n_2166), .A1 (n_3300), .A2 (n_3258));
NOR2_X1 i_1235 (.ZN (n_2165), .A1 (n_3300), .A2 (sgo__n174));
NOR2_X1 i_1234 (.ZN (n_2164), .A1 (n_3300), .A2 (sgo__n201));
NOR2_X1 i_1233 (.ZN (n_2163), .A1 (n_3300), .A2 (sgo__n147));
NOR2_X1 i_1232 (.ZN (n_2162), .A1 (n_3300), .A2 (sgo__n176));
NOR2_X1 i_1231 (.ZN (n_2161), .A1 (n_3300), .A2 (sgo__n162));
NOR2_X1 i_1230 (.ZN (n_2160), .A1 (n_3300), .A2 (sgo__n195));
NOR2_X1 i_1229 (.ZN (n_2159), .A1 (n_3300), .A2 (sgo__n122));
NOR2_X1 i_1228 (.ZN (n_2158), .A1 (n_3300), .A2 (n_3266));
NOR2_X1 i_1227 (.ZN (n_2157), .A1 (n_3300), .A2 (sgo__n99));
NOR2_X1 i_1226 (.ZN (n_2156), .A1 (n_3300), .A2 (n_3268));
NOR2_X1 i_1225 (.ZN (n_2155), .A1 (n_3300), .A2 (n_3269));
NOR2_X1 i_1224 (.ZN (n_2154), .A1 (n_3300), .A2 (n_3270));
NOR2_X1 i_1223 (.ZN (n_2153), .A1 (n_3300), .A2 (n_3271));
NOR2_X1 i_1222 (.ZN (n_2152), .A1 (n_3300), .A2 (n_3272));
NOR2_X1 i_1221 (.ZN (n_2151), .A1 (n_3300), .A2 (n_3273));
NOR2_X1 i_1220 (.ZN (n_2150), .A1 (n_3300), .A2 (n_3274));
NOR2_X1 i_1219 (.ZN (n_2149), .A1 (n_3300), .A2 (n_3275));
NOR2_X1 i_1218 (.ZN (n_2148), .A1 (n_3300), .A2 (n_3276));
NOR2_X1 i_1217 (.ZN (n_2147), .A1 (n_3300), .A2 (n_3277));
NOR2_X1 i_1216 (.ZN (n_2146), .A1 (n_3301), .A2 (n_3246));
NOR2_X1 i_1215 (.ZN (n_2145), .A1 (n_3301), .A2 (n_3247));
NOR2_X1 i_1214 (.ZN (n_2144), .A1 (n_3301), .A2 (n_3248));
NOR2_X1 i_1213 (.ZN (n_2143), .A1 (n_3301), .A2 (n_3249));
NOR2_X1 i_1212 (.ZN (n_2142), .A1 (n_3301), .A2 (n_3250));
NOR2_X1 i_1211 (.ZN (n_2141), .A1 (sgo__n19), .A2 (n_3251));
NOR2_X1 i_1210 (.ZN (n_2140), .A1 (n_3301), .A2 (n_3252));
NOR2_X1 i_1209 (.ZN (n_2139), .A1 (sgo__n19), .A2 (n_3253));
NOR2_X1 i_1208 (.ZN (n_2138), .A1 (sgo__n19), .A2 (n_3254));
NOR2_X1 i_1207 (.ZN (n_2137), .A1 (sgo__n19), .A2 (n_3255));
NOR2_X1 i_1206 (.ZN (n_2136), .A1 (sgo__n19), .A2 (sgo__n182));
NOR2_X1 i_1205 (.ZN (n_2135), .A1 (sgo__n19), .A2 (n_3257));
NOR2_X1 i_1204 (.ZN (n_2134), .A1 (sgo__n19), .A2 (n_3258));
NOR2_X1 i_1203 (.ZN (n_2133), .A1 (sgo__n19), .A2 (sgo__n174));
NOR2_X1 i_1202 (.ZN (n_2132), .A1 (sgo__n19), .A2 (sgo__n201));
NOR2_X1 i_1201 (.ZN (n_2131), .A1 (sgo__n19), .A2 (sgo__n147));
NOR2_X1 i_1200 (.ZN (n_2130), .A1 (sgo__n19), .A2 (sgo__n176));
NOR2_X1 i_1199 (.ZN (n_2129), .A1 (sgo__n19), .A2 (sgo__n162));
NOR2_X1 i_1198 (.ZN (n_2128), .A1 (sgo__n19), .A2 (sgo__n195));
NOR2_X1 i_1197 (.ZN (n_2127), .A1 (sgo__n19), .A2 (sgo__n122));
NOR2_X1 i_1196 (.ZN (n_2126), .A1 (sgo__n19), .A2 (n_3266));
NOR2_X1 i_1195 (.ZN (n_2125), .A1 (sgo__n19), .A2 (sgo__n99));
NOR2_X1 i_1194 (.ZN (n_2124), .A1 (n_3301), .A2 (n_3268));
NOR2_X1 i_1193 (.ZN (n_2123), .A1 (n_3301), .A2 (n_3269));
NOR2_X1 i_1192 (.ZN (n_2122), .A1 (n_3301), .A2 (n_3270));
NOR2_X1 i_1191 (.ZN (n_2121), .A1 (n_3301), .A2 (n_3271));
NOR2_X1 i_1190 (.ZN (n_2120), .A1 (n_3301), .A2 (n_3272));
NOR2_X1 i_1189 (.ZN (n_2119), .A1 (n_3301), .A2 (n_3273));
NOR2_X1 i_1188 (.ZN (n_2118), .A1 (n_3301), .A2 (n_3274));
NOR2_X1 i_1187 (.ZN (n_2117), .A1 (n_3301), .A2 (n_3275));
NOR2_X1 i_1186 (.ZN (n_2116), .A1 (n_3301), .A2 (n_3276));
NOR2_X1 i_1185 (.ZN (n_2115), .A1 (n_3301), .A2 (n_3277));
NOR2_X1 i_1184 (.ZN (n_2114), .A1 (n_3302), .A2 (n_3246));
NOR2_X1 i_1183 (.ZN (n_2113), .A1 (n_3302), .A2 (n_3247));
NOR2_X1 i_1182 (.ZN (n_2112), .A1 (n_3302), .A2 (n_3248));
NOR2_X1 i_1181 (.ZN (n_2111), .A1 (n_3302), .A2 (n_3249));
NOR2_X1 i_1180 (.ZN (n_2110), .A1 (n_3302), .A2 (n_3250));
NOR2_X1 i_1179 (.ZN (n_2109), .A1 (n_3302), .A2 (n_3251));
NOR2_X1 i_1178 (.ZN (n_2108), .A1 (n_3302), .A2 (n_3252));
NOR2_X1 i_1177 (.ZN (n_2107), .A1 (n_3302), .A2 (n_3253));
NOR2_X1 i_1176 (.ZN (n_2106), .A1 (n_3302), .A2 (n_3254));
NOR2_X1 i_1175 (.ZN (n_2105), .A1 (n_3302), .A2 (n_3255));
NOR2_X1 i_1174 (.ZN (n_2104), .A1 (n_3302), .A2 (sgo__n182));
NOR2_X1 i_1173 (.ZN (n_2103), .A1 (n_3302), .A2 (n_3257));
NOR2_X1 i_1172 (.ZN (n_2102), .A1 (n_3302), .A2 (n_3258));
NOR2_X1 i_1171 (.ZN (n_2101), .A1 (n_3302), .A2 (sgo__n174));
NOR2_X1 i_1170 (.ZN (n_2100), .A1 (n_3302), .A2 (sgo__n201));
NOR2_X1 i_1169 (.ZN (n_2099), .A1 (n_3302), .A2 (sgo__n147));
NOR2_X1 i_1168 (.ZN (n_2098), .A1 (n_3302), .A2 (sgo__n176));
NOR2_X1 i_1167 (.ZN (n_2097), .A1 (n_3302), .A2 (sgo__n162));
NOR2_X1 i_1166 (.ZN (n_2096), .A1 (n_3302), .A2 (sgo__n195));
NOR2_X1 i_1165 (.ZN (n_2095), .A1 (n_3302), .A2 (sgo__n122));
NOR2_X1 i_1164 (.ZN (n_2094), .A1 (n_3302), .A2 (n_3266));
NOR2_X1 i_1163 (.ZN (n_2093), .A1 (n_3302), .A2 (n_3267));
NOR2_X1 i_1162 (.ZN (n_2092), .A1 (n_3302), .A2 (n_3268));
NOR2_X1 i_1161 (.ZN (n_2091), .A1 (n_3302), .A2 (n_3269));
NOR2_X1 i_1160 (.ZN (n_2090), .A1 (n_3302), .A2 (n_3270));
NOR2_X1 i_1159 (.ZN (n_2089), .A1 (n_3302), .A2 (n_3271));
NOR2_X1 i_1158 (.ZN (n_2088), .A1 (n_3302), .A2 (n_3272));
NOR2_X1 i_1157 (.ZN (n_2087), .A1 (n_3302), .A2 (n_3273));
NOR2_X1 i_1156 (.ZN (n_2086), .A1 (n_3302), .A2 (n_3274));
NOR2_X1 i_1155 (.ZN (n_2085), .A1 (n_3302), .A2 (n_3275));
NOR2_X1 i_1154 (.ZN (n_2084), .A1 (n_3302), .A2 (n_3276));
NOR2_X1 i_1153 (.ZN (n_2083), .A1 (n_3302), .A2 (n_3277));
NOR2_X1 i_1152 (.ZN (n_2082), .A1 (n_3303), .A2 (n_3246));
NOR2_X1 i_1151 (.ZN (n_2081), .A1 (n_3303), .A2 (n_3247));
NOR2_X1 i_1150 (.ZN (n_2080), .A1 (n_3303), .A2 (n_3248));
NOR2_X1 i_1149 (.ZN (n_2079), .A1 (n_3303), .A2 (n_3249));
NOR2_X1 i_1148 (.ZN (n_2078), .A1 (n_3303), .A2 (n_3250));
NOR2_X1 i_1147 (.ZN (n_2077), .A1 (n_3303), .A2 (n_3251));
NOR2_X1 i_1146 (.ZN (n_2076), .A1 (n_3303), .A2 (n_3252));
NOR2_X1 i_1145 (.ZN (n_2075), .A1 (n_3303), .A2 (n_3253));
NOR2_X1 i_1144 (.ZN (n_2074), .A1 (n_3303), .A2 (n_3254));
NOR2_X1 i_1143 (.ZN (n_2073), .A1 (n_3303), .A2 (n_3255));
NOR2_X1 i_1142 (.ZN (n_2072), .A1 (n_3303), .A2 (sgo__n182));
NOR2_X1 i_1141 (.ZN (n_2071), .A1 (n_3303), .A2 (n_3257));
NOR2_X1 i_1140 (.ZN (n_2070), .A1 (n_3303), .A2 (n_3258));
NOR2_X1 i_1139 (.ZN (n_2069), .A1 (n_3303), .A2 (sgo__n174));
NOR2_X1 i_1138 (.ZN (n_2068), .A1 (n_3303), .A2 (sgo__n201));
NOR2_X1 i_1137 (.ZN (n_2067), .A1 (n_3303), .A2 (sgo__n147));
NOR2_X1 i_1136 (.ZN (n_2066), .A1 (n_3303), .A2 (sgo__n176));
NOR2_X1 i_1135 (.ZN (n_2065), .A1 (n_3303), .A2 (sgo__n162));
NOR2_X1 i_1134 (.ZN (n_2064), .A1 (n_3303), .A2 (n_3264));
NOR2_X1 i_1133 (.ZN (n_2063), .A1 (n_3303), .A2 (n_3265));
NOR2_X1 i_1132 (.ZN (n_2062), .A1 (n_3303), .A2 (n_3266));
NOR2_X1 i_1131 (.ZN (n_2061), .A1 (n_3303), .A2 (n_3267));
NOR2_X1 i_1130 (.ZN (n_2060), .A1 (n_3303), .A2 (n_3268));
NOR2_X1 i_1129 (.ZN (n_2059), .A1 (n_3303), .A2 (n_3269));
NOR2_X1 i_1128 (.ZN (n_2058), .A1 (n_3303), .A2 (n_3270));
NOR2_X1 i_1127 (.ZN (n_2057), .A1 (n_3303), .A2 (n_3271));
NOR2_X1 i_1126 (.ZN (n_2056), .A1 (n_3303), .A2 (n_3272));
NOR2_X1 i_1125 (.ZN (n_2055), .A1 (n_3303), .A2 (n_3273));
NOR2_X1 i_1124 (.ZN (n_2054), .A1 (n_3303), .A2 (n_3274));
NOR2_X1 i_1123 (.ZN (n_2053), .A1 (n_3303), .A2 (n_3275));
NOR2_X1 i_1122 (.ZN (n_2052), .A1 (n_3303), .A2 (n_3276));
NOR2_X1 i_1121 (.ZN (n_2051), .A1 (n_3303), .A2 (n_3277));
NOR2_X1 i_1120 (.ZN (n_2050), .A1 (n_3304), .A2 (n_3246));
NOR2_X1 i_1119 (.ZN (n_2049), .A1 (n_3304), .A2 (n_3247));
NOR2_X1 i_1118 (.ZN (n_2048), .A1 (sgo__n109), .A2 (n_3248));
NOR2_X1 i_1117 (.ZN (n_2047), .A1 (sgo__n109), .A2 (n_3249));
NOR2_X1 i_1116 (.ZN (n_2046), .A1 (sgo__n109), .A2 (n_3250));
NOR2_X1 i_1115 (.ZN (n_2045), .A1 (sgo__n109), .A2 (n_3251));
NOR2_X1 i_1114 (.ZN (n_2044), .A1 (sgo__n109), .A2 (n_3252));
NOR2_X1 i_1113 (.ZN (n_2043), .A1 (sgo__n109), .A2 (n_3253));
NOR2_X1 i_1112 (.ZN (n_2042), .A1 (sgo__n109), .A2 (n_3254));
NOR2_X1 i_1111 (.ZN (n_2041), .A1 (sgo__n109), .A2 (n_3255));
NOR2_X1 i_1110 (.ZN (n_2040), .A1 (sgo__n109), .A2 (sgo__n182));
NOR2_X1 i_1109 (.ZN (n_2039), .A1 (sgo__n109), .A2 (n_3257));
NOR2_X1 i_1108 (.ZN (n_2038), .A1 (sgo__n109), .A2 (n_3258));
NOR2_X1 i_1107 (.ZN (n_2037), .A1 (sgo__n109), .A2 (sgo__n174));
NOR2_X1 i_1106 (.ZN (n_2036), .A1 (sgo__n109), .A2 (sgo__n201));
NOR2_X1 i_1105 (.ZN (n_2035), .A1 (sgo__n109), .A2 (sgo__n147));
NOR2_X1 i_1104 (.ZN (n_2034), .A1 (sgo__n109), .A2 (sgo__n176));
NOR2_X1 i_1103 (.ZN (n_2033), .A1 (sgo__n109), .A2 (n_3263));
NOR2_X1 i_1102 (.ZN (n_2032), .A1 (sgo__n109), .A2 (n_3264));
NOR2_X1 i_1101 (.ZN (n_2031), .A1 (sgo__n109), .A2 (n_3265));
NOR2_X1 i_1100 (.ZN (n_2030), .A1 (sgo__n109), .A2 (n_3266));
NOR2_X1 i_1099 (.ZN (n_2029), .A1 (sgo__n109), .A2 (n_3267));
NOR2_X1 i_1098 (.ZN (n_2028), .A1 (n_3304), .A2 (n_3268));
NOR2_X1 i_1097 (.ZN (n_2027), .A1 (n_3304), .A2 (n_3269));
NOR2_X1 i_1096 (.ZN (n_2026), .A1 (n_3304), .A2 (n_3270));
NOR2_X1 i_1095 (.ZN (n_2025), .A1 (n_3304), .A2 (n_3271));
NOR2_X1 i_1094 (.ZN (n_2024), .A1 (n_3304), .A2 (n_3272));
NOR2_X1 i_1093 (.ZN (n_2023), .A1 (n_3304), .A2 (n_3273));
NOR2_X1 i_1092 (.ZN (n_2022), .A1 (n_3304), .A2 (n_3274));
NOR2_X1 i_1091 (.ZN (n_2021), .A1 (n_3304), .A2 (n_3275));
NOR2_X1 i_1090 (.ZN (n_2020), .A1 (n_3304), .A2 (n_3276));
NOR2_X1 i_1089 (.ZN (n_2019), .A1 (n_3304), .A2 (n_3277));
NOR2_X1 i_1088 (.ZN (n_2018), .A1 (n_3305), .A2 (n_3246));
NOR2_X1 i_1087 (.ZN (n_2017), .A1 (n_3305), .A2 (n_3247));
NOR2_X1 i_1086 (.ZN (n_2016), .A1 (n_3305), .A2 (n_3248));
NOR2_X1 i_1085 (.ZN (n_2015), .A1 (n_3305), .A2 (n_3249));
NOR2_X1 i_1084 (.ZN (n_2014), .A1 (n_3305), .A2 (n_3250));
NOR2_X1 i_1083 (.ZN (n_2013), .A1 (n_3305), .A2 (n_3251));
NOR2_X1 i_1082 (.ZN (n_2012), .A1 (n_3305), .A2 (n_3252));
NOR2_X1 i_1081 (.ZN (n_2011), .A1 (n_3305), .A2 (n_3253));
NOR2_X1 i_1080 (.ZN (n_2010), .A1 (n_3305), .A2 (n_3254));
NOR2_X1 i_1079 (.ZN (n_2009), .A1 (n_3305), .A2 (n_3255));
NOR2_X1 i_1078 (.ZN (n_2008), .A1 (n_3305), .A2 (sgo__n182));
NOR2_X1 i_1077 (.ZN (n_2007), .A1 (n_3305), .A2 (n_3257));
NOR2_X1 i_1076 (.ZN (n_2006), .A1 (n_3305), .A2 (n_3258));
NOR2_X1 i_1075 (.ZN (n_2005), .A1 (n_3305), .A2 (sgo__n174));
NOR2_X1 i_1074 (.ZN (n_2004), .A1 (n_3305), .A2 (sgo__n201));
NOR2_X1 i_1073 (.ZN (n_2003), .A1 (n_3305), .A2 (sgo__n147));
NOR2_X1 i_1072 (.ZN (n_2002), .A1 (n_3305), .A2 (sgo__n176));
NOR2_X1 i_1071 (.ZN (n_2001), .A1 (n_3305), .A2 (n_3263));
NOR2_X1 i_1070 (.ZN (n_2000), .A1 (n_3305), .A2 (n_3264));
NOR2_X1 i_1069 (.ZN (n_1999), .A1 (n_3305), .A2 (n_3265));
NOR2_X1 i_1068 (.ZN (n_1998), .A1 (n_3305), .A2 (n_3266));
NOR2_X1 i_1067 (.ZN (n_1997), .A1 (n_3305), .A2 (n_3267));
NOR2_X1 i_1066 (.ZN (n_1996), .A1 (n_3305), .A2 (n_3268));
NOR2_X1 i_1065 (.ZN (n_1995), .A1 (n_3305), .A2 (n_3269));
NOR2_X1 i_1064 (.ZN (n_1994), .A1 (n_3305), .A2 (n_3270));
NOR2_X1 i_1063 (.ZN (n_1993), .A1 (n_3305), .A2 (n_3271));
NOR2_X1 i_1062 (.ZN (n_1992), .A1 (n_3305), .A2 (n_3272));
NOR2_X1 i_1061 (.ZN (n_1991), .A1 (n_3305), .A2 (n_3273));
NOR2_X1 i_1060 (.ZN (n_1990), .A1 (n_3305), .A2 (n_3274));
NOR2_X1 i_1059 (.ZN (n_1989), .A1 (n_3305), .A2 (n_3275));
NOR2_X1 i_1058 (.ZN (n_1988), .A1 (n_3305), .A2 (n_3276));
NOR2_X1 i_1057 (.ZN (n_1987), .A1 (n_3305), .A2 (n_3277));
NOR2_X1 i_1056 (.ZN (n_1986), .A1 (n_3306), .A2 (n_3246));
NOR2_X1 i_1055 (.ZN (n_1985), .A1 (n_3306), .A2 (n_3247));
NOR2_X1 i_1054 (.ZN (n_1984), .A1 (n_3306), .A2 (n_3248));
NOR2_X1 i_1053 (.ZN (n_1983), .A1 (n_3306), .A2 (n_3249));
NOR2_X1 i_1052 (.ZN (n_1982), .A1 (n_3306), .A2 (n_3250));
NOR2_X1 i_1051 (.ZN (n_1981), .A1 (CLOCK_sgo__n359), .A2 (n_3251));
NOR2_X1 i_1050 (.ZN (n_1980), .A1 (CLOCK_sgo__n359), .A2 (n_3252));
NOR2_X1 i_1049 (.ZN (n_1979), .A1 (CLOCK_sgo__n359), .A2 (n_3253));
NOR2_X1 i_1048 (.ZN (n_1978), .A1 (CLOCK_sgo__n359), .A2 (n_3254));
NOR2_X1 i_1047 (.ZN (n_1977), .A1 (CLOCK_sgo__n359), .A2 (n_3255));
NOR2_X1 i_1046 (.ZN (n_1976), .A1 (CLOCK_sgo__n359), .A2 (sgo__n182));
NOR2_X1 i_1045 (.ZN (n_1975), .A1 (CLOCK_sgo__n359), .A2 (n_3257));
NOR2_X1 i_1044 (.ZN (n_1974), .A1 (CLOCK_sgo__n359), .A2 (n_3258));
NOR2_X1 i_1043 (.ZN (n_1973), .A1 (CLOCK_sgo__n359), .A2 (sgo__n174));
NOR2_X1 i_1042 (.ZN (n_1972), .A1 (CLOCK_sgo__n359), .A2 (sgo__n201));
NOR2_X1 i_1041 (.ZN (n_1971), .A1 (CLOCK_sgo__n359), .A2 (sgo__n147));
NOR2_X1 i_1040 (.ZN (n_1970), .A1 (CLOCK_sgo__n359), .A2 (n_3262));
NOR2_X1 i_1039 (.ZN (n_1969), .A1 (CLOCK_sgo__n359), .A2 (n_3263));
NOR2_X1 i_1038 (.ZN (n_1968), .A1 (n_3306), .A2 (n_3264));
NOR2_X1 i_1037 (.ZN (n_1967), .A1 (n_3306), .A2 (n_3265));
NOR2_X1 i_1036 (.ZN (n_1966), .A1 (n_3306), .A2 (n_3266));
NOR2_X1 i_1035 (.ZN (n_1965), .A1 (n_3306), .A2 (n_3267));
NOR2_X1 i_1034 (.ZN (n_1964), .A1 (CLOCK_sgo__n358), .A2 (n_3268));
NOR2_X1 i_1033 (.ZN (n_1963), .A1 (CLOCK_sgo__n358), .A2 (n_3269));
NOR2_X1 i_1032 (.ZN (n_1962), .A1 (CLOCK_sgo__n358), .A2 (n_3270));
NOR2_X1 i_1031 (.ZN (n_1961), .A1 (CLOCK_sgo__n358), .A2 (n_3271));
NOR2_X1 i_1030 (.ZN (n_1960), .A1 (CLOCK_sgo__n358), .A2 (n_3272));
NOR2_X1 i_1029 (.ZN (n_1959), .A1 (CLOCK_sgo__n358), .A2 (n_3273));
NOR2_X1 i_1028 (.ZN (n_1958), .A1 (CLOCK_sgo__n358), .A2 (n_3274));
NOR2_X1 i_1027 (.ZN (n_1957), .A1 (CLOCK_sgo__n358), .A2 (n_3275));
NOR2_X1 i_1026 (.ZN (n_1956), .A1 (n_3306), .A2 (n_3276));
NOR2_X1 i_1025 (.ZN (n_1955), .A1 (n_3306), .A2 (n_3277));
NOR2_X1 i_1024 (.ZN (n_1954), .A1 (n_3307), .A2 (n_3246));
NOR2_X1 i_1023 (.ZN (n_1953), .A1 (n_3307), .A2 (n_3247));
NOR2_X1 i_1022 (.ZN (n_1952), .A1 (n_3307), .A2 (n_3248));
NOR2_X1 i_1021 (.ZN (n_1951), .A1 (n_3307), .A2 (n_3249));
NOR2_X1 i_1020 (.ZN (n_1950), .A1 (n_3307), .A2 (n_3250));
NOR2_X1 i_1019 (.ZN (n_1949), .A1 (n_3307), .A2 (n_3251));
NOR2_X1 i_1018 (.ZN (n_1948), .A1 (n_3307), .A2 (n_3252));
NOR2_X1 i_1017 (.ZN (n_1947), .A1 (n_3307), .A2 (n_3253));
NOR2_X1 i_1016 (.ZN (n_1946), .A1 (n_3307), .A2 (n_3254));
NOR2_X1 i_1015 (.ZN (n_1945), .A1 (n_3307), .A2 (n_3255));
NOR2_X1 i_1014 (.ZN (n_1944), .A1 (n_3307), .A2 (sgo__n182));
NOR2_X1 i_1013 (.ZN (n_1943), .A1 (n_3307), .A2 (n_3257));
NOR2_X1 i_1012 (.ZN (n_1942), .A1 (n_3307), .A2 (n_3258));
NOR2_X1 i_1011 (.ZN (n_1941), .A1 (n_3307), .A2 (sgo__n174));
NOR2_X1 i_1010 (.ZN (n_1940), .A1 (n_3307), .A2 (n_3260));
NOR2_X1 i_1009 (.ZN (n_1939), .A1 (n_3307), .A2 (sgo__n147));
NOR2_X1 i_1008 (.ZN (n_1938), .A1 (n_3307), .A2 (sgo__n176));
NOR2_X1 i_1007 (.ZN (n_1937), .A1 (n_3307), .A2 (n_3263));
NOR2_X1 i_1006 (.ZN (n_1936), .A1 (n_3307), .A2 (n_3264));
NOR2_X1 i_1005 (.ZN (n_1935), .A1 (n_3307), .A2 (n_3265));
NOR2_X1 i_1004 (.ZN (n_1934), .A1 (n_3307), .A2 (n_3266));
NOR2_X1 i_1003 (.ZN (n_1933), .A1 (n_3307), .A2 (n_3267));
NOR2_X1 i_1002 (.ZN (n_1932), .A1 (n_3307), .A2 (n_3268));
NOR2_X1 i_1001 (.ZN (n_1931), .A1 (n_3307), .A2 (n_3269));
NOR2_X1 i_1000 (.ZN (n_1930), .A1 (n_3307), .A2 (n_3270));
NOR2_X1 i_999 (.ZN (n_1929), .A1 (n_3307), .A2 (n_3271));
NOR2_X1 i_998 (.ZN (n_1928), .A1 (n_3307), .A2 (n_3272));
NOR2_X1 i_997 (.ZN (n_1927), .A1 (n_3307), .A2 (n_3273));
NOR2_X1 i_996 (.ZN (n_1926), .A1 (n_3307), .A2 (n_3274));
NOR2_X1 i_995 (.ZN (n_1925), .A1 (n_3307), .A2 (n_3275));
NOR2_X1 i_994 (.ZN (n_1924), .A1 (n_3307), .A2 (n_3276));
NOR2_X1 i_993 (.ZN (n_1923), .A1 (n_3307), .A2 (n_3277));
NOR2_X1 i_992 (.ZN (n_1922), .A1 (n_3308), .A2 (n_3246));
NOR2_X1 i_991 (.ZN (n_1921), .A1 (n_3308), .A2 (n_3247));
NOR2_X1 i_990 (.ZN (n_1920), .A1 (n_3308), .A2 (n_3248));
NOR2_X1 i_989 (.ZN (n_1919), .A1 (n_3308), .A2 (sgo__n10));
NOR2_X1 i_988 (.ZN (n_1918), .A1 (n_3308), .A2 (n_3250));
NOR2_X1 i_987 (.ZN (n_1917), .A1 (n_3308), .A2 (n_3251));
NOR2_X1 i_986 (.ZN (n_1916), .A1 (n_3308), .A2 (n_3252));
NOR2_X1 i_985 (.ZN (n_1915), .A1 (n_3308), .A2 (n_3253));
NOR2_X1 i_984 (.ZN (n_1914), .A1 (n_3308), .A2 (n_3254));
NOR2_X1 i_983 (.ZN (n_1913), .A1 (n_3308), .A2 (n_3255));
NOR2_X1 i_982 (.ZN (n_1912), .A1 (n_3308), .A2 (sgo__n182));
NOR2_X1 i_981 (.ZN (n_1911), .A1 (n_3308), .A2 (n_3257));
NOR2_X1 i_980 (.ZN (n_1910), .A1 (n_3308), .A2 (n_3258));
NOR2_X1 i_979 (.ZN (n_1909), .A1 (n_3308), .A2 (sgo__n174));
NOR2_X1 i_978 (.ZN (n_1908), .A1 (n_3308), .A2 (n_3260));
NOR2_X1 i_977 (.ZN (n_1907), .A1 (n_3308), .A2 (sgo__n147));
NOR2_X1 i_976 (.ZN (n_1906), .A1 (n_3308), .A2 (sgo__n176));
NOR2_X1 i_975 (.ZN (n_1905), .A1 (n_3308), .A2 (n_3263));
NOR2_X1 i_974 (.ZN (n_1904), .A1 (n_3308), .A2 (n_3264));
NOR2_X1 i_973 (.ZN (n_1903), .A1 (n_3308), .A2 (n_3265));
NOR2_X1 i_972 (.ZN (n_1902), .A1 (n_3308), .A2 (n_3266));
NOR2_X1 i_971 (.ZN (n_1901), .A1 (n_3308), .A2 (n_3267));
NOR2_X1 i_970 (.ZN (n_1900), .A1 (n_3308), .A2 (n_3268));
NOR2_X1 i_969 (.ZN (n_1899), .A1 (n_3308), .A2 (n_3269));
NOR2_X1 i_968 (.ZN (n_1898), .A1 (n_3308), .A2 (n_3270));
NOR2_X1 i_967 (.ZN (n_1897), .A1 (n_3308), .A2 (n_3271));
NOR2_X1 i_966 (.ZN (n_1896), .A1 (n_3308), .A2 (n_3272));
NOR2_X1 i_965 (.ZN (n_1895), .A1 (n_3308), .A2 (n_3273));
NOR2_X1 i_964 (.ZN (n_1894), .A1 (n_3308), .A2 (n_3274));
NOR2_X1 i_963 (.ZN (n_1893), .A1 (n_3308), .A2 (n_3275));
NOR2_X1 i_962 (.ZN (n_1892), .A1 (n_3308), .A2 (n_3276));
NOR2_X1 i_961 (.ZN (n_1891), .A1 (n_3308), .A2 (n_3277));
NOR2_X2 i_960 (.ZN (n_1890), .A1 (n_3309), .A2 (n_3246));
NOR2_X1 i_959 (.ZN (n_1889), .A1 (n_3309), .A2 (n_3247));
NOR2_X1 i_958 (.ZN (n_1888), .A1 (n_3309), .A2 (n_3248));
NOR2_X1 i_957 (.ZN (n_1887), .A1 (n_3309), .A2 (sgo__n10));
NOR2_X1 i_956 (.ZN (n_1886), .A1 (n_3309), .A2 (n_3250));
NOR2_X1 i_955 (.ZN (n_1885), .A1 (n_3309), .A2 (n_3251));
NOR2_X1 i_954 (.ZN (n_1884), .A1 (n_3309), .A2 (n_3252));
NOR2_X1 i_953 (.ZN (n_1883), .A1 (n_3309), .A2 (n_3253));
NOR2_X1 i_952 (.ZN (n_1882), .A1 (n_3309), .A2 (n_3254));
NOR2_X1 i_951 (.ZN (n_1881), .A1 (n_3309), .A2 (n_3255));
NOR2_X1 i_950 (.ZN (n_1880), .A1 (n_3309), .A2 (sgo__n182));
NOR2_X1 i_949 (.ZN (n_1879), .A1 (n_3309), .A2 (n_3257));
NOR2_X1 i_948 (.ZN (n_1878), .A1 (n_3309), .A2 (n_3258));
NOR2_X1 i_947 (.ZN (n_1877), .A1 (n_3309), .A2 (n_3259));
NOR2_X1 i_946 (.ZN (n_1876), .A1 (n_3309), .A2 (n_3260));
NOR2_X1 i_945 (.ZN (n_1875), .A1 (n_3309), .A2 (sgo__n147));
NOR2_X1 i_944 (.ZN (n_1874), .A1 (n_3309), .A2 (n_3262));
NOR2_X1 i_943 (.ZN (n_1873), .A1 (n_3309), .A2 (n_3263));
NOR2_X1 i_942 (.ZN (n_1872), .A1 (n_3309), .A2 (n_3264));
NOR2_X1 i_941 (.ZN (n_1871), .A1 (n_3309), .A2 (n_3265));
NOR2_X1 i_940 (.ZN (n_1870), .A1 (n_3309), .A2 (n_3266));
NOR2_X1 i_939 (.ZN (n_1869), .A1 (n_3309), .A2 (n_3267));
NOR2_X1 i_938 (.ZN (n_1868), .A1 (n_3309), .A2 (n_3268));
NOR2_X1 i_937 (.ZN (n_1867), .A1 (n_3309), .A2 (n_3269));
NOR2_X1 i_936 (.ZN (n_1866), .A1 (n_3309), .A2 (n_3270));
NOR2_X1 i_935 (.ZN (n_1865), .A1 (n_3309), .A2 (n_3271));
NOR2_X1 i_934 (.ZN (n_1864), .A1 (n_3309), .A2 (n_3272));
NOR2_X1 i_933 (.ZN (n_1863), .A1 (n_3309), .A2 (n_3273));
NOR2_X1 i_932 (.ZN (n_1862), .A1 (n_3309), .A2 (n_3274));
NOR2_X1 i_931 (.ZN (n_1861), .A1 (n_3309), .A2 (n_3275));
NOR2_X1 i_930 (.ZN (n_1860), .A1 (n_3309), .A2 (n_3276));
FA_X1 i_929 (.CO (n_1859), .S (n_1858), .A (n_1860), .B (n_1891), .CI (n_1855));
FA_X1 i_928 (.CO (n_1857), .S (n_1856), .A (n_1849), .B (n_1854), .CI (n_1851));
FA_X1 i_927 (.CO (n_1855), .S (n_1854), .A (n_1861), .B (n_1892), .CI (n_1923));
FA_X1 i_926 (.CO (n_1853), .S (n_1852), .A (n_1848), .B (n_1850), .CI (n_1845));
FA_X1 i_925 (.CO (n_1851), .S (n_1850), .A (n_1955), .B (n_1841), .CI (n_1843));
FA_X1 i_924 (.CO (n_1849), .S (n_1848), .A (n_1862), .B (n_1893), .CI (n_1924));
FA_X1 i_923 (.CO (n_1847), .S (n_1846), .A (n_1835), .B (n_1837), .CI (n_1844));
FA_X1 i_922 (.CO (n_1845), .S (n_1844), .A (n_1831), .B (n_1842), .CI (n_1840));
FA_X1 i_921 (.CO (n_1843), .S (n_1842), .A (n_1956), .B (n_1987), .CI (n_1833));
FA_X1 i_920 (.CO (n_1841), .S (n_1840), .A (n_1863), .B (n_1894), .CI (n_1925));
FA_X1 i_919 (.CO (n_1839), .S (n_1838), .A (n_1825), .B (n_1827), .CI (n_1836));
FA_X1 i_918 (.CO (n_1837), .S (n_1836), .A (n_1832), .B (n_1830), .CI (n_1834));
FA_X1 i_917 (.CO (n_1835), .S (n_1834), .A (n_1821), .B (n_1819), .CI (n_1823));
FA_X1 i_916 (.CO (n_1833), .S (n_1832), .A (n_1957), .B (n_1988), .CI (n_2019));
FA_X1 i_915 (.CO (n_1831), .S (n_1830), .A (n_1864), .B (n_1895), .CI (n_1926));
FA_X1 i_914 (.CO (n_1829), .S (n_1828), .A (n_1824), .B (n_1815), .CI (n_1826));
FA_X1 i_913 (.CO (n_1827), .S (n_1826), .A (n_1811), .B (n_1822), .CI (n_1813));
FA_X1 i_912 (.CO (n_1825), .S (n_1824), .A (n_1809), .B (n_1820), .CI (n_1818));
FA_X1 i_911 (.CO (n_1823), .S (n_1822), .A (n_2051), .B (n_1807), .CI (n_1805));
FA_X1 i_910 (.CO (n_1821), .S (n_1820), .A (n_1958), .B (n_1989), .CI (n_2020));
FA_X1 i_909 (.CO (n_1819), .S (n_1818), .A (n_1865), .B (n_1896), .CI (n_1927));
FA_X1 i_908 (.CO (n_1817), .S (n_1816), .A (n_1812), .B (n_1814), .CI (n_1801));
FA_X1 i_907 (.CO (n_1815), .S (n_1814), .A (n_1810), .B (n_1797), .CI (n_1799));
FA_X1 i_906 (.CO (n_1813), .S (n_1812), .A (n_1808), .B (n_1806), .CI (n_1804));
FA_X1 i_905 (.CO (n_1811), .S (n_1810), .A (n_1791), .B (n_1789), .CI (n_1795));
FA_X1 i_904 (.CO (n_1809), .S (n_1808), .A (n_2052), .B (n_2083), .CI (n_1793));
FA_X1 i_903 (.CO (n_1807), .S (n_1806), .A (n_1959), .B (n_1990), .CI (n_2021));
FA_X1 i_902 (.CO (n_1805), .S (n_1804), .A (n_1866), .B (n_1897), .CI (n_1928));
FA_X1 i_901 (.CO (n_1803), .S (n_1802), .A (n_1783), .B (n_1785), .CI (n_1800));
FA_X1 i_900 (.CO (n_1801), .S (n_1800), .A (n_1781), .B (n_1796), .CI (n_1798));
FA_X1 i_899 (.CO (n_1799), .S (n_1798), .A (n_1788), .B (n_1779), .CI (n_1794));
FA_X1 i_898 (.CO (n_1797), .S (n_1796), .A (n_1777), .B (n_1792), .CI (n_1790));
FA_X1 i_897 (.CO (n_1795), .S (n_1794), .A (n_1775), .B (n_1773), .CI (n_1771));
FA_X1 i_896 (.CO (n_1793), .S (n_1792), .A (n_2053), .B (n_2084), .CI (n_2115));
FA_X1 i_895 (.CO (n_1791), .S (n_1790), .A (n_1960), .B (n_1991), .CI (n_2022));
FA_X1 i_894 (.CO (n_1789), .S (n_1788), .A (n_1867), .B (n_1898), .CI (n_1929));
FA_X1 i_893 (.CO (n_1787), .S (n_1786), .A (n_1782), .B (n_1767), .CI (n_1784));
FA_X1 i_892 (.CO (n_1785), .S (n_1784), .A (n_1763), .B (n_1780), .CI (n_1765));
FA_X1 i_891 (.CO (n_1783), .S (n_1782), .A (n_1776), .B (n_1761), .CI (n_1778));
FA_X1 i_890 (.CO (n_1781), .S (n_1780), .A (n_1774), .B (n_1772), .CI (n_1770));
FA_X1 i_889 (.CO (n_1779), .S (n_1778), .A (n_1751), .B (n_1759), .CI (n_1757));
FA_X1 i_888 (.CO (n_1777), .S (n_1776), .A (n_2147), .B (n_1755), .CI (n_1753));
FA_X1 i_887 (.CO (n_1775), .S (n_1774), .A (n_2054), .B (n_2085), .CI (n_2116));
FA_X1 i_886 (.CO (n_1773), .S (n_1772), .A (n_1961), .B (n_1992), .CI (n_2023));
FA_X1 i_885 (.CO (n_1771), .S (n_1770), .A (n_1868), .B (n_1899), .CI (n_1930));
FA_X1 i_884 (.CO (n_1769), .S (n_1768), .A (n_1764), .B (n_1747), .CI (n_1766));
FA_X1 i_883 (.CO (n_1767), .S (n_1766), .A (n_1762), .B (n_1760), .CI (n_1745));
FA_X1 i_882 (.CO (n_1765), .S (n_1764), .A (n_1741), .B (n_1739), .CI (n_1743));
FA_X1 i_881 (.CO (n_1763), .S (n_1762), .A (n_1752), .B (n_1750), .CI (n_1758));
FA_X1 i_880 (.CO (n_1761), .S (n_1760), .A (n_1737), .B (n_1756), .CI (n_1754));
FA_X1 i_879 (.CO (n_1759), .S (n_1758), .A (n_1733), .B (n_1731), .CI (n_1729));
FA_X1 i_878 (.CO (n_1757), .S (n_1756), .A (n_2148), .B (n_2179), .CI (n_1735));
FA_X1 i_877 (.CO (n_1755), .S (n_1754), .A (n_2055), .B (n_2086), .CI (n_2117));
FA_X1 i_876 (.CO (n_1753), .S (n_1752), .A (n_1962), .B (n_1993), .CI (n_2024));
FA_X1 i_875 (.CO (n_1751), .S (n_1750), .A (n_1869), .B (n_1900), .CI (n_1931));
FA_X1 i_874 (.CO (n_1749), .S (n_1748), .A (n_1744), .B (n_1725), .CI (n_1746));
FA_X1 i_873 (.CO (n_1747), .S (n_1746), .A (n_1740), .B (n_1742), .CI (n_1723));
FA_X1 i_872 (.CO (n_1745), .S (n_1744), .A (n_1738), .B (n_1721), .CI (n_1719));
FA_X1 i_871 (.CO (n_1743), .S (n_1742), .A (n_1715), .B (n_1736), .CI (n_1717));
FA_X1 i_870 (.CO (n_1741), .S (n_1740), .A (n_1732), .B (n_1730), .CI (n_1728));
FA_X1 i_869 (.CO (n_1739), .S (n_1738), .A (n_1705), .B (n_1713), .CI (n_1734));
FA_X1 i_868 (.CO (n_1737), .S (n_1736), .A (n_1711), .B (n_1709), .CI (n_1707));
FA_X1 i_867 (.CO (n_1735), .S (n_1734), .A (n_2149), .B (n_2180), .CI (n_2211));
FA_X1 i_866 (.CO (n_1733), .S (n_1732), .A (n_2056), .B (n_2087), .CI (n_2118));
FA_X1 i_865 (.CO (n_1731), .S (n_1730), .A (n_1963), .B (n_1994), .CI (n_2025));
FA_X1 i_864 (.CO (n_1729), .S (n_1728), .A (n_1870), .B (n_1901), .CI (n_1932));
FA_X1 i_863 (.CO (n_1727), .S (n_1726), .A (n_1701), .B (n_1722), .CI (n_1724));
FA_X1 i_862 (.CO (n_1725), .S (n_1724), .A (n_1697), .B (n_1720), .CI (n_1699));
FA_X1 i_861 (.CO (n_1723), .S (n_1722), .A (n_1695), .B (n_1718), .CI (n_1716));
FA_X1 i_860 (.CO (n_1721), .S (n_1720), .A (n_1712), .B (n_1693), .CI (n_1691));
FA_X1 i_859 (.CO (n_1719), .S (n_1718), .A (n_1706), .B (n_1704), .CI (n_1714));
FA_X1 i_858 (.CO (n_1717), .S (n_1716), .A (n_1687), .B (n_1710), .CI (n_1708));
FA_X1 i_857 (.CO (n_1715), .S (n_1714), .A (n_1681), .B (n_1679), .CI (n_1689));
FA_X1 i_856 (.CO (n_1713), .S (n_1712), .A (n_2243), .B (n_1685), .CI (n_1683));
FA_X1 i_855 (.CO (n_1711), .S (n_1710), .A (n_2150), .B (n_2181), .CI (n_2212));
FA_X1 i_854 (.CO (n_1709), .S (n_1708), .A (n_2057), .B (n_2088), .CI (n_2119));
FA_X1 i_853 (.CO (n_1707), .S (n_1706), .A (n_1964), .B (n_1995), .CI (n_2026));
FA_X1 i_852 (.CO (n_1705), .S (n_1704), .A (n_1871), .B (n_1902), .CI (n_1933));
FA_X1 i_851 (.CO (n_1703), .S (n_1702), .A (n_1698), .B (n_1675), .CI (n_1700));
FA_X1 i_850 (.CO (n_1701), .S (n_1700), .A (n_1671), .B (n_1696), .CI (n_1673));
FA_X1 i_849 (.CO (n_1699), .S (n_1698), .A (n_1669), .B (n_1692), .CI (n_1694));
FA_X1 i_848 (.CO (n_1697), .S (n_1696), .A (n_1667), .B (n_1665), .CI (n_1690));
FA_X1 i_847 (.CO (n_1695), .S (n_1694), .A (n_1678), .B (n_1663), .CI (n_1688));
FA_X1 i_846 (.CO (n_1693), .S (n_1692), .A (n_1684), .B (n_1682), .CI (n_1680));
FA_X1 i_845 (.CO (n_1691), .S (n_1690), .A (n_1651), .B (n_1661), .CI (n_1686));
FA_X1 i_844 (.CO (n_1689), .S (n_1688), .A (n_1657), .B (n_1655), .CI (n_1653));
FA_X1 i_843 (.CO (n_1687), .S (n_1686), .A (n_2244), .B (n_2275), .CI (n_1659));
FA_X1 i_842 (.CO (n_1685), .S (n_1684), .A (n_2151), .B (n_2182), .CI (n_2213));
FA_X1 i_841 (.CO (n_1683), .S (n_1682), .A (n_2058), .B (n_2089), .CI (n_2120));
FA_X1 i_840 (.CO (n_1681), .S (n_1680), .A (n_1965), .B (n_1996), .CI (n_2027));
FA_X1 i_839 (.CO (n_1679), .S (n_1678), .A (n_1872), .B (n_1903), .CI (n_1934));
FA_X1 i_838 (.CO (n_1677), .S (n_1676), .A (n_1672), .B (n_1647), .CI (n_1674));
FA_X1 i_837 (.CO (n_1675), .S (n_1674), .A (n_1668), .B (n_1670), .CI (n_1645));
FA_X1 i_836 (.CO (n_1673), .S (n_1672), .A (n_1666), .B (n_1664), .CI (n_1643));
FA_X1 i_835 (.CO (n_1671), .S (n_1670), .A (n_1635), .B (n_1641), .CI (n_1639));
FA_X1 i_834 (.CO (n_1669), .S (n_1668), .A (n_1662), .B (n_1660), .CI (n_1637));
FA_X1 i_833 (.CO (n_1667), .S (n_1666), .A (n_1654), .B (n_1652), .CI (n_1650));
FA_X1 i_832 (.CO (n_1665), .S (n_1664), .A (n_1631), .B (n_1658), .CI (n_1656));
FA_X1 i_831 (.CO (n_1663), .S (n_1662), .A (n_1623), .B (n_1621), .CI (n_1633));
FA_X1 i_830 (.CO (n_1661), .S (n_1660), .A (n_1629), .B (n_1627), .CI (n_1625));
FA_X1 i_829 (.CO (n_1659), .S (n_1658), .A (n_2245), .B (n_2276), .CI (n_2307));
FA_X1 i_828 (.CO (n_1657), .S (n_1656), .A (n_2152), .B (n_2183), .CI (n_2214));
FA_X1 i_827 (.CO (n_1655), .S (n_1654), .A (n_2059), .B (n_2090), .CI (n_2121));
FA_X1 i_826 (.CO (n_1653), .S (n_1652), .A (n_1966), .B (n_1997), .CI (n_2028));
FA_X1 i_825 (.CO (n_1651), .S (n_1650), .A (n_1873), .B (n_1904), .CI (n_1935));
FA_X1 i_824 (.CO (n_1649), .S (n_1648), .A (n_1644), .B (n_1617), .CI (n_1646));
FA_X1 i_823 (.CO (n_1647), .S (n_1646), .A (n_1613), .B (n_1642), .CI (n_1615));
FA_X1 i_822 (.CO (n_1645), .S (n_1644), .A (n_1636), .B (n_1638), .CI (n_1640));
FA_X1 i_821 (.CO (n_1643), .S (n_1642), .A (n_1634), .B (n_1609), .CI (n_1611));
FA_X1 i_820 (.CO (n_1641), .S (n_1640), .A (n_1630), .B (n_1607), .CI (n_1605));
FA_X1 i_819 (.CO (n_1639), .S (n_1638), .A (n_1620), .B (n_1603), .CI (n_1632));
FA_X1 i_818 (.CO (n_1637), .S (n_1636), .A (n_1626), .B (n_1624), .CI (n_1622));
FA_X1 i_817 (.CO (n_1635), .S (n_1634), .A (n_1601), .B (n_1599), .CI (n_1628));
FA_X1 i_816 (.CO (n_1633), .S (n_1632), .A (n_1593), .B (n_1591), .CI (n_1589));
FA_X1 i_815 (.CO (n_1631), .S (n_1630), .A (n_2339), .B (n_1597), .CI (n_1595));
FA_X1 i_814 (.CO (n_1629), .S (n_1628), .A (n_2246), .B (n_2277), .CI (n_2308));
FA_X1 i_813 (.CO (n_1627), .S (n_1626), .A (n_2153), .B (n_2184), .CI (n_2215));
FA_X1 i_812 (.CO (n_1625), .S (n_1624), .A (n_2060), .B (n_2091), .CI (n_2122));
FA_X1 i_811 (.CO (n_1623), .S (n_1622), .A (n_1967), .B (n_1998), .CI (n_2029));
FA_X1 i_810 (.CO (n_1621), .S (n_1620), .A (n_1874), .B (n_1905), .CI (n_1936));
FA_X1 i_809 (.CO (n_1619), .S (n_1618), .A (n_1614), .B (n_1585), .CI (n_1616));
FA_X1 i_808 (.CO (n_1617), .S (n_1616), .A (n_1581), .B (n_1612), .CI (n_1583));
FA_X1 i_807 (.CO (n_1615), .S (n_1614), .A (n_1579), .B (n_1610), .CI (n_1608));
FA_X1 i_806 (.CO (n_1613), .S (n_1612), .A (n_1577), .B (n_1606), .CI (n_1604));
FA_X1 i_805 (.CO (n_1611), .S (n_1610), .A (n_1573), .B (n_1571), .CI (n_1575));
FA_X1 i_804 (.CO (n_1609), .S (n_1608), .A (n_1588), .B (n_1602), .CI (n_1600));
FA_X1 i_803 (.CO (n_1607), .S (n_1606), .A (n_1594), .B (n_1592), .CI (n_1590));
FA_X1 i_802 (.CO (n_1605), .S (n_1604), .A (n_1567), .B (n_1598), .CI (n_1596));
FA_X1 i_801 (.CO (n_1603), .S (n_1602), .A (n_1557), .B (n_1555), .CI (n_1569));
FA_X1 i_800 (.CO (n_1601), .S (n_1600), .A (n_1563), .B (n_1561), .CI (n_1559));
FA_X1 i_799 (.CO (n_1599), .S (n_1598), .A (n_2340), .B (n_2371), .CI (n_1565));
FA_X1 i_798 (.CO (n_1597), .S (n_1596), .A (n_2247), .B (n_2278), .CI (n_2309));
FA_X1 i_797 (.CO (n_1595), .S (n_1594), .A (n_2154), .B (n_2185), .CI (n_2216));
FA_X1 i_796 (.CO (n_1593), .S (n_1592), .A (n_2061), .B (n_2092), .CI (n_2123));
FA_X1 i_795 (.CO (n_1591), .S (n_1590), .A (n_1968), .B (n_1999), .CI (n_2030));
FA_X1 i_794 (.CO (n_1589), .S (n_1588), .A (n_1875), .B (n_1906), .CI (n_1937));
FA_X1 i_793 (.CO (n_1587), .S (n_1586), .A (n_1582), .B (n_1551), .CI (n_1584));
FA_X1 i_792 (.CO (n_1585), .S (n_1584), .A (n_1547), .B (n_1580), .CI (n_1549));
FA_X1 i_791 (.CO (n_1583), .S (n_1582), .A (n_1576), .B (n_1545), .CI (n_1578));
FA_X1 i_790 (.CO (n_1581), .S (n_1580), .A (n_1541), .B (n_1574), .CI (n_1572));
FA_X1 i_789 (.CO (n_1579), .S (n_1578), .A (n_1537), .B (n_1570), .CI (n_1543));
FA_X1 i_788 (.CO (n_1577), .S (n_1576), .A (n_1568), .B (n_1566), .CI (n_1539));
FA_X1 i_787 (.CO (n_1575), .S (n_1574), .A (n_1556), .B (n_1554), .CI (n_1535));
FA_X1 i_786 (.CO (n_1573), .S (n_1572), .A (n_1562), .B (n_1560), .CI (n_1558));
FA_X1 i_785 (.CO (n_1571), .S (n_1570), .A (n_1533), .B (n_1531), .CI (n_1564));
FA_X1 i_784 (.CO (n_1569), .S (n_1568), .A (n_1523), .B (n_1521), .CI (n_1519));
FA_X1 i_783 (.CO (n_1567), .S (n_1566), .A (n_1529), .B (n_1527), .CI (n_1525));
FA_X1 i_782 (.CO (n_1565), .S (n_1564), .A (n_2341), .B (n_2372), .CI (n_2403));
FA_X1 i_781 (.CO (n_1563), .S (n_1562), .A (n_2248), .B (n_2279), .CI (n_2310));
FA_X1 i_780 (.CO (n_1561), .S (n_1560), .A (n_2155), .B (n_2186), .CI (n_2217));
FA_X1 i_779 (.CO (n_1559), .S (n_1558), .A (n_2062), .B (n_2093), .CI (n_2124));
FA_X1 i_778 (.CO (n_1557), .S (n_1556), .A (n_1969), .B (n_2000), .CI (n_2031));
FA_X1 i_777 (.CO (n_1555), .S (n_1554), .A (n_1876), .B (n_1907), .CI (n_1938));
FA_X1 i_776 (.CO (n_1553), .S (n_1552), .A (n_1548), .B (n_1515), .CI (n_1550));
FA_X1 i_775 (.CO (n_1551), .S (n_1550), .A (n_1511), .B (n_1546), .CI (n_1513));
FA_X1 i_774 (.CO (n_1549), .S (n_1548), .A (n_1540), .B (n_1509), .CI (n_1544));
FA_X1 i_773 (.CO (n_1547), .S (n_1546), .A (n_1536), .B (n_1507), .CI (n_1542));
FA_X1 i_772 (.CO (n_1545), .S (n_1544), .A (n_1534), .B (n_1505), .CI (n_1538));
FA_X1 i_771 (.CO (n_1543), .S (n_1542), .A (n_1503), .B (n_1501), .CI (n_1499));
FA_X1 i_770 (.CO (n_1541), .S (n_1540), .A (n_1518), .B (n_1532), .CI (n_1530));
FA_X1 i_769 (.CO (n_1539), .S (n_1538), .A (n_1524), .B (n_1522), .CI (n_1520));
FA_X1 i_768 (.CO (n_1537), .S (n_1536), .A (n_1493), .B (n_1528), .CI (n_1526));
FA_X1 i_767 (.CO (n_1535), .S (n_1534), .A (n_1481), .B (n_1497), .CI (n_1495));
FA_X1 i_766 (.CO (n_1533), .S (n_1532), .A (n_1487), .B (n_1485), .CI (n_1483));
FA_X1 i_765 (.CO (n_1531), .S (n_1530), .A (n_2435), .B (n_1491), .CI (n_1489));
FA_X1 i_764 (.CO (n_1529), .S (n_1528), .A (n_2342), .B (n_2373), .CI (n_2404));
FA_X1 i_763 (.CO (n_1527), .S (n_1526), .A (n_2249), .B (n_2280), .CI (n_2311));
FA_X1 i_762 (.CO (n_1525), .S (n_1524), .A (n_2156), .B (n_2187), .CI (n_2218));
FA_X1 i_761 (.CO (n_1523), .S (n_1522), .A (n_2063), .B (n_2094), .CI (n_2125));
FA_X1 i_760 (.CO (n_1521), .S (n_1520), .A (n_1970), .B (n_2001), .CI (n_2032));
FA_X1 i_759 (.CO (n_1519), .S (n_1518), .A (n_1877), .B (n_1908), .CI (n_1939));
FA_X1 i_758 (.CO (n_1517), .S (n_1516), .A (n_1512), .B (n_1477), .CI (n_1514));
FA_X1 i_757 (.CO (n_1515), .S (n_1514), .A (n_1473), .B (n_1510), .CI (n_1475));
FA_X1 i_756 (.CO (n_1513), .S (n_1512), .A (n_1504), .B (n_1471), .CI (n_1508));
FA_X1 i_755 (.CO (n_1511), .S (n_1510), .A (n_1500), .B (n_1469), .CI (n_1506));
FA_X1 i_754 (.CO (n_1509), .S (n_1508), .A (n_1467), .B (n_1465), .CI (n_1502));
FA_X1 i_753 (.CO (n_1507), .S (n_1506), .A (n_1463), .B (n_1461), .CI (n_1498));
FA_X1 i_752 (.CO (n_1505), .S (n_1504), .A (n_1459), .B (n_1496), .CI (n_1494));
FA_X1 i_751 (.CO (n_1503), .S (n_1502), .A (n_1484), .B (n_1482), .CI (n_1480));
FA_X1 i_750 (.CO (n_1501), .S (n_1500), .A (n_1490), .B (n_1488), .CI (n_1486));
FA_X1 i_749 (.CO (n_1499), .S (n_1498), .A (n_1457), .B (n_1455), .CI (n_1492));
FA_X1 i_748 (.CO (n_1497), .S (n_1496), .A (n_1445), .B (n_1443), .CI (n_1441));
FA_X1 i_747 (.CO (n_1495), .S (n_1494), .A (n_1451), .B (n_1449), .CI (n_1447));
FA_X1 i_746 (.CO (n_1493), .S (n_1492), .A (n_2436), .B (n_2467), .CI (n_1453));
FA_X1 i_745 (.CO (n_1491), .S (n_1490), .A (n_2343), .B (n_2374), .CI (n_2405));
FA_X1 i_744 (.CO (n_1489), .S (n_1488), .A (n_2250), .B (n_2281), .CI (n_2312));
FA_X1 i_743 (.CO (n_1487), .S (n_1486), .A (n_2157), .B (n_2188), .CI (n_2219));
FA_X1 i_742 (.CO (n_1485), .S (n_1484), .A (n_2064), .B (n_2095), .CI (n_2126));
FA_X1 i_741 (.CO (n_1483), .S (n_1482), .A (n_1971), .B (n_2002), .CI (n_2033));
FA_X1 i_740 (.CO (n_1481), .S (n_1480), .A (n_1878), .B (n_1909), .CI (n_1940));
FA_X1 i_739 (.CO (n_1479), .S (n_1478), .A (n_1474), .B (n_1437), .CI (n_1476));
FA_X1 i_738 (.CO (n_1477), .S (n_1476), .A (n_1470), .B (n_1472), .CI (n_1435));
FA_X1 i_737 (.CO (n_1475), .S (n_1474), .A (n_1431), .B (n_1468), .CI (n_1433));
FA_X1 i_736 (.CO (n_1473), .S (n_1472), .A (n_1464), .B (n_1429), .CI (n_1466));
FA_X1 i_735 (.CO (n_1471), .S (n_1470), .A (n_1425), .B (n_1462), .CI (n_1460));
FA_X1 i_734 (.CO (n_1469), .S (n_1468), .A (n_1419), .B (n_1458), .CI (n_1427));
FA_X1 i_733 (.CO (n_1467), .S (n_1466), .A (n_1454), .B (n_1423), .CI (n_1421));
FA_X1 i_732 (.CO (n_1465), .S (n_1464), .A (n_1440), .B (n_1417), .CI (n_1456));
FA_X1 i_731 (.CO (n_1463), .S (n_1462), .A (n_1446), .B (n_1444), .CI (n_1442));
FA_X1 i_730 (.CO (n_1461), .S (n_1460), .A (n_1452), .B (n_1450), .CI (n_1448));
FA_X1 i_729 (.CO (n_1459), .S (n_1458), .A (n_1399), .B (n_1415), .CI (n_1413));
FA_X1 i_728 (.CO (n_1457), .S (n_1456), .A (n_1405), .B (n_1403), .CI (n_1401));
FA_X1 i_727 (.CO (n_1455), .S (n_1454), .A (n_1411), .B (n_1409), .CI (n_1407));
FA_X1 i_726 (.CO (n_1453), .S (n_1452), .A (n_2437), .B (n_2468), .CI (n_2499));
FA_X1 i_725 (.CO (n_1451), .S (n_1450), .A (n_2344), .B (n_2375), .CI (n_2406));
FA_X1 i_724 (.CO (n_1449), .S (n_1448), .A (n_2251), .B (n_2282), .CI (n_2313));
FA_X1 i_723 (.CO (n_1447), .S (n_1446), .A (n_2158), .B (n_2189), .CI (n_2220));
FA_X1 i_722 (.CO (n_1445), .S (n_1444), .A (n_2065), .B (n_2096), .CI (n_2127));
FA_X1 i_721 (.CO (n_1443), .S (n_1442), .A (n_1972), .B (n_2003), .CI (n_2034));
FA_X1 i_720 (.CO (n_1441), .S (n_1440), .A (n_1879), .B (n_1910), .CI (n_1941));
FA_X1 i_719 (.CO (n_1439), .S (n_1438), .A (n_1434), .B (n_1395), .CI (n_1436));
FA_X1 i_718 (.CO (n_1437), .S (n_1436), .A (n_1430), .B (n_1393), .CI (n_1432));
FA_X1 i_717 (.CO (n_1435), .S (n_1434), .A (n_1389), .B (n_1428), .CI (n_1391));
FA_X1 i_716 (.CO (n_1433), .S (n_1432), .A (n_1426), .B (n_1424), .CI (n_1387));
FA_X1 i_715 (.CO (n_1431), .S (n_1430), .A (n_1422), .B (n_1420), .CI (n_1385));
FA_X1 i_714 (.CO (n_1429), .S (n_1428), .A (n_1381), .B (n_1418), .CI (n_1383));
FA_X1 i_713 (.CO (n_1427), .S (n_1426), .A (n_1412), .B (n_1379), .CI (n_1377));
FA_X1 i_712 (.CO (n_1425), .S (n_1424), .A (n_1375), .B (n_1416), .CI (n_1414));
FA_X1 i_711 (.CO (n_1423), .S (n_1422), .A (n_1402), .B (n_1400), .CI (n_1398));
FA_X1 i_710 (.CO (n_1421), .S (n_1420), .A (n_1408), .B (n_1406), .CI (n_1404));
FA_X1 i_709 (.CO (n_1419), .S (n_1418), .A (n_1371), .B (n_1369), .CI (n_1410));
FA_X1 i_708 (.CO (n_1417), .S (n_1416), .A (n_1357), .B (n_1355), .CI (n_1373));
FA_X1 i_707 (.CO (n_1415), .S (n_1414), .A (n_1363), .B (n_1361), .CI (n_1359));
FA_X1 i_706 (.CO (n_1413), .S (n_1412), .A (n_2531), .B (n_1367), .CI (n_1365));
FA_X1 i_705 (.CO (n_1411), .S (n_1410), .A (n_2438), .B (n_2469), .CI (n_2500));
FA_X1 i_704 (.CO (n_1409), .S (n_1408), .A (n_2345), .B (n_2376), .CI (n_2407));
FA_X1 i_703 (.CO (n_1407), .S (n_1406), .A (n_2252), .B (n_2283), .CI (n_2314));
FA_X1 i_702 (.CO (n_1405), .S (n_1404), .A (n_2159), .B (n_2190), .CI (n_2221));
FA_X1 i_701 (.CO (n_1403), .S (n_1402), .A (n_2066), .B (n_2097), .CI (n_2128));
FA_X1 i_700 (.CO (n_1401), .S (n_1400), .A (n_1973), .B (n_2004), .CI (n_2035));
FA_X1 i_699 (.CO (n_1399), .S (n_1398), .A (n_1880), .B (n_1911), .CI (n_1942));
FA_X1 i_698 (.CO (n_1397), .S (n_1396), .A (n_1392), .B (n_1351), .CI (n_1394));
FA_X1 i_697 (.CO (n_1395), .S (n_1394), .A (n_1388), .B (n_1390), .CI (n_1349));
FA_X1 i_696 (.CO (n_1393), .S (n_1392), .A (n_1345), .B (n_1386), .CI (n_1347));
FA_X1 i_695 (.CO (n_1391), .S (n_1390), .A (n_1384), .B (n_1382), .CI (n_1343));
FA_X1 i_694 (.CO (n_1389), .S (n_1388), .A (n_1378), .B (n_1376), .CI (n_1341));
FA_X1 i_693 (.CO (n_1387), .S (n_1386), .A (n_1339), .B (n_1337), .CI (n_1380));
FA_X1 i_692 (.CO (n_1385), .S (n_1384), .A (n_1333), .B (n_1331), .CI (n_1374));
FA_X1 i_691 (.CO (n_1383), .S (n_1382), .A (n_1372), .B (n_1370), .CI (n_1335));
FA_X1 i_690 (.CO (n_1381), .S (n_1380), .A (n_1356), .B (n_1354), .CI (n_1329));
FA_X1 i_689 (.CO (n_1379), .S (n_1378), .A (n_1362), .B (n_1360), .CI (n_1358));
FA_X1 i_688 (.CO (n_1377), .S (n_1376), .A (n_1368), .B (n_1366), .CI (n_1364));
FA_X1 i_687 (.CO (n_1375), .S (n_1374), .A (n_1309), .B (n_1327), .CI (n_1325));
FA_X1 i_686 (.CO (n_1373), .S (n_1372), .A (n_1315), .B (n_1313), .CI (n_1311));
FA_X1 i_685 (.CO (n_1371), .S (n_1370), .A (n_1321), .B (n_1319), .CI (n_1317));
FA_X1 i_684 (.CO (n_1369), .S (n_1368), .A (n_2532), .B (n_2563), .CI (n_1323));
FA_X1 i_683 (.CO (n_1367), .S (n_1366), .A (n_2439), .B (n_2470), .CI (n_2501));
FA_X1 i_682 (.CO (n_1365), .S (n_1364), .A (n_2346), .B (n_2377), .CI (n_2408));
FA_X1 i_681 (.CO (n_1363), .S (n_1362), .A (n_2253), .B (n_2284), .CI (n_2315));
FA_X1 i_680 (.CO (n_1361), .S (n_1360), .A (n_2160), .B (n_2191), .CI (n_2222));
FA_X1 i_679 (.CO (n_1359), .S (n_1358), .A (n_2067), .B (n_2098), .CI (n_2129));
FA_X1 i_678 (.CO (n_1357), .S (n_1356), .A (n_1974), .B (n_2005), .CI (n_2036));
FA_X1 i_677 (.CO (n_1355), .S (n_1354), .A (n_1881), .B (n_1912), .CI (n_1943));
FA_X1 i_676 (.CO (n_1353), .S (n_1352), .A (n_1348), .B (n_1305), .CI (n_1350));
FA_X1 i_675 (.CO (n_1351), .S (n_1350), .A (n_1301), .B (n_1346), .CI (n_1303));
FA_X1 i_674 (.CO (n_1349), .S (n_1348), .A (n_1342), .B (n_1299), .CI (n_1344));
FA_X1 i_673 (.CO (n_1347), .S (n_1346), .A (n_1338), .B (n_1297), .CI (n_1340));
FA_X1 i_672 (.CO (n_1345), .S (n_1344), .A (n_1332), .B (n_1336), .CI (n_1295));
FA_X1 i_671 (.CO (n_1343), .S (n_1342), .A (n_1293), .B (n_1291), .CI (n_1334));
FA_X1 i_670 (.CO (n_1341), .S (n_1340), .A (n_1285), .B (n_1289), .CI (n_1330));
FA_X1 i_669 (.CO (n_1339), .S (n_1338), .A (n_1326), .B (n_1324), .CI (n_1287));
FA_X1 i_668 (.CO (n_1337), .S (n_1336), .A (n_1308), .B (n_1283), .CI (n_1328));
FA_X1 i_667 (.CO (n_1335), .S (n_1334), .A (n_1314), .B (n_1312), .CI (n_1310));
FA_X1 i_666 (.CO (n_1333), .S (n_1332), .A (n_1320), .B (n_1318), .CI (n_1316));
FA_X1 i_665 (.CO (n_1331), .S (n_1330), .A (n_1279), .B (n_1277), .CI (n_1322));
FA_X1 i_664 (.CO (n_1329), .S (n_1328), .A (n_1263), .B (n_1261), .CI (n_1281));
FA_X1 i_663 (.CO (n_1327), .S (n_1326), .A (n_1269), .B (n_1267), .CI (n_1265));
FA_X1 i_662 (.CO (n_1325), .S (n_1324), .A (n_1275), .B (n_1273), .CI (n_1271));
FA_X1 i_661 (.CO (n_1323), .S (n_1322), .A (n_2533), .B (n_2564), .CI (n_2595));
FA_X1 i_660 (.CO (n_1321), .S (n_1320), .A (n_2440), .B (n_2471), .CI (n_2502));
FA_X1 i_659 (.CO (n_1319), .S (n_1318), .A (n_2347), .B (n_2378), .CI (n_2409));
FA_X1 i_658 (.CO (n_1317), .S (n_1316), .A (n_2254), .B (n_2285), .CI (n_2316));
FA_X1 i_657 (.CO (n_1315), .S (n_1314), .A (n_2161), .B (n_2192), .CI (n_2223));
FA_X1 i_656 (.CO (n_1313), .S (n_1312), .A (n_2068), .B (n_2099), .CI (n_2130));
FA_X1 i_655 (.CO (n_1311), .S (n_1310), .A (n_1975), .B (n_2006), .CI (n_2037));
FA_X1 i_654 (.CO (n_1309), .S (n_1308), .A (n_1882), .B (n_1913), .CI (n_1944));
FA_X1 i_653 (.CO (n_1307), .S (n_1306), .A (n_1257), .B (n_1302), .CI (n_1304));
FA_X1 i_652 (.CO (n_1305), .S (n_1304), .A (n_1253), .B (n_1300), .CI (n_1255));
FA_X1 i_651 (.CO (n_1303), .S (n_1302), .A (n_1251), .B (n_1296), .CI (n_1298));
FA_X1 i_650 (.CO (n_1301), .S (n_1300), .A (n_1290), .B (n_1249), .CI (n_1294));
FA_X1 i_649 (.CO (n_1299), .S (n_1298), .A (n_1284), .B (n_1247), .CI (n_1292));
FA_X1 i_648 (.CO (n_1297), .S (n_1296), .A (n_1243), .B (n_1288), .CI (n_1286));
FA_X1 i_647 (.CO (n_1295), .S (n_1294), .A (n_1241), .B (n_1282), .CI (n_1245));
FA_X1 i_646 (.CO (n_1293), .S (n_1292), .A (n_1239), .B (n_1237), .CI (n_1235));
FA_X1 i_645 (.CO (n_1291), .S (n_1290), .A (n_1280), .B (n_1278), .CI (n_1276));
FA_X1 i_644 (.CO (n_1289), .S (n_1288), .A (n_1262), .B (n_1260), .CI (n_1233));
FA_X1 i_643 (.CO (n_1287), .S (n_1286), .A (n_1268), .B (n_1266), .CI (n_1264));
FA_X1 i_642 (.CO (n_1285), .S (n_1284), .A (n_1274), .B (n_1272), .CI (n_1270));
FA_X1 i_641 (.CO (n_1283), .S (n_1282), .A (n_1231), .B (n_1229), .CI (n_1227));
FA_X1 i_640 (.CO (n_1281), .S (n_1280), .A (n_1215), .B (n_1213), .CI (n_1211));
FA_X1 i_639 (.CO (n_1279), .S (n_1278), .A (n_1221), .B (n_1219), .CI (n_1217));
FA_X1 i_638 (.CO (n_1277), .S (n_1276), .A (n_2627), .B (n_1225), .CI (n_1223));
FA_X1 i_637 (.CO (n_1275), .S (n_1274), .A (n_2534), .B (n_2565), .CI (n_2596));
FA_X1 i_636 (.CO (n_1273), .S (n_1272), .A (n_2441), .B (n_2472), .CI (n_2503));
FA_X1 i_635 (.CO (n_1271), .S (n_1270), .A (n_2348), .B (n_2379), .CI (n_2410));
FA_X1 i_634 (.CO (n_1269), .S (n_1268), .A (n_2255), .B (n_2286), .CI (n_2317));
FA_X1 i_633 (.CO (n_1267), .S (n_1266), .A (n_2162), .B (n_2193), .CI (n_2224));
FA_X1 i_632 (.CO (n_1265), .S (n_1264), .A (n_2069), .B (n_2100), .CI (n_2131));
FA_X1 i_631 (.CO (n_1263), .S (n_1262), .A (n_1976), .B (n_2007), .CI (n_2038));
FA_X1 i_630 (.CO (n_1261), .S (n_1260), .A (n_1883), .B (n_1914), .CI (n_1945));
FA_X1 i_629 (.CO (n_1259), .S (n_1258), .A (n_1254), .B (n_1207), .CI (n_1256));
FA_X1 i_628 (.CO (n_1257), .S (n_1256), .A (n_1250), .B (n_1252), .CI (n_1205));
FA_X1 i_627 (.CO (n_1255), .S (n_1254), .A (n_1201), .B (n_1248), .CI (n_1203));
FA_X1 i_626 (.CO (n_1253), .S (n_1252), .A (n_1197), .B (n_1199), .CI (n_1246));
FA_X1 i_625 (.CO (n_1251), .S (n_1250), .A (n_1195), .B (n_1244), .CI (n_1242));
FA_X1 i_624 (.CO (n_1249), .S (n_1248), .A (n_1240), .B (n_1238), .CI (n_1236));
FA_X1 i_623 (.CO (n_1247), .S (n_1246), .A (n_1234), .B (n_1193), .CI (n_1191));
FA_X1 i_622 (.CO (n_1245), .S (n_1244), .A (n_1189), .B (n_1187), .CI (n_1185));
FA_X1 i_621 (.CO (n_1243), .S (n_1242), .A (n_1232), .B (n_1230), .CI (n_1228));
FA_X1 i_620 (.CO (n_1241), .S (n_1240), .A (n_1212), .B (n_1210), .CI (n_1183));
FA_X1 i_619 (.CO (n_1239), .S (n_1238), .A (n_1218), .B (n_1216), .CI (n_1214));
FA_X1 i_618 (.CO (n_1237), .S (n_1236), .A (n_1224), .B (n_1222), .CI (n_1220));
FA_X1 i_617 (.CO (n_1235), .S (n_1234), .A (n_1179), .B (n_1177), .CI (n_1226));
FA_X1 i_616 (.CO (n_1233), .S (n_1232), .A (n_1161), .B (n_1159), .CI (n_1181));
FA_X1 i_615 (.CO (n_1231), .S (n_1230), .A (n_1167), .B (n_1165), .CI (n_1163));
FA_X1 i_614 (.CO (n_1229), .S (n_1228), .A (n_1173), .B (n_1171), .CI (n_1169));
FA_X1 i_613 (.CO (n_1227), .S (n_1226), .A (n_2628), .B (n_2659), .CI (n_1175));
FA_X1 i_612 (.CO (n_1225), .S (n_1224), .A (n_2535), .B (n_2566), .CI (n_2597));
FA_X1 i_611 (.CO (n_1223), .S (n_1222), .A (n_2442), .B (n_2473), .CI (n_2504));
FA_X1 i_610 (.CO (n_1221), .S (n_1220), .A (n_2349), .B (n_2380), .CI (n_2411));
FA_X1 i_609 (.CO (n_1219), .S (n_1218), .A (n_2256), .B (n_2287), .CI (n_2318));
FA_X1 i_608 (.CO (n_1217), .S (n_1216), .A (n_2163), .B (n_2194), .CI (n_2225));
FA_X1 i_607 (.CO (n_1215), .S (n_1214), .A (n_2070), .B (n_2101), .CI (n_2132));
FA_X1 i_606 (.CO (n_1213), .S (n_1212), .A (n_1977), .B (n_2008), .CI (n_2039));
FA_X1 i_605 (.CO (n_1211), .S (n_1210), .A (n_1884), .B (n_1915), .CI (n_1946));
FA_X1 i_604 (.CO (n_1209), .S (n_1208), .A (n_1204), .B (n_1155), .CI (n_1206));
FA_X1 i_603 (.CO (n_1207), .S (n_1206), .A (n_1200), .B (n_1202), .CI (n_1153));
FA_X1 i_602 (.CO (n_1205), .S (n_1204), .A (n_1149), .B (n_1198), .CI (n_1151));
FA_X1 i_601 (.CO (n_1203), .S (n_1202), .A (n_1194), .B (n_1147), .CI (n_1196));
FA_X1 i_600 (.CO (n_1201), .S (n_1200), .A (n_1192), .B (n_1190), .CI (n_1145));
FA_X1 i_599 (.CO (n_1199), .S (n_1198), .A (n_1186), .B (n_1184), .CI (n_1143));
FA_X1 i_598 (.CO (n_1197), .S (n_1196), .A (n_1141), .B (n_1139), .CI (n_1188));
FA_X1 i_597 (.CO (n_1195), .S (n_1194), .A (n_1131), .B (n_1137), .CI (n_1182));
FA_X1 i_596 (.CO (n_1193), .S (n_1192), .A (n_1176), .B (n_1135), .CI (n_1133));
FA_X1 i_595 (.CO (n_1191), .S (n_1190), .A (n_1129), .B (n_1180), .CI (n_1178));
FA_X1 i_594 (.CO (n_1189), .S (n_1188), .A (n_1162), .B (n_1160), .CI (n_1158));
FA_X1 i_593 (.CO (n_1187), .S (n_1186), .A (n_1168), .B (n_1166), .CI (n_1164));
FA_X1 i_592 (.CO (n_1185), .S (n_1184), .A (n_1174), .B (n_1172), .CI (n_1170));
FA_X1 i_591 (.CO (n_1183), .S (n_1182), .A (n_1127), .B (n_1125), .CI (n_1123));
FA_X1 i_590 (.CO (n_1181), .S (n_1180), .A (n_1109), .B (n_1107), .CI (n_1105));
FA_X1 i_589 (.CO (n_1179), .S (n_1178), .A (n_1115), .B (n_1113), .CI (n_1111));
FA_X1 i_588 (.CO (n_1177), .S (n_1176), .A (n_1121), .B (n_1119), .CI (n_1117));
FA_X1 i_587 (.CO (n_1175), .S (n_1174), .A (n_2629), .B (n_2660), .CI (n_2691));
FA_X1 i_586 (.CO (n_1173), .S (n_1172), .A (n_2536), .B (n_2567), .CI (n_2598));
FA_X1 i_585 (.CO (n_1171), .S (n_1170), .A (n_2443), .B (n_2474), .CI (n_2505));
FA_X1 i_584 (.CO (n_1169), .S (n_1168), .A (n_2350), .B (n_2381), .CI (n_2412));
FA_X1 i_583 (.CO (n_1167), .S (n_1166), .A (n_2257), .B (n_2288), .CI (n_2319));
FA_X1 i_582 (.CO (n_1165), .S (n_1164), .A (n_2164), .B (n_2195), .CI (n_2226));
FA_X1 i_581 (.CO (n_1163), .S (n_1162), .A (n_2071), .B (n_2102), .CI (n_2133));
FA_X1 i_580 (.CO (n_1161), .S (n_1160), .A (n_1978), .B (n_2009), .CI (n_2040));
FA_X1 i_579 (.CO (n_1159), .S (n_1158), .A (n_1885), .B (n_1916), .CI (n_1947));
FA_X1 i_578 (.CO (n_1157), .S (n_1156), .A (n_1152), .B (n_1101), .CI (n_1154));
FA_X1 i_577 (.CO (n_1155), .S (n_1154), .A (n_1097), .B (n_1150), .CI (n_1099));
FA_X1 i_576 (.CO (n_1153), .S (n_1152), .A (n_1144), .B (n_1146), .CI (n_1148));
FA_X1 i_575 (.CO (n_1151), .S (n_1150), .A (n_1142), .B (n_1095), .CI (n_1093));
FA_X1 i_574 (.CO (n_1149), .S (n_1148), .A (n_1140), .B (n_1138), .CI (n_1091));
FA_X1 i_573 (.CO (n_1147), .S (n_1146), .A (n_1134), .B (n_1132), .CI (n_1089));
FA_X1 i_572 (.CO (n_1145), .S (n_1144), .A (n_1083), .B (n_1087), .CI (n_1136));
FA_X1 i_571 (.CO (n_1143), .S (n_1142), .A (n_1130), .B (n_1128), .CI (n_1085));
FA_X1 i_570 (.CO (n_1141), .S (n_1140), .A (n_1081), .B (n_1079), .CI (n_1077));
FA_X1 i_569 (.CO (n_1139), .S (n_1138), .A (n_1126), .B (n_1124), .CI (n_1122));
FA_X1 i_568 (.CO (n_1137), .S (n_1136), .A (n_1106), .B (n_1104), .CI (n_1075));
FA_X1 i_567 (.CO (n_1135), .S (n_1134), .A (n_1112), .B (n_1110), .CI (n_1108));
FA_X1 i_566 (.CO (n_1133), .S (n_1132), .A (n_1118), .B (n_1116), .CI (n_1114));
FA_X1 i_565 (.CO (n_1131), .S (n_1130), .A (n_1069), .B (n_1067), .CI (n_1120));
FA_X1 i_564 (.CO (n_1129), .S (n_1128), .A (n_1049), .B (n_1073), .CI (n_1071));
FA_X1 i_563 (.CO (n_1127), .S (n_1126), .A (n_1055), .B (n_1053), .CI (n_1051));
FA_X1 i_562 (.CO (n_1125), .S (n_1124), .A (n_1061), .B (n_1059), .CI (n_1057));
FA_X1 i_561 (.CO (n_1123), .S (n_1122), .A (n_2723), .B (n_1065), .CI (n_1063));
FA_X1 i_560 (.CO (n_1121), .S (n_1120), .A (n_2630), .B (n_2661), .CI (n_2692));
FA_X1 i_559 (.CO (n_1119), .S (n_1118), .A (n_2537), .B (n_2568), .CI (n_2599));
FA_X1 i_558 (.CO (n_1117), .S (n_1116), .A (n_2444), .B (n_2475), .CI (n_2506));
FA_X1 i_557 (.CO (n_1115), .S (n_1114), .A (n_2351), .B (n_2382), .CI (n_2413));
FA_X1 i_556 (.CO (n_1113), .S (n_1112), .A (n_2258), .B (n_2289), .CI (n_2320));
FA_X1 i_555 (.CO (n_1111), .S (n_1110), .A (n_2165), .B (n_2196), .CI (n_2227));
FA_X1 i_554 (.CO (n_1109), .S (n_1108), .A (n_2072), .B (n_2103), .CI (n_2134));
FA_X1 i_553 (.CO (n_1107), .S (n_1106), .A (n_1979), .B (n_2010), .CI (n_2041));
FA_X1 i_552 (.CO (n_1105), .S (n_1104), .A (n_1886), .B (n_1917), .CI (n_1948));
FA_X1 i_551 (.CO (n_1103), .S (n_1102), .A (n_1098), .B (n_1045), .CI (n_1100));
FA_X1 i_550 (.CO (n_1101), .S (n_1100), .A (n_1041), .B (n_1096), .CI (n_1043));
FA_X1 i_549 (.CO (n_1099), .S (n_1098), .A (n_1092), .B (n_1039), .CI (n_1094));
FA_X1 i_548 (.CO (n_1097), .S (n_1096), .A (n_1088), .B (n_1037), .CI (n_1090));
FA_X1 i_547 (.CO (n_1095), .S (n_1094), .A (n_1084), .B (n_1035), .CI (n_1033));
FA_X1 i_546 (.CO (n_1093), .S (n_1092), .A (n_1082), .B (n_1031), .CI (n_1086));
FA_X1 i_545 (.CO (n_1091), .S (n_1090), .A (n_1080), .B (n_1078), .CI (n_1076));
FA_X1 i_544 (.CO (n_1089), .S (n_1088), .A (n_1074), .B (n_1029), .CI (n_1027));
FA_X1 i_543 (.CO (n_1087), .S (n_1086), .A (n_1021), .B (n_1019), .CI (n_1025));
FA_X1 i_542 (.CO (n_1085), .S (n_1084), .A (n_1070), .B (n_1068), .CI (n_1023));
FA_X1 i_541 (.CO (n_1083), .S (n_1082), .A (n_1048), .B (n_1017), .CI (n_1072));
FA_X1 i_540 (.CO (n_1081), .S (n_1080), .A (n_1054), .B (n_1052), .CI (n_1050));
FA_X1 i_539 (.CO (n_1079), .S (n_1078), .A (n_1060), .B (n_1058), .CI (n_1056));
FA_X1 i_538 (.CO (n_1077), .S (n_1076), .A (n_1066), .B (n_1064), .CI (n_1062));
FA_X1 i_537 (.CO (n_1075), .S (n_1074), .A (n_1015), .B (n_1013), .CI (n_1011));
FA_X1 i_536 (.CO (n_1073), .S (n_1072), .A (n_995), .B (n_993), .CI (n_991));
FA_X1 i_535 (.CO (n_1071), .S (n_1070), .A (n_1001), .B (n_999), .CI (n_997));
FA_X1 i_534 (.CO (n_1069), .S (n_1068), .A (n_1007), .B (n_1005), .CI (n_1003));
FA_X1 i_533 (.CO (n_1067), .S (n_1066), .A (n_2724), .B (n_2755), .CI (n_1009));
FA_X1 i_532 (.CO (n_1065), .S (n_1064), .A (n_2631), .B (n_2662), .CI (n_2693));
FA_X1 i_531 (.CO (n_1063), .S (n_1062), .A (n_2538), .B (n_2569), .CI (n_2600));
FA_X1 i_530 (.CO (n_1061), .S (n_1060), .A (n_2445), .B (n_2476), .CI (n_2507));
FA_X1 i_529 (.CO (n_1059), .S (n_1058), .A (n_2352), .B (n_2383), .CI (n_2414));
FA_X1 i_528 (.CO (n_1057), .S (n_1056), .A (n_2259), .B (n_2290), .CI (n_2321));
FA_X1 i_527 (.CO (n_1055), .S (n_1054), .A (n_2166), .B (n_2197), .CI (n_2228));
FA_X1 i_526 (.CO (n_1053), .S (n_1052), .A (n_2073), .B (n_2104), .CI (n_2135));
FA_X1 i_525 (.CO (n_1051), .S (n_1050), .A (n_1980), .B (n_2011), .CI (n_2042));
FA_X1 i_524 (.CO (n_1049), .S (n_1048), .A (n_1887), .B (n_1918), .CI (n_1949));
FA_X1 i_523 (.CO (n_1047), .S (n_1046), .A (n_1042), .B (n_1044), .CI (n_987));
FA_X1 i_522 (.CO (n_1045), .S (n_1044), .A (n_983), .B (n_1040), .CI (n_985));
FA_X1 i_521 (.CO (n_1043), .S (n_1042), .A (n_981), .B (n_1036), .CI (n_1038));
FA_X1 i_520 (.CO (n_1041), .S (n_1040), .A (n_1030), .B (n_979), .CI (n_1034));
FA_X1 i_519 (.CO (n_1039), .S (n_1038), .A (n_975), .B (n_977), .CI (n_1032));
FA_X1 i_518 (.CO (n_1037), .S (n_1036), .A (n_973), .B (n_1028), .CI (n_1026));
FA_X1 i_517 (.CO (n_1035), .S (n_1034), .A (n_1022), .B (n_1020), .CI (n_1018));
FA_X1 i_516 (.CO (n_1033), .S (n_1032), .A (n_969), .B (n_967), .CI (n_1024));
FA_X1 i_515 (.CO (n_1031), .S (n_1030), .A (n_961), .B (n_1016), .CI (n_971));
FA_X1 i_514 (.CO (n_1029), .S (n_1028), .A (n_1010), .B (n_965), .CI (n_963));
FA_X1 i_513 (.CO (n_1027), .S (n_1026), .A (n_957), .B (n_1014), .CI (n_1012));
FA_X1 i_512 (.CO (n_1025), .S (n_1024), .A (n_992), .B (n_990), .CI (n_959));
FA_X1 i_511 (.CO (n_1023), .S (n_1022), .A (n_998), .B (n_996), .CI (n_994));
FA_X1 i_510 (.CO (n_1021), .S (n_1020), .A (n_1004), .B (n_1002), .CI (n_1000));
FA_X1 i_509 (.CO (n_1019), .S (n_1018), .A (n_951), .B (n_1008), .CI (n_1006));
FA_X1 i_508 (.CO (n_1017), .S (n_1016), .A (n_931), .B (n_955), .CI (n_953));
FA_X1 i_507 (.CO (n_1015), .S (n_1014), .A (n_937), .B (n_935), .CI (n_933));
FA_X1 i_506 (.CO (n_1013), .S (n_1012), .A (n_943), .B (n_941), .CI (n_939));
FA_X1 i_505 (.CO (n_1011), .S (n_1010), .A (n_949), .B (n_947), .CI (n_945));
FA_X1 i_504 (.CO (n_1009), .S (n_1008), .A (n_2725), .B (n_2756), .CI (n_2787));
FA_X1 i_503 (.CO (n_1007), .S (n_1006), .A (n_2632), .B (n_2663), .CI (n_2694));
FA_X1 i_502 (.CO (n_1005), .S (n_1004), .A (n_2539), .B (n_2570), .CI (n_2601));
FA_X1 i_501 (.CO (n_1003), .S (n_1002), .A (n_2446), .B (n_2477), .CI (n_2508));
FA_X1 i_500 (.CO (n_1001), .S (n_1000), .A (n_2353), .B (n_2384), .CI (n_2415));
FA_X1 i_499 (.CO (n_999), .S (n_998), .A (n_2260), .B (n_2291), .CI (n_2322));
FA_X1 i_498 (.CO (n_997), .S (n_996), .A (n_2167), .B (n_2198), .CI (n_2229));
FA_X1 i_497 (.CO (n_995), .S (n_994), .A (n_2074), .B (n_2105), .CI (n_2136));
FA_X1 i_496 (.CO (n_993), .S (n_992), .A (n_1981), .B (n_2012), .CI (n_2043));
FA_X1 i_495 (.CO (n_991), .S (n_990), .A (n_1888), .B (n_1919), .CI (n_1950));
HA_X1 i_494 (.CO (n_989), .S (n_988), .A (n_927), .B (n_986));
FA_X1 i_493 (.CO (n_987), .S (n_986), .A (n_982), .B (n_925), .CI (n_984));
FA_X1 i_492 (.CO (n_985), .S (n_984), .A (n_978), .B (n_923), .CI (n_980));
FA_X1 i_491 (.CO (n_983), .S (n_982), .A (n_974), .B (n_976), .CI (n_921));
FA_X1 i_490 (.CO (n_981), .S (n_980), .A (n_917), .B (n_972), .CI (n_919));
FA_X1 i_489 (.CO (n_979), .S (n_978), .A (n_970), .B (n_968), .CI (n_915));
FA_X1 i_488 (.CO (n_977), .S (n_976), .A (n_960), .B (n_966), .CI (n_913));
FA_X1 i_487 (.CO (n_975), .S (n_974), .A (n_909), .B (n_964), .CI (n_962));
FA_X1 i_486 (.CO (n_973), .S (n_972), .A (n_907), .B (n_958), .CI (n_911));
FA_X1 i_485 (.CO (n_971), .S (n_970), .A (n_905), .B (n_903), .CI (n_901));
FA_X1 i_484 (.CO (n_969), .S (n_968), .A (n_954), .B (n_952), .CI (n_950));
FA_X1 i_483 (.CO (n_967), .S (n_966), .A (n_930), .B (n_899), .CI (n_956));
FA_X1 i_482 (.CO (n_965), .S (n_964), .A (n_936), .B (n_934), .CI (n_932));
FA_X1 i_481 (.CO (n_963), .S (n_962), .A (n_942), .B (n_940), .CI (n_938));
FA_X1 i_480 (.CO (n_961), .S (n_960), .A (n_948), .B (n_946), .CI (n_944));
FA_X1 i_479 (.CO (n_959), .S (n_958), .A (n_895), .B (n_893), .CI (n_891));
FA_X1 i_478 (.CO (n_957), .S (n_956), .A (n_873), .B (n_871), .CI (n_897));
FA_X1 i_477 (.CO (n_955), .S (n_954), .A (n_879), .B (n_877), .CI (n_875));
FA_X1 i_476 (.CO (n_953), .S (n_952), .A (n_885), .B (n_883), .CI (n_881));
FA_X1 i_475 (.CO (n_951), .S (n_950), .A (n_2819), .B (n_889), .CI (n_887));
FA_X1 i_474 (.CO (n_949), .S (n_948), .A (n_2726), .B (n_2757), .CI (n_2788));
FA_X1 i_473 (.CO (n_947), .S (n_946), .A (n_2633), .B (n_2664), .CI (n_2695));
FA_X1 i_472 (.CO (n_945), .S (n_944), .A (n_2540), .B (n_2571), .CI (n_2602));
FA_X1 i_471 (.CO (n_943), .S (n_942), .A (n_2447), .B (n_2478), .CI (n_2509));
FA_X1 i_470 (.CO (n_941), .S (n_940), .A (n_2354), .B (n_2385), .CI (n_2416));
FA_X1 i_469 (.CO (n_939), .S (n_938), .A (n_2261), .B (n_2292), .CI (n_2323));
FA_X1 i_468 (.CO (n_937), .S (n_936), .A (n_2168), .B (n_2199), .CI (n_2230));
FA_X1 i_467 (.CO (n_935), .S (n_934), .A (n_2075), .B (n_2106), .CI (n_2137));
FA_X1 i_466 (.CO (n_933), .S (n_932), .A (n_1982), .B (n_2013), .CI (n_2044));
FA_X1 i_465 (.CO (n_931), .S (n_930), .A (n_1889), .B (n_1920), .CI (n_1951));
HA_X1 i_464 (.CO (n_929), .S (n_928), .A (n_867), .B (n_926));
FA_X1 i_463 (.CO (n_927), .S (n_926), .A (n_865), .B (n_922), .CI (n_924));
FA_X1 i_462 (.CO (n_925), .S (n_924), .A (n_918), .B (n_863), .CI (n_920));
FA_X1 i_461 (.CO (n_923), .S (n_922), .A (n_916), .B (n_914), .CI (n_861));
FA_X1 i_460 (.CO (n_921), .S (n_920), .A (n_857), .B (n_912), .CI (n_859));
FA_X1 i_459 (.CO (n_919), .S (n_918), .A (n_853), .B (n_910), .CI (n_908));
FA_X1 i_458 (.CO (n_917), .S (n_916), .A (n_902), .B (n_900), .CI (n_855));
FA_X1 i_457 (.CO (n_915), .S (n_914), .A (n_849), .B (n_906), .CI (n_904));
FA_X1 i_456 (.CO (n_913), .S (n_912), .A (n_841), .B (n_898), .CI (n_851));
FA_X1 i_455 (.CO (n_911), .S (n_910), .A (n_847), .B (n_845), .CI (n_843));
FA_X1 i_454 (.CO (n_909), .S (n_908), .A (n_896), .B (n_894), .CI (n_892));
FA_X1 i_453 (.CO (n_907), .S (n_906), .A (n_872), .B (n_870), .CI (n_839));
FA_X1 i_452 (.CO (n_905), .S (n_904), .A (n_878), .B (n_876), .CI (n_874));
FA_X1 i_451 (.CO (n_903), .S (n_902), .A (n_884), .B (n_882), .CI (n_880));
FA_X1 i_450 (.CO (n_901), .S (n_900), .A (n_890), .B (n_888), .CI (n_886));
FA_X1 i_449 (.CO (n_899), .S (n_898), .A (n_837), .B (n_835), .CI (n_833));
FA_X1 i_448 (.CO (n_897), .S (n_896), .A (n_817), .B (n_815), .CI (n_813));
FA_X1 i_447 (.CO (n_895), .S (n_894), .A (n_823), .B (n_821), .CI (n_819));
FA_X1 i_446 (.CO (n_893), .S (n_892), .A (n_829), .B (n_827), .CI (n_825));
FA_X1 i_445 (.CO (n_891), .S (n_890), .A (n_2820), .B (n_2849), .CI (n_831));
FA_X1 i_444 (.CO (n_889), .S (n_888), .A (n_2727), .B (n_2758), .CI (n_2789));
FA_X1 i_443 (.CO (n_887), .S (n_886), .A (n_2634), .B (n_2665), .CI (n_2696));
FA_X1 i_442 (.CO (n_885), .S (n_884), .A (n_2541), .B (n_2572), .CI (n_2603));
FA_X1 i_441 (.CO (n_883), .S (n_882), .A (n_2448), .B (n_2479), .CI (n_2510));
FA_X1 i_440 (.CO (n_881), .S (n_880), .A (n_2355), .B (n_2386), .CI (n_2417));
FA_X1 i_439 (.CO (n_879), .S (n_878), .A (n_2262), .B (n_2293), .CI (n_2324));
FA_X1 i_438 (.CO (n_877), .S (n_876), .A (n_2169), .B (n_2200), .CI (n_2231));
FA_X1 i_437 (.CO (n_875), .S (n_874), .A (n_2076), .B (n_2107), .CI (n_2138));
FA_X1 i_436 (.CO (n_873), .S (n_872), .A (n_1983), .B (n_2014), .CI (n_2045));
FA_X1 i_435 (.CO (n_871), .S (n_870), .A (n_1890), .B (n_1921), .CI (n_1952));
HA_X1 i_434 (.CO (n_869), .S (n_868), .A (n_809), .B (n_866));
FA_X1 i_433 (.CO (n_867), .S (n_866), .A (n_807), .B (n_862), .CI (n_864));
FA_X1 i_432 (.CO (n_865), .S (n_864), .A (n_860), .B (n_858), .CI (n_805));
FA_X1 i_431 (.CO (n_863), .S (n_862), .A (n_801), .B (n_856), .CI (n_803));
FA_X1 i_430 (.CO (n_861), .S (n_860), .A (n_848), .B (n_799), .CI (n_854));
FA_X1 i_429 (.CO (n_859), .S (n_858), .A (n_797), .B (n_852), .CI (n_850));
FA_X1 i_428 (.CO (n_857), .S (n_856), .A (n_846), .B (n_844), .CI (n_842));
FA_X1 i_427 (.CO (n_855), .S (n_854), .A (n_795), .B (n_793), .CI (n_791));
FA_X1 i_426 (.CO (n_853), .S (n_852), .A (n_787), .B (n_785), .CI (n_840));
FA_X1 i_425 (.CO (n_851), .S (n_850), .A (n_834), .B (n_832), .CI (n_789));
FA_X1 i_424 (.CO (n_849), .S (n_848), .A (n_783), .B (n_838), .CI (n_836));
FA_X1 i_423 (.CO (n_847), .S (n_846), .A (n_816), .B (n_814), .CI (n_812));
FA_X1 i_422 (.CO (n_845), .S (n_844), .A (n_822), .B (n_820), .CI (n_818));
FA_X1 i_421 (.CO (n_843), .S (n_842), .A (n_828), .B (n_826), .CI (n_824));
FA_X1 i_420 (.CO (n_841), .S (n_840), .A (n_779), .B (n_777), .CI (n_830));
FA_X1 i_419 (.CO (n_839), .S (n_838), .A (n_759), .B (n_757), .CI (n_781));
FA_X1 i_418 (.CO (n_837), .S (n_836), .A (n_765), .B (n_763), .CI (n_761));
FA_X1 i_417 (.CO (n_835), .S (n_834), .A (n_771), .B (n_769), .CI (n_767));
FA_X1 i_416 (.CO (n_833), .S (n_832), .A (n_2850), .B (n_775), .CI (n_773));
FA_X1 i_415 (.CO (n_831), .S (n_830), .A (n_2759), .B (n_2790), .CI (n_2821));
FA_X1 i_414 (.CO (n_829), .S (n_828), .A (n_2666), .B (n_2697), .CI (n_2728));
FA_X1 i_413 (.CO (n_827), .S (n_826), .A (n_2573), .B (n_2604), .CI (n_2635));
FA_X1 i_412 (.CO (n_825), .S (n_824), .A (n_2480), .B (n_2511), .CI (n_2542));
FA_X1 i_411 (.CO (n_823), .S (n_822), .A (n_2387), .B (n_2418), .CI (n_2449));
FA_X1 i_410 (.CO (n_821), .S (n_820), .A (n_2294), .B (n_2325), .CI (n_2356));
FA_X1 i_409 (.CO (n_819), .S (n_818), .A (n_2201), .B (n_2232), .CI (n_2263));
FA_X1 i_408 (.CO (n_817), .S (n_816), .A (n_2108), .B (n_2139), .CI (n_2170));
FA_X1 i_407 (.CO (n_815), .S (n_814), .A (n_2015), .B (n_2046), .CI (n_2077));
FA_X1 i_406 (.CO (n_813), .S (n_812), .A (n_1922), .B (n_1953), .CI (n_1984));
HA_X1 i_405 (.CO (n_811), .S (n_810), .A (n_753), .B (n_808));
FA_X1 i_404 (.CO (n_809), .S (n_808), .A (n_751), .B (n_804), .CI (n_806));
FA_X1 i_403 (.CO (n_807), .S (n_806), .A (n_800), .B (n_802), .CI (n_749));
FA_X1 i_402 (.CO (n_805), .S (n_804), .A (n_745), .B (n_747), .CI (n_798));
FA_X1 i_401 (.CO (n_803), .S (n_802), .A (n_792), .B (n_743), .CI (n_796));
FA_X1 i_400 (.CO (n_801), .S (n_800), .A (n_790), .B (n_741), .CI (n_794));
FA_X1 i_399 (.CO (n_799), .S (n_798), .A (n_788), .B (n_786), .CI (n_784));
FA_X1 i_398 (.CO (n_797), .S (n_796), .A (n_782), .B (n_739), .CI (n_737));
FA_X1 i_397 (.CO (n_795), .S (n_794), .A (n_733), .B (n_731), .CI (n_729));
FA_X1 i_396 (.CO (n_793), .S (n_792), .A (n_778), .B (n_776), .CI (n_735));
FA_X1 i_395 (.CO (n_791), .S (n_790), .A (n_756), .B (n_727), .CI (n_780));
FA_X1 i_394 (.CO (n_789), .S (n_788), .A (n_762), .B (n_760), .CI (n_758));
FA_X1 i_393 (.CO (n_787), .S (n_786), .A (n_768), .B (n_766), .CI (n_764));
FA_X1 i_392 (.CO (n_785), .S (n_784), .A (n_774), .B (n_772), .CI (n_770));
FA_X1 i_391 (.CO (n_783), .S (n_782), .A (n_725), .B (n_723), .CI (n_721));
FA_X1 i_390 (.CO (n_781), .S (n_780), .A (n_707), .B (n_705), .CI (n_703));
FA_X1 i_389 (.CO (n_779), .S (n_778), .A (n_713), .B (n_711), .CI (n_709));
FA_X1 i_388 (.CO (n_777), .S (n_776), .A (n_719), .B (n_717), .CI (n_715));
FA_X1 i_387 (.CO (n_775), .S (n_774), .A (n_2791), .B (n_2822), .CI (n_2851));
FA_X1 i_386 (.CO (n_773), .S (n_772), .A (n_2698), .B (n_2729), .CI (n_2760));
FA_X1 i_385 (.CO (n_771), .S (n_770), .A (n_2605), .B (n_2636), .CI (n_2667));
FA_X1 i_384 (.CO (n_769), .S (n_768), .A (n_2512), .B (n_2543), .CI (n_2574));
FA_X1 i_383 (.CO (n_767), .S (n_766), .A (n_2419), .B (n_2450), .CI (n_2481));
FA_X1 i_382 (.CO (n_765), .S (n_764), .A (n_2326), .B (n_2357), .CI (n_2388));
FA_X1 i_381 (.CO (n_763), .S (n_762), .A (n_2233), .B (n_2264), .CI (n_2295));
FA_X1 i_380 (.CO (n_761), .S (n_760), .A (n_2140), .B (n_2171), .CI (n_2202));
FA_X1 i_379 (.CO (n_759), .S (n_758), .A (n_2047), .B (n_2078), .CI (n_2109));
FA_X1 i_378 (.CO (n_757), .S (n_756), .A (n_1954), .B (n_1985), .CI (n_2016));
HA_X1 i_377 (.CO (n_755), .S (n_754), .A (n_699), .B (n_752));
FA_X1 i_376 (.CO (n_753), .S (n_752), .A (n_748), .B (n_697), .CI (n_750));
FA_X1 i_375 (.CO (n_751), .S (n_750), .A (n_744), .B (n_695), .CI (n_746));
FA_X1 i_374 (.CO (n_749), .S (n_748), .A (n_740), .B (n_693), .CI (n_742));
FA_X1 i_373 (.CO (n_747), .S (n_746), .A (n_736), .B (n_689), .CI (n_691));
FA_X1 i_372 (.CO (n_745), .S (n_744), .A (n_730), .B (n_687), .CI (n_738));
FA_X1 i_371 (.CO (n_743), .S (n_742), .A (n_683), .B (n_734), .CI (n_732));
FA_X1 i_370 (.CO (n_741), .S (n_740), .A (n_677), .B (n_728), .CI (n_685));
FA_X1 i_369 (.CO (n_739), .S (n_738), .A (n_722), .B (n_681), .CI (n_679));
FA_X1 i_368 (.CO (n_737), .S (n_736), .A (n_675), .B (n_726), .CI (n_724));
FA_X1 i_367 (.CO (n_735), .S (n_734), .A (n_706), .B (n_704), .CI (n_702));
FA_X1 i_366 (.CO (n_733), .S (n_732), .A (n_712), .B (n_710), .CI (n_708));
FA_X1 i_365 (.CO (n_731), .S (n_730), .A (n_718), .B (n_716), .CI (n_714));
FA_X1 i_364 (.CO (n_729), .S (n_728), .A (n_671), .B (n_669), .CI (n_720));
FA_X1 i_363 (.CO (n_727), .S (n_726), .A (n_653), .B (n_651), .CI (n_673));
FA_X1 i_362 (.CO (n_725), .S (n_724), .A (n_659), .B (n_657), .CI (n_655));
FA_X1 i_361 (.CO (n_723), .S (n_722), .A (n_665), .B (n_663), .CI (n_661));
FA_X1 i_360 (.CO (n_721), .S (n_720), .A (n_2823), .B (n_2852), .CI (n_667));
FA_X1 i_359 (.CO (n_719), .S (n_718), .A (n_2730), .B (n_2761), .CI (n_2792));
FA_X1 i_358 (.CO (n_717), .S (n_716), .A (n_2637), .B (n_2668), .CI (n_2699));
FA_X1 i_357 (.CO (n_715), .S (n_714), .A (n_2544), .B (n_2575), .CI (n_2606));
FA_X1 i_356 (.CO (n_713), .S (n_712), .A (n_2451), .B (n_2482), .CI (n_2513));
FA_X1 i_355 (.CO (n_711), .S (n_710), .A (n_2358), .B (n_2389), .CI (n_2420));
FA_X1 i_354 (.CO (n_709), .S (n_708), .A (n_2265), .B (n_2296), .CI (n_2327));
FA_X1 i_353 (.CO (n_707), .S (n_706), .A (n_2172), .B (n_2203), .CI (n_2234));
FA_X1 i_352 (.CO (n_705), .S (n_704), .A (n_2079), .B (n_2110), .CI (n_2141));
FA_X1 i_351 (.CO (n_703), .S (n_702), .A (n_1986), .B (n_2017), .CI (n_2048));
HA_X1 i_350 (.CO (n_701), .S (n_700), .A (n_647), .B (n_698));
FA_X1 i_349 (.CO (n_699), .S (n_698), .A (n_694), .B (n_645), .CI (n_696));
FA_X1 i_348 (.CO (n_697), .S (n_696), .A (n_690), .B (n_643), .CI (n_692));
FA_X1 i_347 (.CO (n_695), .S (n_694), .A (n_686), .B (n_688), .CI (n_641));
FA_X1 i_346 (.CO (n_693), .S (n_692), .A (n_684), .B (n_682), .CI (n_639));
FA_X1 i_345 (.CO (n_691), .S (n_690), .A (n_678), .B (n_676), .CI (n_637));
FA_X1 i_344 (.CO (n_689), .S (n_688), .A (n_635), .B (n_633), .CI (n_680));
FA_X1 i_343 (.CO (n_687), .S (n_686), .A (n_625), .B (n_631), .CI (n_674));
FA_X1 i_342 (.CO (n_685), .S (n_684), .A (n_668), .B (n_629), .CI (n_627));
FA_X1 i_341 (.CO (n_683), .S (n_682), .A (n_623), .B (n_672), .CI (n_670));
FA_X1 i_340 (.CO (n_681), .S (n_680), .A (n_654), .B (n_652), .CI (n_650));
FA_X1 i_339 (.CO (n_679), .S (n_678), .A (n_660), .B (n_658), .CI (n_656));
FA_X1 i_338 (.CO (n_677), .S (n_676), .A (n_666), .B (n_664), .CI (n_662));
FA_X1 i_337 (.CO (n_675), .S (n_674), .A (n_601), .B (n_621), .CI (n_619));
FA_X1 i_336 (.CO (n_673), .S (n_672), .A (n_607), .B (n_605), .CI (n_603));
FA_X1 i_335 (.CO (n_671), .S (n_670), .A (n_613), .B (n_611), .CI (n_609));
FA_X1 i_334 (.CO (n_669), .S (n_668), .A (n_2853), .B (n_617), .CI (n_615));
FA_X1 i_333 (.CO (n_667), .S (n_666), .A (n_2762), .B (n_2793), .CI (n_2824));
FA_X1 i_332 (.CO (n_665), .S (n_664), .A (n_2669), .B (n_2700), .CI (n_2731));
FA_X1 i_331 (.CO (n_663), .S (n_662), .A (n_2576), .B (n_2607), .CI (n_2638));
FA_X1 i_330 (.CO (n_661), .S (n_660), .A (n_2483), .B (n_2514), .CI (n_2545));
FA_X1 i_329 (.CO (n_659), .S (n_658), .A (n_2390), .B (n_2421), .CI (n_2452));
FA_X1 i_328 (.CO (n_657), .S (n_656), .A (n_2297), .B (n_2328), .CI (n_2359));
FA_X1 i_327 (.CO (n_655), .S (n_654), .A (n_2204), .B (n_2235), .CI (n_2266));
FA_X1 i_326 (.CO (n_653), .S (n_652), .A (n_2111), .B (n_2142), .CI (n_2173));
FA_X1 i_325 (.CO (n_651), .S (n_650), .A (n_2018), .B (n_2049), .CI (n_2080));
HA_X1 i_324 (.CO (n_649), .S (n_648), .A (n_597), .B (n_646));
FA_X1 i_323 (.CO (n_647), .S (n_646), .A (n_642), .B (n_595), .CI (n_644));
FA_X1 i_322 (.CO (n_645), .S (n_644), .A (n_638), .B (n_593), .CI (n_640));
FA_X1 i_321 (.CO (n_643), .S (n_642), .A (n_589), .B (n_636), .CI (n_591));
FA_X1 i_320 (.CO (n_641), .S (n_640), .A (n_587), .B (n_634), .CI (n_632));
FA_X1 i_319 (.CO (n_639), .S (n_638), .A (n_630), .B (n_628), .CI (n_626));
FA_X1 i_318 (.CO (n_637), .S (n_636), .A (n_624), .B (n_585), .CI (n_583));
FA_X1 i_317 (.CO (n_635), .S (n_634), .A (n_581), .B (n_579), .CI (n_577));
FA_X1 i_316 (.CO (n_633), .S (n_632), .A (n_622), .B (n_620), .CI (n_618));
FA_X1 i_315 (.CO (n_631), .S (n_630), .A (n_602), .B (n_600), .CI (n_575));
FA_X1 i_314 (.CO (n_629), .S (n_628), .A (n_608), .B (n_606), .CI (n_604));
FA_X1 i_313 (.CO (n_627), .S (n_626), .A (n_614), .B (n_612), .CI (n_610));
FA_X1 i_312 (.CO (n_625), .S (n_624), .A (n_571), .B (n_569), .CI (n_616));
FA_X1 i_311 (.CO (n_623), .S (n_622), .A (n_555), .B (n_553), .CI (n_573));
FA_X1 i_310 (.CO (n_621), .S (n_620), .A (n_561), .B (n_559), .CI (n_557));
FA_X1 i_309 (.CO (n_619), .S (n_618), .A (n_567), .B (n_565), .CI (n_563));
FA_X1 i_308 (.CO (n_617), .S (n_616), .A (n_2794), .B (n_2825), .CI (n_2854));
FA_X1 i_307 (.CO (n_615), .S (n_614), .A (n_2701), .B (n_2732), .CI (n_2763));
FA_X1 i_306 (.CO (n_613), .S (n_612), .A (n_2608), .B (n_2639), .CI (n_2670));
FA_X1 i_305 (.CO (n_611), .S (n_610), .A (n_2515), .B (n_2546), .CI (n_2577));
FA_X1 i_304 (.CO (n_609), .S (n_608), .A (n_2422), .B (n_2453), .CI (n_2484));
FA_X1 i_303 (.CO (n_607), .S (n_606), .A (n_2329), .B (n_2360), .CI (n_2391));
FA_X1 i_302 (.CO (n_605), .S (n_604), .A (n_2236), .B (n_2267), .CI (n_2298));
FA_X1 i_301 (.CO (n_603), .S (n_602), .A (n_2143), .B (n_2174), .CI (n_2205));
FA_X1 i_300 (.CO (n_601), .S (n_600), .A (n_2050), .B (n_2081), .CI (n_2112));
HA_X1 i_299 (.CO (n_599), .S (n_598), .A (n_549), .B (n_551));
FA_X1 i_298 (.CO (n_597), .S (n_596), .A (n_547), .B (n_592), .CI (n_594));
FA_X1 i_297 (.CO (n_595), .S (n_594), .A (n_545), .B (n_588), .CI (n_590));
FA_X1 i_296 (.CO (n_593), .S (n_592), .A (n_541), .B (n_586), .CI (n_543));
FA_X1 i_295 (.CO (n_591), .S (n_590), .A (n_539), .B (n_584), .CI (n_582));
FA_X1 i_294 (.CO (n_589), .S (n_588), .A (n_580), .B (n_578), .CI (n_576));
FA_X1 i_293 (.CO (n_587), .S (n_586), .A (n_574), .B (n_537), .CI (n_535));
FA_X1 i_292 (.CO (n_585), .S (n_584), .A (n_533), .B (n_531), .CI (n_529));
FA_X1 i_291 (.CO (n_583), .S (n_582), .A (n_552), .B (n_572), .CI (n_570));
FA_X1 i_290 (.CO (n_581), .S (n_580), .A (n_558), .B (n_556), .CI (n_554));
FA_X1 i_289 (.CO (n_579), .S (n_578), .A (n_564), .B (n_562), .CI (n_560));
FA_X1 i_288 (.CO (n_577), .S (n_576), .A (n_523), .B (n_568), .CI (n_566));
FA_X1 i_287 (.CO (n_575), .S (n_574), .A (n_507), .B (n_527), .CI (n_525));
FA_X1 i_286 (.CO (n_573), .S (n_572), .A (n_513), .B (n_511), .CI (n_509));
FA_X1 i_285 (.CO (n_571), .S (n_570), .A (n_519), .B (n_517), .CI (n_515));
FA_X1 i_284 (.CO (n_569), .S (n_568), .A (n_2826), .B (n_2855), .CI (n_521));
FA_X1 i_283 (.CO (n_567), .S (n_566), .A (n_2733), .B (n_2764), .CI (n_2795));
FA_X1 i_282 (.CO (n_565), .S (n_564), .A (n_2640), .B (n_2671), .CI (n_2702));
FA_X1 i_281 (.CO (n_563), .S (n_562), .A (n_2547), .B (n_2578), .CI (n_2609));
FA_X1 i_280 (.CO (n_561), .S (n_560), .A (n_2454), .B (n_2485), .CI (n_2516));
FA_X1 i_279 (.CO (n_559), .S (n_558), .A (n_2361), .B (n_2392), .CI (n_2423));
FA_X1 i_278 (.CO (n_557), .S (n_556), .A (n_2268), .B (n_2299), .CI (n_2330));
FA_X1 i_277 (.CO (n_555), .S (n_554), .A (n_2175), .B (n_2206), .CI (n_2237));
FA_X1 i_276 (.CO (n_553), .S (n_552), .A (n_2082), .B (n_2113), .CI (n_2144));
HA_X1 i_275 (.CO (n_551), .S (n_550), .A (n_503), .B (n_548));
FA_X1 i_274 (.CO (n_549), .S (n_548), .A (n_544), .B (n_501), .CI (n_546));
FA_X1 i_273 (.CO (n_547), .S (n_546), .A (n_499), .B (n_540), .CI (n_542));
FA_X1 i_272 (.CO (n_545), .S (n_544), .A (n_536), .B (n_495), .CI (n_497));
FA_X1 i_271 (.CO (n_543), .S (n_542), .A (n_534), .B (n_493), .CI (n_538));
FA_X1 i_270 (.CO (n_541), .S (n_540), .A (n_491), .B (n_532), .CI (n_530));
FA_X1 i_269 (.CO (n_539), .S (n_538), .A (n_487), .B (n_485), .CI (n_528));
FA_X1 i_268 (.CO (n_537), .S (n_536), .A (n_524), .B (n_522), .CI (n_489));
FA_X1 i_267 (.CO (n_535), .S (n_534), .A (n_506), .B (n_483), .CI (n_526));
FA_X1 i_266 (.CO (n_533), .S (n_532), .A (n_512), .B (n_510), .CI (n_508));
FA_X1 i_265 (.CO (n_531), .S (n_530), .A (n_518), .B (n_516), .CI (n_514));
FA_X1 i_264 (.CO (n_529), .S (n_528), .A (n_481), .B (n_479), .CI (n_520));
FA_X1 i_263 (.CO (n_527), .S (n_526), .A (n_467), .B (n_465), .CI (n_463));
FA_X1 i_262 (.CO (n_525), .S (n_524), .A (n_473), .B (n_471), .CI (n_469));
FA_X1 i_261 (.CO (n_523), .S (n_522), .A (n_2856), .B (n_477), .CI (n_475));
FA_X1 i_260 (.CO (n_521), .S (n_520), .A (n_2765), .B (n_2796), .CI (n_2827));
FA_X1 i_259 (.CO (n_519), .S (n_518), .A (n_2672), .B (n_2703), .CI (n_2734));
FA_X1 i_258 (.CO (n_517), .S (n_516), .A (n_2579), .B (n_2610), .CI (n_2641));
FA_X1 i_257 (.CO (n_515), .S (n_514), .A (n_2486), .B (n_2517), .CI (n_2548));
FA_X1 i_256 (.CO (n_513), .S (n_512), .A (n_2393), .B (n_2424), .CI (n_2455));
FA_X1 i_255 (.CO (n_511), .S (n_510), .A (n_2300), .B (n_2331), .CI (n_2362));
FA_X1 i_254 (.CO (n_509), .S (n_508), .A (n_2207), .B (n_2238), .CI (n_2269));
FA_X1 i_253 (.CO (n_507), .S (n_506), .A (n_2114), .B (n_2145), .CI (n_2176));
HA_X1 i_252 (.CO (n_505), .S (n_504), .A (n_459), .B (n_502));
FA_X1 i_251 (.CO (n_503), .S (n_502), .A (n_498), .B (n_457), .CI (n_500));
FA_X1 i_250 (.CO (n_501), .S (n_500), .A (n_494), .B (n_455), .CI (n_496));
FA_X1 i_249 (.CO (n_499), .S (n_498), .A (n_492), .B (n_490), .CI (n_453));
FA_X1 i_248 (.CO (n_497), .S (n_496), .A (n_486), .B (n_484), .CI (n_451));
FA_X1 i_247 (.CO (n_495), .S (n_494), .A (n_449), .B (n_447), .CI (n_488));
FA_X1 i_246 (.CO (n_493), .S (n_492), .A (n_443), .B (n_441), .CI (n_482));
FA_X1 i_245 (.CO (n_491), .S (n_490), .A (n_480), .B (n_478), .CI (n_445));
FA_X1 i_244 (.CO (n_489), .S (n_488), .A (n_466), .B (n_464), .CI (n_462));
FA_X1 i_243 (.CO (n_487), .S (n_486), .A (n_472), .B (n_470), .CI (n_468));
FA_X1 i_242 (.CO (n_485), .S (n_484), .A (n_435), .B (n_476), .CI (n_474));
FA_X1 i_241 (.CO (n_483), .S (n_482), .A (n_421), .B (n_439), .CI (n_437));
FA_X1 i_240 (.CO (n_481), .S (n_480), .A (n_427), .B (n_425), .CI (n_423));
FA_X1 i_239 (.CO (n_479), .S (n_478), .A (n_433), .B (n_431), .CI (n_429));
FA_X1 i_238 (.CO (n_477), .S (n_476), .A (n_2797), .B (n_2828), .CI (n_2857));
FA_X1 i_237 (.CO (n_475), .S (n_474), .A (n_2704), .B (n_2735), .CI (n_2766));
FA_X1 i_236 (.CO (n_473), .S (n_472), .A (n_2611), .B (n_2642), .CI (n_2673));
FA_X1 i_235 (.CO (n_471), .S (n_470), .A (n_2518), .B (n_2549), .CI (n_2580));
FA_X1 i_234 (.CO (n_469), .S (n_468), .A (n_2425), .B (n_2456), .CI (n_2487));
FA_X1 i_233 (.CO (n_467), .S (n_466), .A (n_2332), .B (n_2363), .CI (n_2394));
FA_X1 i_232 (.CO (n_465), .S (n_464), .A (n_2239), .B (n_2270), .CI (n_2301));
FA_X1 i_231 (.CO (n_463), .S (n_462), .A (n_2146), .B (n_2177), .CI (n_2208));
HA_X1 i_230 (.CO (n_461), .S (n_460), .A (n_417), .B (n_458));
FA_X1 i_229 (.CO (n_459), .S (n_458), .A (n_454), .B (n_415), .CI (n_456));
FA_X1 i_228 (.CO (n_457), .S (n_456), .A (n_450), .B (n_413), .CI (n_452));
FA_X1 i_227 (.CO (n_455), .S (n_454), .A (n_409), .B (n_448), .CI (n_411));
FA_X1 i_226 (.CO (n_453), .S (n_452), .A (n_444), .B (n_442), .CI (n_446));
FA_X1 i_225 (.CO (n_451), .S (n_450), .A (n_440), .B (n_407), .CI (n_405));
FA_X1 i_224 (.CO (n_449), .S (n_448), .A (n_436), .B (n_403), .CI (n_401));
FA_X1 i_223 (.CO (n_447), .S (n_446), .A (n_420), .B (n_399), .CI (n_438));
FA_X1 i_222 (.CO (n_445), .S (n_444), .A (n_426), .B (n_424), .CI (n_422));
FA_X1 i_221 (.CO (n_443), .S (n_442), .A (n_432), .B (n_430), .CI (n_428));
FA_X1 i_220 (.CO (n_441), .S (n_440), .A (n_397), .B (n_395), .CI (n_434));
FA_X1 i_219 (.CO (n_439), .S (n_438), .A (n_385), .B (n_383), .CI (n_381));
FA_X1 i_218 (.CO (n_437), .S (n_436), .A (n_391), .B (n_389), .CI (n_387));
FA_X1 i_217 (.CO (n_435), .S (n_434), .A (n_2829), .B (n_2858), .CI (n_393));
FA_X1 i_216 (.CO (n_433), .S (n_432), .A (n_2736), .B (n_2767), .CI (n_2798));
FA_X1 i_215 (.CO (n_431), .S (n_430), .A (n_2643), .B (n_2674), .CI (n_2705));
FA_X1 i_214 (.CO (n_429), .S (n_428), .A (n_2550), .B (n_2581), .CI (n_2612));
FA_X1 i_213 (.CO (n_427), .S (n_426), .A (n_2457), .B (n_2488), .CI (n_2519));
FA_X1 i_212 (.CO (n_425), .S (n_424), .A (n_2364), .B (n_2395), .CI (n_2426));
FA_X1 i_211 (.CO (n_423), .S (n_422), .A (n_2271), .B (n_2302), .CI (n_2333));
FA_X1 i_210 (.CO (n_421), .S (n_420), .A (n_2178), .B (n_2209), .CI (n_2240));
HA_X1 i_209 (.CO (n_419), .S (n_418), .A (n_377), .B (n_416));
FA_X1 i_208 (.CO (n_417), .S (n_416), .A (n_375), .B (n_412), .CI (n_414));
FA_X1 i_207 (.CO (n_415), .S (n_414), .A (n_371), .B (n_373), .CI (n_410));
FA_X1 i_206 (.CO (n_413), .S (n_412), .A (n_369), .B (n_408), .CI (n_406));
FA_X1 i_205 (.CO (n_411), .S (n_410), .A (n_404), .B (n_402), .CI (n_400));
FA_X1 i_204 (.CO (n_409), .S (n_408), .A (n_363), .B (n_361), .CI (n_367));
FA_X1 i_203 (.CO (n_407), .S (n_406), .A (n_396), .B (n_394), .CI (n_365));
FA_X1 i_202 (.CO (n_405), .S (n_404), .A (n_382), .B (n_380), .CI (n_398));
FA_X1 i_201 (.CO (n_403), .S (n_402), .A (n_388), .B (n_386), .CI (n_384));
FA_X1 i_200 (.CO (n_401), .S (n_400), .A (n_357), .B (n_392), .CI (n_390));
FA_X1 i_199 (.CO (n_399), .S (n_398), .A (n_345), .B (n_343), .CI (n_359));
FA_X1 i_198 (.CO (n_397), .S (n_396), .A (n_351), .B (n_349), .CI (n_347));
FA_X1 i_197 (.CO (n_395), .S (n_394), .A (n_2859), .B (n_355), .CI (n_353));
FA_X1 i_196 (.CO (n_393), .S (n_392), .A (n_2768), .B (n_2799), .CI (n_2830));
FA_X1 i_195 (.CO (n_391), .S (n_390), .A (n_2675), .B (n_2706), .CI (n_2737));
FA_X1 i_194 (.CO (n_389), .S (n_388), .A (n_2582), .B (n_2613), .CI (n_2644));
FA_X1 i_193 (.CO (n_387), .S (n_386), .A (n_2489), .B (n_2520), .CI (n_2551));
FA_X1 i_192 (.CO (n_385), .S (n_384), .A (n_2396), .B (n_2427), .CI (n_2458));
FA_X1 i_191 (.CO (n_383), .S (n_382), .A (n_2303), .B (n_2334), .CI (n_2365));
FA_X1 i_190 (.CO (n_381), .S (n_380), .A (n_2210), .B (n_2241), .CI (n_2272));
HA_X1 i_189 (.CO (n_379), .S (n_378), .A (n_339), .B (n_341));
FA_X1 i_188 (.CO (n_377), .S (n_376), .A (n_337), .B (n_372), .CI (n_374));
FA_X1 i_187 (.CO (n_375), .S (n_374), .A (n_333), .B (n_335), .CI (n_370));
FA_X1 i_186 (.CO (n_373), .S (n_372), .A (n_362), .B (n_368), .CI (n_366));
FA_X1 i_185 (.CO (n_371), .S (n_370), .A (n_331), .B (n_329), .CI (n_364));
FA_X1 i_184 (.CO (n_369), .S (n_368), .A (n_327), .B (n_325), .CI (n_360));
FA_X1 i_183 (.CO (n_367), .S (n_366), .A (n_323), .B (n_358), .CI (n_356));
FA_X1 i_182 (.CO (n_365), .S (n_364), .A (n_346), .B (n_344), .CI (n_342));
FA_X1 i_181 (.CO (n_363), .S (n_362), .A (n_352), .B (n_350), .CI (n_348));
FA_X1 i_180 (.CO (n_361), .S (n_360), .A (n_321), .B (n_319), .CI (n_354));
FA_X1 i_179 (.CO (n_359), .S (n_358), .A (n_311), .B (n_309), .CI (n_307));
FA_X1 i_178 (.CO (n_357), .S (n_356), .A (n_317), .B (n_315), .CI (n_313));
FA_X1 i_177 (.CO (n_355), .S (n_354), .A (n_2800), .B (n_2831), .CI (n_2860));
FA_X1 i_176 (.CO (n_353), .S (n_352), .A (n_2707), .B (n_2738), .CI (n_2769));
FA_X1 i_175 (.CO (n_351), .S (n_350), .A (n_2614), .B (n_2645), .CI (n_2676));
FA_X1 i_174 (.CO (n_349), .S (n_348), .A (n_2521), .B (n_2552), .CI (n_2583));
FA_X1 i_173 (.CO (n_347), .S (n_346), .A (n_2428), .B (n_2459), .CI (n_2490));
FA_X1 i_172 (.CO (n_345), .S (n_344), .A (n_2335), .B (n_2366), .CI (n_2397));
FA_X1 i_171 (.CO (n_343), .S (n_342), .A (n_2242), .B (n_2273), .CI (n_2304));
HA_X1 i_170 (.CO (n_341), .S (n_340), .A (n_303), .B (n_338));
FA_X1 i_169 (.CO (n_339), .S (n_338), .A (n_334), .B (n_301), .CI (n_336));
FA_X1 i_168 (.CO (n_337), .S (n_336), .A (n_330), .B (n_299), .CI (n_332));
FA_X1 i_167 (.CO (n_335), .S (n_334), .A (n_326), .B (n_324), .CI (n_297));
FA_X1 i_166 (.CO (n_333), .S (n_332), .A (n_293), .B (n_295), .CI (n_328));
FA_X1 i_165 (.CO (n_331), .S (n_330), .A (n_320), .B (n_291), .CI (n_289));
FA_X1 i_164 (.CO (n_329), .S (n_328), .A (n_308), .B (n_306), .CI (n_322));
FA_X1 i_163 (.CO (n_327), .S (n_326), .A (n_314), .B (n_312), .CI (n_310));
FA_X1 i_162 (.CO (n_325), .S (n_324), .A (n_285), .B (n_318), .CI (n_316));
FA_X1 i_161 (.CO (n_323), .S (n_322), .A (n_275), .B (n_273), .CI (n_287));
FA_X1 i_160 (.CO (n_321), .S (n_320), .A (n_281), .B (n_279), .CI (n_277));
FA_X1 i_159 (.CO (n_319), .S (n_318), .A (n_2832), .B (n_2861), .CI (n_283));
FA_X1 i_158 (.CO (n_317), .S (n_316), .A (n_2739), .B (n_2770), .CI (n_2801));
FA_X1 i_157 (.CO (n_315), .S (n_314), .A (n_2646), .B (n_2677), .CI (n_2708));
FA_X1 i_156 (.CO (n_313), .S (n_312), .A (n_2553), .B (n_2584), .CI (n_2615));
FA_X1 i_155 (.CO (n_311), .S (n_310), .A (n_2460), .B (n_2491), .CI (n_2522));
FA_X1 i_154 (.CO (n_309), .S (n_308), .A (n_2367), .B (n_2398), .CI (n_2429));
FA_X1 i_153 (.CO (n_307), .S (n_306), .A (n_2274), .B (n_2305), .CI (n_2336));
HA_X1 i_152 (.CO (n_305), .S (n_304), .A (n_269), .B (n_302));
FA_X1 i_151 (.CO (n_303), .S (n_302), .A (n_267), .B (n_298), .CI (n_300));
FA_X1 i_150 (.CO (n_301), .S (n_300), .A (n_294), .B (n_265), .CI (n_296));
FA_X1 i_149 (.CO (n_299), .S (n_298), .A (n_261), .B (n_292), .CI (n_290));
FA_X1 i_148 (.CO (n_297), .S (n_296), .A (n_257), .B (n_288), .CI (n_263));
FA_X1 i_147 (.CO (n_295), .S (n_294), .A (n_286), .B (n_284), .CI (n_259));
FA_X1 i_146 (.CO (n_293), .S (n_292), .A (n_274), .B (n_272), .CI (n_255));
FA_X1 i_145 (.CO (n_291), .S (n_290), .A (n_280), .B (n_278), .CI (n_276));
FA_X1 i_144 (.CO (n_289), .S (n_288), .A (n_241), .B (n_253), .CI (n_282));
FA_X1 i_143 (.CO (n_287), .S (n_286), .A (n_247), .B (n_245), .CI (n_243));
FA_X1 i_142 (.CO (n_285), .S (n_284), .A (n_2862), .B (n_251), .CI (n_249));
FA_X1 i_141 (.CO (n_283), .S (n_282), .A (n_2771), .B (n_2802), .CI (n_2833));
FA_X1 i_140 (.CO (n_281), .S (n_280), .A (n_2678), .B (n_2709), .CI (n_2740));
FA_X1 i_139 (.CO (n_279), .S (n_278), .A (n_2585), .B (n_2616), .CI (n_2647));
FA_X1 i_138 (.CO (n_277), .S (n_276), .A (n_2492), .B (n_2523), .CI (n_2554));
FA_X1 i_137 (.CO (n_275), .S (n_274), .A (n_2399), .B (n_2430), .CI (n_2461));
FA_X1 i_136 (.CO (n_273), .S (n_272), .A (n_2306), .B (n_2337), .CI (n_2368));
HA_X1 i_135 (.CO (n_271), .S (n_270), .A (n_237), .B (n_239));
FA_X1 i_134 (.CO (n_269), .S (n_268), .A (n_235), .B (n_264), .CI (n_266));
FA_X1 i_133 (.CO (n_267), .S (n_266), .A (n_260), .B (n_262), .CI (n_233));
FA_X1 i_132 (.CO (n_265), .S (n_264), .A (n_231), .B (n_258), .CI (n_256));
FA_X1 i_131 (.CO (n_263), .S (n_262), .A (n_252), .B (n_229), .CI (n_227));
FA_X1 i_130 (.CO (n_261), .S (n_260), .A (n_240), .B (n_225), .CI (n_254));
FA_X1 i_129 (.CO (n_259), .S (n_258), .A (n_246), .B (n_244), .CI (n_242));
FA_X1 i_128 (.CO (n_257), .S (n_256), .A (n_221), .B (n_250), .CI (n_248));
FA_X1 i_127 (.CO (n_255), .S (n_254), .A (n_213), .B (n_211), .CI (n_223));
FA_X1 i_126 (.CO (n_253), .S (n_252), .A (n_219), .B (n_217), .CI (n_215));
FA_X1 i_125 (.CO (n_251), .S (n_250), .A (n_2803), .B (n_2834), .CI (n_2863));
FA_X1 i_124 (.CO (n_249), .S (n_248), .A (n_2710), .B (n_2741), .CI (n_2772));
FA_X1 i_123 (.CO (n_247), .S (n_246), .A (n_2617), .B (n_2648), .CI (n_2679));
FA_X1 i_122 (.CO (n_245), .S (n_244), .A (n_2524), .B (n_2555), .CI (n_2586));
FA_X1 i_121 (.CO (n_243), .S (n_242), .A (n_2431), .B (n_2462), .CI (n_2493));
FA_X1 i_120 (.CO (n_241), .S (n_240), .A (n_2338), .B (n_2369), .CI (n_2400));
HA_X1 i_119 (.CO (n_239), .S (n_238), .A (n_207), .B (n_209));
FA_X1 i_118 (.CO (n_237), .S (n_236), .A (n_232), .B (n_205), .CI (n_234));
FA_X1 i_117 (.CO (n_235), .S (n_234), .A (n_226), .B (n_230), .CI (n_203));
FA_X1 i_116 (.CO (n_233), .S (n_232), .A (n_224), .B (n_201), .CI (n_228));
FA_X1 i_115 (.CO (n_231), .S (n_230), .A (n_222), .B (n_199), .CI (n_197));
FA_X1 i_114 (.CO (n_229), .S (n_228), .A (n_214), .B (n_212), .CI (n_210));
FA_X1 i_113 (.CO (n_227), .S (n_226), .A (n_220), .B (n_218), .CI (n_216));
FA_X1 i_112 (.CO (n_225), .S (n_224), .A (n_183), .B (n_195), .CI (n_193));
FA_X1 i_111 (.CO (n_223), .S (n_222), .A (n_189), .B (n_187), .CI (n_185));
FA_X1 i_110 (.CO (n_221), .S (n_220), .A (n_2835), .B (n_2864), .CI (n_191));
FA_X1 i_109 (.CO (n_219), .S (n_218), .A (n_2742), .B (n_2773), .CI (n_2804));
FA_X1 i_108 (.CO (n_217), .S (n_216), .A (n_2649), .B (n_2680), .CI (n_2711));
FA_X1 i_107 (.CO (n_215), .S (n_214), .A (n_2556), .B (n_2587), .CI (n_2618));
FA_X1 i_106 (.CO (n_213), .S (n_212), .A (n_2463), .B (n_2494), .CI (n_2525));
FA_X1 i_105 (.CO (n_211), .S (n_210), .A (n_2370), .B (n_2401), .CI (n_2432));
HA_X1 i_104 (.CO (n_209), .S (n_208), .A (n_179), .B (n_181));
FA_X1 i_103 (.CO (n_207), .S (n_206), .A (n_177), .B (n_202), .CI (n_204));
FA_X1 i_102 (.CO (n_205), .S (n_204), .A (n_196), .B (n_175), .CI (n_200));
FA_X1 i_101 (.CO (n_203), .S (n_202), .A (n_171), .B (n_173), .CI (n_198));
FA_X1 i_100 (.CO (n_201), .S (n_200), .A (n_169), .B (n_194), .CI (n_192));
FA_X1 i_99 (.CO (n_199), .S (n_198), .A (n_186), .B (n_184), .CI (n_182));
FA_X1 i_98 (.CO (n_197), .S (n_196), .A (n_167), .B (n_190), .CI (n_188));
FA_X1 i_97 (.CO (n_195), .S (n_194), .A (n_161), .B (n_159), .CI (n_157));
FA_X1 i_96 (.CO (n_193), .S (n_192), .A (n_2865), .B (n_165), .CI (n_163));
FA_X1 i_95 (.CO (n_191), .S (n_190), .A (n_2774), .B (n_2805), .CI (n_2836));
FA_X1 i_94 (.CO (n_189), .S (n_188), .A (n_2681), .B (n_2712), .CI (n_2743));
FA_X1 i_93 (.CO (n_187), .S (n_186), .A (n_2588), .B (n_2619), .CI (n_2650));
FA_X1 i_92 (.CO (n_185), .S (n_184), .A (n_2495), .B (n_2526), .CI (n_2557));
FA_X1 i_91 (.CO (n_183), .S (n_182), .A (n_2402), .B (n_2433), .CI (n_2464));
HA_X1 i_90 (.CO (n_181), .S (n_180), .A (n_153), .B (n_155));
FA_X1 i_89 (.CO (n_179), .S (n_178), .A (n_174), .B (n_151), .CI (n_176));
FA_X1 i_88 (.CO (n_177), .S (n_176), .A (n_149), .B (n_172), .CI (n_170));
FA_X1 i_87 (.CO (n_175), .S (n_174), .A (n_147), .B (n_145), .CI (n_168));
FA_X1 i_86 (.CO (n_173), .S (n_172), .A (n_158), .B (n_156), .CI (n_166));
FA_X1 i_85 (.CO (n_171), .S (n_170), .A (n_164), .B (n_162), .CI (n_160));
FA_X1 i_84 (.CO (n_169), .S (n_168), .A (n_133), .B (n_143), .CI (n_141));
FA_X1 i_83 (.CO (n_167), .S (n_166), .A (n_139), .B (n_137), .CI (n_135));
FA_X1 i_82 (.CO (n_165), .S (n_164), .A (n_2806), .B (n_2837), .CI (n_2866));
FA_X1 i_81 (.CO (n_163), .S (n_162), .A (n_2713), .B (n_2744), .CI (n_2775));
FA_X1 i_80 (.CO (n_161), .S (n_160), .A (n_2620), .B (n_2651), .CI (n_2682));
FA_X1 i_79 (.CO (n_159), .S (n_158), .A (n_2527), .B (n_2558), .CI (n_2589));
FA_X1 i_78 (.CO (n_157), .S (n_156), .A (n_2434), .B (n_2465), .CI (n_2496));
HA_X1 i_77 (.CO (n_155), .S (n_154), .A (n_150), .B (n_131));
FA_X1 i_76 (.CO (n_153), .S (n_152), .A (n_148), .B (n_127), .CI (n_129));
FA_X1 i_75 (.CO (n_151), .S (n_150), .A (n_125), .B (n_146), .CI (n_144));
FA_X1 i_74 (.CO (n_149), .S (n_148), .A (n_121), .B (n_142), .CI (n_123));
FA_X1 i_73 (.CO (n_147), .S (n_146), .A (n_136), .B (n_134), .CI (n_132));
FA_X1 i_72 (.CO (n_145), .S (n_144), .A (n_119), .B (n_140), .CI (n_138));
FA_X1 i_71 (.CO (n_143), .S (n_142), .A (n_115), .B (n_113), .CI (n_111));
FA_X1 i_70 (.CO (n_141), .S (n_140), .A (n_2838), .B (n_2867), .CI (n_117));
FA_X1 i_69 (.CO (n_139), .S (n_138), .A (n_2745), .B (n_2776), .CI (n_2807));
FA_X1 i_68 (.CO (n_137), .S (n_136), .A (n_2652), .B (n_2683), .CI (n_2714));
FA_X1 i_67 (.CO (n_135), .S (n_134), .A (n_2559), .B (n_2590), .CI (n_2621));
FA_X1 i_66 (.CO (n_133), .S (n_132), .A (n_2466), .B (n_2497), .CI (n_2528));
HA_X1 i_65 (.CO (n_131), .S (n_130), .A (n_107), .B (n_109));
FA_X1 i_64 (.CO (n_129), .S (n_128), .A (n_105), .B (n_124), .CI (n_126));
FA_X1 i_63 (.CO (n_127), .S (n_126), .A (n_101), .B (n_103), .CI (n_122));
FA_X1 i_62 (.CO (n_125), .S (n_124), .A (n_110), .B (n_120), .CI (n_118));
FA_X1 i_61 (.CO (n_123), .S (n_122), .A (n_116), .B (n_114), .CI (n_112));
FA_X1 i_60 (.CO (n_121), .S (n_120), .A (n_93), .B (n_91), .CI (n_99));
FA_X1 i_59 (.CO (n_119), .S (n_118), .A (n_2868), .B (n_97), .CI (n_95));
FA_X1 i_58 (.CO (n_117), .S (n_116), .A (n_2777), .B (n_2808), .CI (n_2839));
FA_X1 i_57 (.CO (n_115), .S (n_114), .A (n_2684), .B (n_2715), .CI (n_2746));
FA_X1 i_56 (.CO (n_113), .S (n_112), .A (n_2591), .B (n_2622), .CI (n_2653));
FA_X1 i_55 (.CO (n_111), .S (n_110), .A (n_2498), .B (n_2529), .CI (n_2560));
HA_X1 i_54 (.CO (n_109), .S (n_108), .A (n_89), .B (n_87));
FA_X1 i_53 (.CO (n_107), .S (n_106), .A (n_102), .B (n_100), .CI (n_104));
FA_X1 i_52 (.CO (n_105), .S (n_104), .A (n_98), .B (n_83), .CI (n_85));
FA_X1 i_51 (.CO (n_103), .S (n_102), .A (n_92), .B (n_90), .CI (n_81));
FA_X1 i_50 (.CO (n_101), .S (n_100), .A (n_79), .B (n_96), .CI (n_94));
FA_X1 i_49 (.CO (n_99), .S (n_98), .A (n_77), .B (n_75), .CI (n_73));
FA_X1 i_48 (.CO (n_97), .S (n_96), .A (n_2809), .B (n_2840), .CI (n_2869));
FA_X1 i_47 (.CO (n_95), .S (n_94), .A (n_2716), .B (n_2747), .CI (n_2778));
FA_X1 i_46 (.CO (n_93), .S (n_92), .A (n_2623), .B (n_2654), .CI (n_2685));
FA_X1 i_45 (.CO (n_91), .S (n_90), .A (n_2530), .B (n_2561), .CI (n_2592));
HA_X1 i_44 (.CO (n_89), .S (n_88), .A (n_71), .B (n_69));
FA_X1 i_43 (.CO (n_87), .S (n_86), .A (n_67), .B (n_82), .CI (n_84));
FA_X1 i_42 (.CO (n_85), .S (n_84), .A (n_72), .B (n_80), .CI (n_65));
FA_X1 i_41 (.CO (n_83), .S (n_82), .A (n_78), .B (n_76), .CI (n_74));
FA_X1 i_40 (.CO (n_81), .S (n_80), .A (n_59), .B (n_57), .CI (n_63));
FA_X1 i_39 (.CO (n_79), .S (n_78), .A (n_2841), .B (n_2870), .CI (n_61));
FA_X1 i_38 (.CO (n_77), .S (n_76), .A (n_2748), .B (n_2779), .CI (n_2810));
FA_X1 i_37 (.CO (n_75), .S (n_74), .A (n_2655), .B (n_2686), .CI (n_2717));
FA_X1 i_36 (.CO (n_73), .S (n_72), .A (n_2562), .B (n_2593), .CI (n_2624));
HA_X1 i_35 (.CO (n_71), .S (n_70), .A (n_55), .B (n_53));
FA_X1 i_34 (.CO (n_69), .S (n_68), .A (n_51), .B (n_64), .CI (n_66));
FA_X1 i_33 (.CO (n_67), .S (n_66), .A (n_56), .B (n_49), .CI (n_62));
FA_X1 i_32 (.CO (n_65), .S (n_64), .A (n_43), .B (n_60), .CI (n_58));
FA_X1 i_31 (.CO (n_63), .S (n_62), .A (n_2871), .B (n_47), .CI (n_45));
FA_X1 i_30 (.CO (n_61), .S (n_60), .A (n_2780), .B (n_2811), .CI (n_2842));
FA_X1 i_29 (.CO (n_59), .S (n_58), .A (n_2687), .B (n_2718), .CI (n_2749));
FA_X1 i_28 (.CO (n_57), .S (n_56), .A (n_2594), .B (n_2625), .CI (n_2656));
HA_X1 i_27 (.CO (n_55), .S (n_54), .A (n_39), .B (n_50));
FA_X1 i_26 (.CO (n_53), .S (n_52), .A (n_48), .B (n_37), .CI (n_41));
FA_X1 i_25 (.CO (n_51), .S (n_50), .A (n_46), .B (n_44), .CI (n_42));
FA_X1 i_24 (.CO (n_49), .S (n_48), .A (n_33), .B (n_31), .CI (n_35));
FA_X1 i_23 (.CO (n_47), .S (n_46), .A (n_2812), .B (n_2843), .CI (n_2872));
FA_X1 i_22 (.CO (n_45), .S (n_44), .A (n_2719), .B (n_2750), .CI (n_2781));
FA_X1 i_21 (.CO (n_43), .S (n_42), .A (n_2626), .B (n_2657), .CI (n_2688));
HA_X1 i_20 (.CO (n_41), .S (n_40), .A (n_36), .B (n_27));
FA_X1 i_19 (.CO (n_39), .S (n_38), .A (n_32), .B (n_30), .CI (n_29));
FA_X1 i_18 (.CO (n_37), .S (n_36), .A (n_21), .B (n_25), .CI (n_34));
FA_X1 i_17 (.CO (n_35), .S (n_34), .A (n_2844), .B (n_2873), .CI (n_23));
FA_X1 i_16 (.CO (n_33), .S (n_32), .A (n_2751), .B (n_2782), .CI (n_2813));
FA_X1 i_15 (.CO (n_31), .S (n_30), .A (n_2658), .B (n_2689), .CI (n_2720));
HA_X1 i_14 (.CO (n_29), .S (n_28), .A (n_19), .B (n_17));
FA_X1 i_13 (.CO (n_27), .S (n_26), .A (n_22), .B (n_20), .CI (n_24));
FA_X1 i_12 (.CO (n_25), .S (n_24), .A (n_2874), .B (n_15), .CI (n_13));
FA_X1 i_11 (.CO (n_23), .S (n_22), .A (n_2783), .B (n_2814), .CI (n_2845));
FA_X1 i_10 (.CO (n_21), .S (n_20), .A (n_2690), .B (n_2721), .CI (n_2752));
HA_X1 i_9 (.CO (n_19), .S (n_18), .A (n_12), .B (n_11));
FA_X1 i_8 (.CO (n_17), .S (n_16), .A (n_7), .B (n_9), .CI (n_14));
FA_X1 i_7 (.CO (n_15), .S (n_14), .A (n_2815), .B (n_2846), .CI (n_2875));
FA_X1 i_6 (.CO (n_13), .S (n_12), .A (n_2722), .B (n_2753), .CI (n_2784));
HA_X1 i_5 (.CO (n_11), .S (n_10), .A (n_3), .B (n_8));
FA_X1 i_4 (.CO (n_9), .S (n_8), .A (n_2847), .B (n_2876), .CI (n_5));
FA_X1 i_3 (.CO (n_7), .S (n_6), .A (n_2754), .B (n_2785), .CI (n_2816));
HA_X1 i_2 (.CO (n_5), .S (n_4), .A (n_2877), .B (n_1));
FA_X1 i_1 (.CO (n_3), .S (n_2), .A (n_2786), .B (n_2817), .CI (n_2848));
HA_X1 i_0 (.CO (n_1), .S (n_0), .A (n_2818), .B (n_3231));
CLKBUF_X2 sgo__L1_c3 (.Z (sgo__n3), .A (n_3298));
CLKBUF_X1 sgo__L1_c5 (.Z (sgo__n5), .A (n_3298));
BUF_X8 sgo__L1_c208 (.Z (sgo__n208), .A (n_3118));
CLKBUF_X1 sgo__L1_c10 (.Z (sgo__n10), .A (n_3249));
CLKBUF_X3 sgo__L1_c19 (.Z (sgo__n19), .A (n_3301));
OR2_X1 sgo__sro_c219 (.ZN (sgo__sro_n217), .A1 (n_3165), .A2 (n_3132));
OAI221_X1 sgo__sro_c220 (.ZN (sgo__sro_n216), .A (sgo__sro_n217), .B1 (n_3155), .B2 (n_3120)
    , .C1 (n_3154), .C2 (n_3138));
INV_X1 sgo__sro_c230 (.ZN (sgo__sro_n227), .A (n_3044));
NOR2_X1 sgo__sro_c231 (.ZN (sgo__sro_n226), .A1 (n_3040), .A2 (n_3043));
NAND2_X1 sgo__sro_c232 (.ZN (sgo__sro_n225), .A1 (sgo__sro_n227), .A2 (sgo__sro_n226));
NOR2_X2 sgo__sro_c233 (.ZN (sgo__sro_n224), .A1 (n_3047), .A2 (sgo__sro_n225));
CLKBUF_X1 sgo__L1_c43 (.Z (sgo__n43), .A (n_3297));
CLKBUF_X1 sgo__L1_c78 (.Z (sgo__n78), .A (n_3295));
CLKBUF_X1 sgo__L1_c98 (.Z (sgo__n98), .A (n_3296));
CLKBUF_X2 sgo__L1_c99 (.Z (sgo__n99), .A (n_3267));
CLKBUF_X3 sgo__L1_c109 (.Z (sgo__n109), .A (n_3304));
CLKBUF_X2 sgo__L1_c122 (.Z (sgo__n122), .A (n_3265));
CLKBUF_X1 CLOCK_sgo__L1_c364 (.Z (CLOCK_sgo__n358), .A (n_3306));
CLKBUF_X1 sgo__L1_c134 (.Z (sgo__n134), .A (n_3257));
CLKBUF_X1 sgo__L1_c141 (.Z (sgo__n141), .A (n_3289));
CLKBUF_X2 sgo__L1_c147 (.Z (sgo__n147), .A (n_3261));
CLKBUF_X1 sgo__L1_c148 (.Z (sgo__n148), .A (n_3261));
CLKBUF_X1 sgo__L1_c150 (.Z (sgo__n150), .A (n_3261));
CLKBUF_X1 sgo__L2_c162 (.Z (sgo__n162), .A (n_3263));
CLKBUF_X1 sgo__L1_c164 (.Z (sgo__n164), .A (n_3286));
CLKBUF_X1 sgo__L1_c168 (.Z (sgo__n168), .A (n_3269));
CLKBUF_X1 sgo__L1_c170 (.Z (sgo__n170), .A (n_3268));
CLKBUF_X2 sgo__L1_c172 (.Z (sgo__n172), .A (n_3268));
CLKBUF_X1 sgo__L1_c174 (.Z (sgo__n174), .A (n_3259));
CLKBUF_X3 CLOCK_sgo__L1_c365 (.Z (CLOCK_sgo__n359), .A (n_3306));
CLKBUF_X2 sgo__L1_c176 (.Z (sgo__n176), .A (n_3262));
CLKBUF_X1 sgo__L1_c177 (.Z (sgo__n177), .A (n_3255));
BUF_X1 sgo__L1_c178 (.Z (sgo__n178), .A (n_3255));
CLKBUF_X1 sgo__L1_c180 (.Z (sgo__n180), .A (n_3255));
BUF_X1 sgo__L1_c182 (.Z (sgo__n182), .A (n_3256));
BUF_X4 CLOCK_opt_ipo_c363 (.Z (CLOCK_opt_ipo_n357), .A (n_3054));
CLKBUF_X1 sgo__L1_c195 (.Z (sgo__n195), .A (n_3264));
CLKBUF_X1 sgo__L1_c201 (.Z (sgo__n201), .A (n_3260));
CLKBUF_X1 sgo__L1_c203 (.Z (sgo__n203), .A (n_3270));

endmodule //datapath

module multOperator (clk_CTS_0_PP_0, clk_CTS_0_PP_9, clk_CTS_0_PP_10, clk, rst, a, 
    b, c);

output [63:0] c;
output clk_CTS_0_PP_0;
output clk_CTS_0_PP_9;
input [31:0] a;
input [31:0] b;
input clk;
input rst;
input clk_CTS_0_PP_10;
wire n_64;
wire n_0;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire hfn_ipo_n5;
wire hfn_ipo_n6;
wire CTS_n_tid0_18;
wire CTS_n_tid0_60;


datapath i_1 (.p_0 ({n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
    n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
    n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, 
    n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, 
    n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1})
    , .a ({a[31], a[30], a[29], a[28], a[27], a[26], a[25], a[24], a[23], a[22], 
    a[21], a[20], a[19], a[18], a[17], a[16], a[15], a[14], a[13], a[12], a[11], 
    a[10], a[9], a[8], a[7], a[6], a[5], a[4], a[3], a[2], a[1], a[0]}), .b ({b[31], 
    b[30], b[29], b[28], b[27], b[26], b[25], b[24], b[23], b[22], b[21], b[20], 
    b[19], b[18], b[17], b[16], b[15], b[14], b[13], b[12], b[11], b[10], b[9], b[8], 
    b[7], b[6], b[5], b[4], b[3], b[2], b[1], b[0]}));
DFFR_X1 \c_reg[0]  (.Q (c[0]), .CK (CTS_n_tid0_60), .D (n_1), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[1]  (.Q (c[1]), .CK (CTS_n_tid0_60), .D (n_2), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[2]  (.Q (c[2]), .CK (CTS_n_tid0_60), .D (n_3), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[3]  (.Q (c[3]), .CK (CTS_n_tid0_60), .D (n_4), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[4]  (.Q (c[4]), .CK (CTS_n_tid0_60), .D (n_5), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[5]  (.Q (c[5]), .CK (CTS_n_tid0_60), .D (n_6), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[6]  (.Q (c[6]), .CK (CTS_n_tid0_60), .D (n_7), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[7]  (.Q (c[7]), .CK (CTS_n_tid0_60), .D (n_8), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[8]  (.Q (c[8]), .CK (CTS_n_tid0_60), .D (n_9), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[9]  (.Q (c[9]), .CK (CTS_n_tid0_60), .D (n_10), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[10]  (.Q (c[10]), .CK (CTS_n_tid0_60), .D (n_11), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[11]  (.Q (c[11]), .CK (CTS_n_tid0_60), .D (n_12), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[12]  (.Q (c[12]), .CK (CTS_n_tid0_60), .D (n_13), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[13]  (.Q (c[13]), .CK (CTS_n_tid0_60), .D (n_14), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[14]  (.Q (c[14]), .CK (CTS_n_tid0_60), .D (n_15), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[15]  (.Q (c[15]), .CK (CTS_n_tid0_60), .D (n_16), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[16]  (.Q (c[16]), .CK (CTS_n_tid0_18), .D (n_17), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[17]  (.Q (c[17]), .CK (CTS_n_tid0_18), .D (n_18), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[18]  (.Q (c[18]), .CK (CTS_n_tid0_18), .D (n_19), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[19]  (.Q (c[19]), .CK (CTS_n_tid0_18), .D (n_20), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[20]  (.Q (c[20]), .CK (CTS_n_tid0_18), .D (n_21), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[21]  (.Q (c[21]), .CK (CTS_n_tid0_18), .D (n_22), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[22]  (.Q (c[22]), .CK (CTS_n_tid0_18), .D (n_23), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[23]  (.Q (c[23]), .CK (CTS_n_tid0_18), .D (n_24), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[24]  (.Q (c[24]), .CK (CTS_n_tid0_18), .D (n_25), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[25]  (.Q (c[25]), .CK (CTS_n_tid0_18), .D (n_26), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[26]  (.Q (c[26]), .CK (CTS_n_tid0_18), .D (n_27), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[27]  (.Q (c[27]), .CK (CTS_n_tid0_18), .D (n_28), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[28]  (.Q (c[28]), .CK (CTS_n_tid0_18), .D (n_29), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[29]  (.Q (c[29]), .CK (CTS_n_tid0_18), .D (n_30), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[30]  (.Q (c[30]), .CK (CTS_n_tid0_18), .D (n_31), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[31]  (.Q (c[31]), .CK (CTS_n_tid0_18), .D (n_32), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[32]  (.Q (c[32]), .CK (CTS_n_tid0_18), .D (n_33), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[33]  (.Q (c[33]), .CK (CTS_n_tid0_60), .D (n_34), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[34]  (.Q (c[34]), .CK (CTS_n_tid0_60), .D (n_35), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[35]  (.Q (c[35]), .CK (CTS_n_tid0_60), .D (n_36), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[36]  (.Q (c[36]), .CK (CTS_n_tid0_60), .D (n_37), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[37]  (.Q (c[37]), .CK (CTS_n_tid0_60), .D (n_38), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[38]  (.Q (c[38]), .CK (CTS_n_tid0_60), .D (n_39), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[39]  (.Q (c[39]), .CK (CTS_n_tid0_60), .D (n_40), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[40]  (.Q (c[40]), .CK (CTS_n_tid0_60), .D (n_41), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[41]  (.Q (c[41]), .CK (CTS_n_tid0_60), .D (n_42), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[42]  (.Q (c[42]), .CK (CTS_n_tid0_60), .D (n_43), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[43]  (.Q (c[43]), .CK (CTS_n_tid0_60), .D (n_44), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[44]  (.Q (c[44]), .CK (CTS_n_tid0_60), .D (n_45), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[45]  (.Q (c[45]), .CK (CTS_n_tid0_60), .D (n_46), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[46]  (.Q (c[46]), .CK (CTS_n_tid0_60), .D (n_47), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[47]  (.Q (c[47]), .CK (CTS_n_tid0_60), .D (n_48), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[48]  (.Q (c[48]), .CK (CTS_n_tid0_60), .D (n_49), .RN (hfn_ipo_n5));
DFFR_X1 \c_reg[49]  (.Q (c[49]), .CK (CTS_n_tid0_18), .D (n_50), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[50]  (.Q (c[50]), .CK (CTS_n_tid0_18), .D (n_51), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[51]  (.Q (c[51]), .CK (CTS_n_tid0_18), .D (n_52), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[52]  (.Q (c[52]), .CK (CTS_n_tid0_18), .D (n_53), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[53]  (.Q (c[53]), .CK (CTS_n_tid0_18), .D (n_54), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[54]  (.Q (c[54]), .CK (CTS_n_tid0_18), .D (n_55), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[55]  (.Q (c[55]), .CK (CTS_n_tid0_18), .D (n_56), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[56]  (.Q (c[56]), .CK (CTS_n_tid0_18), .D (n_57), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[57]  (.Q (c[57]), .CK (CTS_n_tid0_18), .D (n_58), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[58]  (.Q (c[58]), .CK (CTS_n_tid0_18), .D (n_59), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[59]  (.Q (c[59]), .CK (CTS_n_tid0_18), .D (n_60), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[60]  (.Q (c[60]), .CK (CTS_n_tid0_18), .D (n_61), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[61]  (.Q (c[61]), .CK (CTS_n_tid0_60), .D (n_62), .RN (hfn_ipo_n6));
DFFR_X1 \c_reg[62]  (.Q (c[62]), .CK (CTS_n_tid0_60), .D (n_63), .RN (hfn_ipo_n6));
INV_X1 i_0_0 (.ZN (n_0), .A (rst));
DFFR_X1 \c_reg[63]  (.Q (c[63]), .CK (CTS_n_tid0_60), .D (n_64), .RN (hfn_ipo_n6));
BUF_X4 hfn_ipo_c5 (.Z (hfn_ipo_n5), .A (n_0));
CLKBUF_X2 hfn_ipo_c6 (.Z (hfn_ipo_n6), .A (n_0));
CLKBUF_X2 CTS_L3_c_tid0_17 (.Z (CTS_n_tid0_18), .A (clk_CTS_0_PP_0));
CLKBUF_X2 CTS_L2_c_tid0_64 (.Z (clk_CTS_0_PP_0), .A (clk_CTS_0_PP_9));
CLKBUF_X1 CTS_L1_c_tid0_77 (.Z (clk_CTS_0_PP_9), .A (clk_CTS_0_PP_10));
CLKBUF_X3 CTS_L3_c_tid0_59 (.Z (CTS_n_tid0_60), .A (clk_CTS_0_PP_0));

endmodule //multOperator

module buffer (clk_CTS_0_PP_0, clk, rst, en, D, Q);

output [31:0] Q;
input [31:0] D;
input clk;
input en;
input rst;
input clk_CTS_0_PP_0;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_2;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid1_3;
wire CLOCK_slh__n101;
wire CLOCK_slh__n107;
wire CLOCK_slh__n102;
wire CLOCK_slh__n103;
wire CLOCK_slh__n108;
wire CLOCK_slh__n109;
wire CLOCK_slh__n113;
wire CLOCK_slh__n114;
wire CLOCK_slh__n115;
wire CLOCK_slh__n119;
wire CLOCK_slh__n120;
wire CLOCK_slh__n121;
wire CLOCK_slh__n125;
wire CLOCK_slh__n126;
wire CLOCK_slh__n127;
wire CLOCK_slh__n131;
wire CLOCK_slh__n132;
wire CLOCK_slh__n133;
wire CLOCK_slh__n137;
wire CLOCK_slh__n138;
wire CLOCK_slh__n139;
wire CLOCK_slh__n143;
wire CLOCK_slh__n144;
wire CLOCK_slh__n145;
wire CLOCK_slh__n149;
wire CLOCK_slh__n150;
wire CLOCK_slh__n151;
wire CLOCK_slh__n155;
wire CLOCK_slh__n156;
wire CLOCK_slh__n157;
wire CLOCK_slh__n161;
wire CLOCK_slh__n162;
wire CLOCK_slh__n163;
wire CLOCK_slh__n167;
wire CLOCK_slh__n168;
wire CLOCK_slh__n169;
wire CLOCK_slh__n173;
wire CLOCK_slh__n174;
wire CLOCK_slh__n175;
wire CLOCK_slh__n179;
wire CLOCK_slh__n180;
wire CLOCK_slh__n181;
wire CLOCK_slh__n185;
wire CLOCK_slh__n186;
wire CLOCK_slh__n187;
wire CLOCK_slh__n191;
wire CLOCK_slh__n192;
wire CLOCK_slh__n193;
wire CLOCK_slh__n197;
wire CLOCK_slh__n198;
wire CLOCK_slh__n199;
wire CLOCK_slh__n203;
wire CLOCK_slh__n205;
wire CLOCK_slh__n207;
wire CLOCK_slh__n208;
wire CLOCK_slh__n209;
wire CLOCK_slh__n213;
wire CLOCK_slh__n214;
wire CLOCK_slh__n215;
wire CLOCK_slh__n219;
wire CLOCK_slh__n220;
wire CLOCK_slh__n221;
wire CLOCK_slh__n225;
wire CLOCK_slh__n226;
wire CLOCK_slh__n227;
wire CLOCK_slh__n231;
wire CLOCK_slh__n232;
wire CLOCK_slh__n233;
wire CLOCK_slh__n237;
wire CLOCK_slh__n238;
wire CLOCK_slh__n239;
wire CLOCK_slh__n243;
wire CLOCK_slh__n244;
wire CLOCK_slh__n245;
wire CLOCK_slh__n249;
wire CLOCK_slh__n250;
wire CLOCK_slh__n251;
wire CLOCK_slh__n255;
wire CLOCK_slh__n256;
wire CLOCK_slh__n257;
wire CLOCK_slh__n261;
wire CLOCK_slh__n262;
wire CLOCK_slh__n263;
wire CLOCK_slh__n267;
wire CLOCK_slh__n268;
wire CLOCK_slh__n269;
wire CLOCK_slh__n270;
wire CLOCK_slh__n271;
wire CLOCK_slh__n272;
wire CLOCK_slh__n273;
wire CLOCK_slh__n274;
wire CLOCK_slh__n275;
wire CLOCK_slh__n276;
wire CLOCK_slh__n277;
wire CLOCK_slh__n278;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n125), .A1 (n_0_0), .A2 (D[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n161), .A1 (n_0_0), .A2 (D[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n155), .A1 (n_0_0), .A2 (D[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n167), .A1 (n_0_0), .A2 (D[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n173), .A1 (n_0_0), .A2 (D[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n267), .A1 (n_0_0), .A2 (D[26]));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n131), .A1 (n_0_0), .A2 (D[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n119), .A1 (n_0_0), .A2 (D[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n137), .A1 (n_0_0), .A2 (D[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n179), .A1 (n_0_0), .A2 (D[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n197), .A1 (n_0_0), .A2 (CLOCK_slh__n205));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n207), .A1 (n_0_0), .A2 (D[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n191), .A1 (n_0_0), .A2 (CLOCK_slh__n203));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n213), .A1 (n_0_0), .A2 (D[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n225), .A1 (n_0_0), .A2 (D[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n219), .A1 (n_0_0), .A2 (D[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n185), .A1 (n_0_0), .A2 (D[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n273), .A1 (n_0_0), .A2 (D[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n249), .A1 (n_0_0), .A2 (D[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n237), .A1 (n_0_0), .A2 (D[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n231), .A1 (n_0_0), .A2 (D[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n275), .A1 (n_0_0), .A2 (D[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n277), .A1 (n_0_0), .A2 (D[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n270), .A1 (n_0_0), .A2 (D[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n243), .A1 (n_0_0), .A2 (D[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n261), .A1 (n_0_0), .A2 (D[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n255), .A1 (n_0_0), .A2 (D[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n149), .A1 (n_0_0), .A2 (D[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n113), .A1 (n_0_0), .A2 (D[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n143), .A1 (n_0_0), .A2 (D[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n107), .A1 (n_0_0), .A2 (D[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n101), .A1 (n_0_0), .A2 (D[0]));
INV_X2 i_0_1 (.ZN (n_0_0), .A (rst));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (rst));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (CTS_n_tid1_2), .D (n_2));
DFF_X1 \Q_reg[1]  (.Q (Q[1]), .CK (CTS_n_tid1_2), .D (n_3));
DFF_X1 \Q_reg[2]  (.Q (Q[2]), .CK (CTS_n_tid1_2), .D (n_4));
DFF_X1 \Q_reg[3]  (.Q (Q[3]), .CK (CTS_n_tid1_2), .D (n_5));
DFF_X1 \Q_reg[4]  (.Q (Q[4]), .CK (CTS_n_tid1_2), .D (n_6));
DFF_X1 \Q_reg[5]  (.Q (Q[5]), .CK (CTS_n_tid1_2), .D (n_7));
DFF_X1 \Q_reg[6]  (.Q (Q[6]), .CK (CTS_n_tid1_2), .D (n_8));
DFF_X1 \Q_reg[7]  (.Q (Q[7]), .CK (CTS_n_tid1_2), .D (n_9));
DFF_X1 \Q_reg[8]  (.Q (Q[8]), .CK (CTS_n_tid1_2), .D (n_10));
DFF_X1 \Q_reg[9]  (.Q (Q[9]), .CK (CTS_n_tid1_2), .D (n_11));
DFF_X1 \Q_reg[10]  (.Q (Q[10]), .CK (CTS_n_tid1_2), .D (n_12));
DFF_X1 \Q_reg[11]  (.Q (Q[11]), .CK (CTS_n_tid1_2), .D (n_13));
DFF_X1 \Q_reg[12]  (.Q (Q[12]), .CK (CTS_n_tid1_2), .D (n_14));
DFF_X1 \Q_reg[13]  (.Q (Q[13]), .CK (CTS_n_tid1_2), .D (n_15));
DFF_X1 \Q_reg[14]  (.Q (Q[14]), .CK (CTS_n_tid1_2), .D (n_16));
DFF_X1 \Q_reg[15]  (.Q (Q[15]), .CK (CTS_n_tid1_2), .D (n_17));
DFF_X1 \Q_reg[16]  (.Q (Q[16]), .CK (CTS_n_tid1_2), .D (n_18));
DFF_X1 \Q_reg[17]  (.Q (Q[17]), .CK (CTS_n_tid1_2), .D (n_19));
DFF_X1 \Q_reg[18]  (.Q (Q[18]), .CK (CTS_n_tid1_2), .D (n_20));
DFF_X1 \Q_reg[19]  (.Q (Q[19]), .CK (CTS_n_tid1_2), .D (n_21));
DFF_X1 \Q_reg[20]  (.Q (Q[20]), .CK (CTS_n_tid1_2), .D (n_22));
DFF_X1 \Q_reg[21]  (.Q (Q[21]), .CK (CTS_n_tid1_2), .D (n_23));
DFF_X1 \Q_reg[22]  (.Q (Q[22]), .CK (CTS_n_tid1_2), .D (n_24));
DFF_X1 \Q_reg[23]  (.Q (Q[23]), .CK (CTS_n_tid1_2), .D (n_25));
DFF_X1 \Q_reg[24]  (.Q (Q[24]), .CK (CTS_n_tid1_2), .D (n_26));
DFF_X1 \Q_reg[25]  (.Q (Q[25]), .CK (CTS_n_tid1_2), .D (n_27));
DFF_X1 \Q_reg[26]  (.Q (Q[26]), .CK (CTS_n_tid1_2), .D (n_28));
DFF_X1 \Q_reg[27]  (.Q (Q[27]), .CK (CTS_n_tid1_2), .D (n_29));
DFF_X1 \Q_reg[28]  (.Q (Q[28]), .CK (CTS_n_tid1_2), .D (n_30));
DFF_X1 \Q_reg[29]  (.Q (Q[29]), .CK (CTS_n_tid1_2), .D (n_31));
DFF_X1 \Q_reg[30]  (.Q (Q[30]), .CK (CTS_n_tid1_2), .D (n_32));
DFF_X1 \Q_reg[31]  (.Q (Q[31]), .CK (CTS_n_tid1_2), .D (n_33));
CLKGATETST_X8 clk_gate_Q_reg (.GCK (CTS_n_tid1_3), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
CLKBUF_X3 CTS_L4_c_tid1_3 (.Z (CTS_n_tid1_2), .A (CTS_n_tid1_3));
CLKBUF_X1 CLOCK_slh__c42 (.Z (CLOCK_slh__n102), .A (CLOCK_slh__n101));
CLKBUF_X1 CLOCK_slh__c43 (.Z (CLOCK_slh__n103), .A (CLOCK_slh__n102));
CLKBUF_X1 CLOCK_slh__c44 (.Z (n_2), .A (CLOCK_slh__n103));
CLKBUF_X1 CLOCK_slh__c48 (.Z (CLOCK_slh__n108), .A (CLOCK_slh__n107));
CLKBUF_X1 CLOCK_slh__c49 (.Z (CLOCK_slh__n109), .A (CLOCK_slh__n108));
CLKBUF_X1 CLOCK_slh__c50 (.Z (n_3), .A (CLOCK_slh__n109));
CLKBUF_X1 CLOCK_slh__c54 (.Z (CLOCK_slh__n114), .A (CLOCK_slh__n113));
CLKBUF_X1 CLOCK_slh__c55 (.Z (CLOCK_slh__n115), .A (CLOCK_slh__n114));
CLKBUF_X1 CLOCK_slh__c56 (.Z (n_5), .A (CLOCK_slh__n115));
CLKBUF_X1 CLOCK_slh__c60 (.Z (CLOCK_slh__n120), .A (CLOCK_slh__n119));
CLKBUF_X1 CLOCK_slh__c61 (.Z (CLOCK_slh__n121), .A (CLOCK_slh__n120));
CLKBUF_X1 CLOCK_slh__c62 (.Z (n_26), .A (CLOCK_slh__n121));
CLKBUF_X1 CLOCK_slh__c66 (.Z (CLOCK_slh__n126), .A (CLOCK_slh__n125));
CLKBUF_X1 CLOCK_slh__c67 (.Z (CLOCK_slh__n127), .A (CLOCK_slh__n126));
CLKBUF_X1 CLOCK_slh__c68 (.Z (n_33), .A (CLOCK_slh__n127));
CLKBUF_X1 CLOCK_slh__c72 (.Z (CLOCK_slh__n132), .A (CLOCK_slh__n131));
CLKBUF_X1 CLOCK_slh__c73 (.Z (CLOCK_slh__n133), .A (CLOCK_slh__n132));
CLKBUF_X1 CLOCK_slh__c74 (.Z (n_27), .A (CLOCK_slh__n133));
CLKBUF_X1 CLOCK_slh__c78 (.Z (CLOCK_slh__n138), .A (CLOCK_slh__n137));
CLKBUF_X1 CLOCK_slh__c79 (.Z (CLOCK_slh__n139), .A (CLOCK_slh__n138));
CLKBUF_X1 CLOCK_slh__c80 (.Z (n_25), .A (CLOCK_slh__n139));
CLKBUF_X1 CLOCK_slh__c84 (.Z (CLOCK_slh__n144), .A (CLOCK_slh__n143));
CLKBUF_X1 CLOCK_slh__c85 (.Z (CLOCK_slh__n145), .A (CLOCK_slh__n144));
CLKBUF_X1 CLOCK_slh__c86 (.Z (n_4), .A (CLOCK_slh__n145));
CLKBUF_X1 CLOCK_slh__c90 (.Z (CLOCK_slh__n150), .A (CLOCK_slh__n149));
CLKBUF_X1 CLOCK_slh__c91 (.Z (CLOCK_slh__n151), .A (CLOCK_slh__n150));
CLKBUF_X1 CLOCK_slh__c92 (.Z (n_6), .A (CLOCK_slh__n151));
CLKBUF_X1 CLOCK_slh__c96 (.Z (CLOCK_slh__n156), .A (CLOCK_slh__n155));
CLKBUF_X1 CLOCK_slh__c97 (.Z (CLOCK_slh__n157), .A (CLOCK_slh__n156));
CLKBUF_X1 CLOCK_slh__c98 (.Z (n_31), .A (CLOCK_slh__n157));
CLKBUF_X1 CLOCK_slh__c102 (.Z (CLOCK_slh__n162), .A (CLOCK_slh__n161));
CLKBUF_X1 CLOCK_slh__c103 (.Z (CLOCK_slh__n163), .A (CLOCK_slh__n162));
CLKBUF_X1 CLOCK_slh__c104 (.Z (n_32), .A (CLOCK_slh__n163));
CLKBUF_X1 CLOCK_slh__c108 (.Z (CLOCK_slh__n168), .A (CLOCK_slh__n167));
CLKBUF_X1 CLOCK_slh__c109 (.Z (CLOCK_slh__n169), .A (CLOCK_slh__n168));
CLKBUF_X1 CLOCK_slh__c110 (.Z (n_30), .A (CLOCK_slh__n169));
CLKBUF_X1 CLOCK_slh__c114 (.Z (CLOCK_slh__n174), .A (CLOCK_slh__n173));
CLKBUF_X1 CLOCK_slh__c115 (.Z (CLOCK_slh__n175), .A (CLOCK_slh__n174));
CLKBUF_X1 CLOCK_slh__c116 (.Z (n_29), .A (CLOCK_slh__n175));
CLKBUF_X1 CLOCK_slh__c120 (.Z (CLOCK_slh__n180), .A (CLOCK_slh__n179));
CLKBUF_X1 CLOCK_slh__c121 (.Z (CLOCK_slh__n181), .A (CLOCK_slh__n180));
CLKBUF_X1 CLOCK_slh__c122 (.Z (n_24), .A (CLOCK_slh__n181));
CLKBUF_X1 CLOCK_slh__c126 (.Z (CLOCK_slh__n186), .A (CLOCK_slh__n185));
CLKBUF_X1 CLOCK_slh__c127 (.Z (CLOCK_slh__n187), .A (CLOCK_slh__n186));
CLKBUF_X1 CLOCK_slh__c128 (.Z (n_17), .A (CLOCK_slh__n187));
CLKBUF_X1 CLOCK_slh__c132 (.Z (CLOCK_slh__n192), .A (CLOCK_slh__n191));
CLKBUF_X1 CLOCK_slh__c133 (.Z (CLOCK_slh__n193), .A (CLOCK_slh__n192));
CLKBUF_X1 CLOCK_slh__c134 (.Z (n_21), .A (CLOCK_slh__n193));
CLKBUF_X1 CLOCK_slh__c138 (.Z (CLOCK_slh__n198), .A (CLOCK_slh__n197));
CLKBUF_X1 CLOCK_slh__c139 (.Z (CLOCK_slh__n199), .A (CLOCK_slh__n198));
CLKBUF_X1 CLOCK_slh__c140 (.Z (n_23), .A (CLOCK_slh__n199));
CLKBUF_X1 CLOCK_slh__c144 (.Z (CLOCK_slh__n203), .A (D[19]));
CLKBUF_X1 CLOCK_slh__c146 (.Z (CLOCK_slh__n205), .A (D[21]));
CLKBUF_X1 CLOCK_slh__c148 (.Z (CLOCK_slh__n208), .A (CLOCK_slh__n207));
CLKBUF_X1 CLOCK_slh__c149 (.Z (CLOCK_slh__n209), .A (CLOCK_slh__n208));
CLKBUF_X1 CLOCK_slh__c150 (.Z (n_22), .A (CLOCK_slh__n209));
CLKBUF_X1 CLOCK_slh__c154 (.Z (CLOCK_slh__n214), .A (CLOCK_slh__n213));
CLKBUF_X1 CLOCK_slh__c155 (.Z (CLOCK_slh__n215), .A (CLOCK_slh__n214));
CLKBUF_X1 CLOCK_slh__c156 (.Z (n_20), .A (CLOCK_slh__n215));
CLKBUF_X1 CLOCK_slh__c160 (.Z (CLOCK_slh__n220), .A (CLOCK_slh__n219));
CLKBUF_X1 CLOCK_slh__c161 (.Z (CLOCK_slh__n221), .A (CLOCK_slh__n220));
CLKBUF_X1 CLOCK_slh__c162 (.Z (n_18), .A (CLOCK_slh__n221));
CLKBUF_X1 CLOCK_slh__c166 (.Z (CLOCK_slh__n226), .A (CLOCK_slh__n225));
CLKBUF_X1 CLOCK_slh__c167 (.Z (CLOCK_slh__n227), .A (CLOCK_slh__n226));
CLKBUF_X1 CLOCK_slh__c168 (.Z (n_19), .A (CLOCK_slh__n227));
CLKBUF_X1 CLOCK_slh__c172 (.Z (CLOCK_slh__n232), .A (CLOCK_slh__n231));
CLKBUF_X1 CLOCK_slh__c173 (.Z (CLOCK_slh__n233), .A (CLOCK_slh__n232));
CLKBUF_X1 CLOCK_slh__c174 (.Z (n_13), .A (CLOCK_slh__n233));
CLKBUF_X1 CLOCK_slh__c178 (.Z (CLOCK_slh__n238), .A (CLOCK_slh__n237));
CLKBUF_X1 CLOCK_slh__c179 (.Z (CLOCK_slh__n239), .A (CLOCK_slh__n238));
CLKBUF_X1 CLOCK_slh__c180 (.Z (n_14), .A (CLOCK_slh__n239));
CLKBUF_X1 CLOCK_slh__c184 (.Z (CLOCK_slh__n244), .A (CLOCK_slh__n243));
CLKBUF_X1 CLOCK_slh__c185 (.Z (CLOCK_slh__n245), .A (CLOCK_slh__n244));
CLKBUF_X1 CLOCK_slh__c186 (.Z (n_9), .A (CLOCK_slh__n245));
CLKBUF_X1 CLOCK_slh__c190 (.Z (CLOCK_slh__n250), .A (CLOCK_slh__n249));
CLKBUF_X1 CLOCK_slh__c191 (.Z (CLOCK_slh__n251), .A (CLOCK_slh__n250));
CLKBUF_X1 CLOCK_slh__c192 (.Z (n_15), .A (CLOCK_slh__n251));
CLKBUF_X1 CLOCK_slh__c196 (.Z (CLOCK_slh__n256), .A (CLOCK_slh__n255));
CLKBUF_X1 CLOCK_slh__c197 (.Z (CLOCK_slh__n257), .A (CLOCK_slh__n256));
CLKBUF_X1 CLOCK_slh__c198 (.Z (n_7), .A (CLOCK_slh__n257));
CLKBUF_X1 CLOCK_slh__c202 (.Z (CLOCK_slh__n262), .A (CLOCK_slh__n261));
CLKBUF_X1 CLOCK_slh__c203 (.Z (CLOCK_slh__n263), .A (CLOCK_slh__n262));
CLKBUF_X1 CLOCK_slh__c204 (.Z (n_8), .A (CLOCK_slh__n263));
CLKBUF_X1 CLOCK_slh__c208 (.Z (CLOCK_slh__n268), .A (CLOCK_slh__n267));
CLKBUF_X1 CLOCK_slh__c209 (.Z (CLOCK_slh__n269), .A (CLOCK_slh__n268));
CLKBUF_X1 CLOCK_slh__c210 (.Z (n_28), .A (CLOCK_slh__n269));
CLKBUF_X1 CLOCK_slh__c211 (.Z (CLOCK_slh__n271), .A (CLOCK_slh__n270));
CLKBUF_X1 CLOCK_slh__c212 (.Z (CLOCK_slh__n272), .A (CLOCK_slh__n271));
CLKBUF_X1 CLOCK_slh__c213 (.Z (n_10), .A (CLOCK_slh__n272));
CLKBUF_X1 CLOCK_slh__c214 (.Z (CLOCK_slh__n274), .A (CLOCK_slh__n273));
CLKBUF_X1 CLOCK_slh__c215 (.Z (n_16), .A (CLOCK_slh__n274));
CLKBUF_X1 CLOCK_slh__c216 (.Z (CLOCK_slh__n276), .A (CLOCK_slh__n275));
CLKBUF_X1 CLOCK_slh__c217 (.Z (n_12), .A (CLOCK_slh__n276));
CLKBUF_X1 CLOCK_slh__c218 (.Z (CLOCK_slh__n278), .A (CLOCK_slh__n277));
CLKBUF_X1 CLOCK_slh__c219 (.Z (n_11), .A (CLOCK_slh__n278));

endmodule //buffer

module buffer__0_68 (clk_CTS_0_PP_0, clk, rst, en, D, Q);

output [31:0] Q;
input [31:0] D;
input clk;
input en;
input rst;
input clk_CTS_0_PP_0;
wire n_0_0;
wire n_1;
wire CTS_n_tid0_2;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid0_3;
wire CLOCK_slh__n377;
wire CLOCK_slh__n382;
wire CLOCK_slh__n383;
wire CLOCK_slh__n376;
wire CLOCK_slh__n378;
wire CLOCK_slh__n384;
wire CLOCK_slh__n388;
wire CLOCK_slh__n389;
wire CLOCK_slh__n390;
wire CLOCK_slh__n394;
wire CLOCK_slh__n395;
wire CLOCK_slh__n396;
wire CLOCK_slh__n400;
wire CLOCK_slh__n401;
wire CLOCK_slh__n402;
wire CLOCK_slh__n406;
wire CLOCK_slh__n407;
wire CLOCK_slh__n408;
wire CLOCK_slh__n412;
wire CLOCK_slh__n413;
wire CLOCK_slh__n414;
wire CLOCK_slh__n418;
wire CLOCK_slh__n420;
wire CLOCK_slh__n422;
wire CLOCK_slh__n424;
wire CLOCK_slh__n425;
wire CLOCK_slh__n426;
wire CLOCK_slh__n430;
wire CLOCK_slh__n431;
wire CLOCK_slh__n432;
wire CLOCK_slh__n436;
wire CLOCK_slh__n437;
wire CLOCK_slh__n438;
wire CLOCK_slh__n442;
wire CLOCK_slh__n443;
wire CLOCK_slh__n444;
wire CLOCK_slh__n448;
wire CLOCK_slh__n449;
wire CLOCK_slh__n450;
wire CLOCK_slh__n454;
wire CLOCK_slh__n455;
wire CLOCK_slh__n456;
wire CLOCK_slh__n460;
wire CLOCK_slh__n461;
wire CLOCK_slh__n462;
wire CLOCK_slh__n466;
wire CLOCK_slh__n467;
wire CLOCK_slh__n468;
wire CLOCK_slh__n472;
wire CLOCK_slh__n473;
wire CLOCK_slh__n474;
wire CLOCK_slh__n478;
wire CLOCK_slh__n480;
wire CLOCK_slh__n481;
wire CLOCK_slh__n482;
wire CLOCK_slh__n486;
wire CLOCK_slh__n487;
wire CLOCK_slh__n488;
wire CLOCK_slh__n492;
wire CLOCK_slh__n494;
wire CLOCK_slh__n495;
wire CLOCK_slh__n496;
wire CLOCK_slh__n500;
wire CLOCK_slh__n501;
wire CLOCK_slh__n502;
wire CLOCK_slh__n506;
wire CLOCK_slh__n507;
wire CLOCK_slh__n508;
wire CLOCK_slh__n512;
wire CLOCK_slh__n513;
wire CLOCK_slh__n514;
wire CLOCK_slh__n518;
wire CLOCK_slh__n519;
wire CLOCK_slh__n520;
wire CLOCK_slh__n524;
wire CLOCK_slh__n525;
wire CLOCK_slh__n526;
wire CLOCK_slh__n530;
wire CLOCK_slh__n531;
wire CLOCK_slh__n532;
wire CLOCK_slh__n533;
wire CLOCK_slh__n534;
wire CLOCK_slh__n535;
wire CLOCK_slh__n536;
wire CLOCK_slh__n537;
wire CLOCK_slh__n538;
wire CLOCK_slh__n539;
wire CLOCK_slh__n540;
wire CLOCK_slh__n541;
wire CLOCK_slh__n542;
wire CLOCK_slh__n543;
wire CLOCK_slh__n544;
wire CLOCK_slh__n545;
wire CLOCK_slh__n546;
wire CLOCK_slh__n547;
wire CLOCK_slh__n548;
wire CLOCK_slh__n549;
wire CLOCK_slh__n550;
wire CLOCK_slh__n551;
wire CLOCK_slh__n552;
wire CLOCK_slh__n553;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n412), .A1 (n_0_0), .A2 (CLOCK_slh__n422));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n406), .A1 (n_0_0), .A2 (CLOCK_slh__n418));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n480), .A1 (n_0_0), .A2 (CLOCK_slh__n492));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n400), .A1 (n_0_0), .A2 (CLOCK_slh__n420));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n494), .A1 (n_0_0), .A2 (D[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n436), .A1 (n_0_0), .A2 (CLOCK_slh__n478));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n536), .A1 (n_0_0), .A2 (D[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n530), .A1 (n_0_0), .A2 (D[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n533), .A1 (n_0_0), .A2 (D[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n548), .A1 (n_0_0), .A2 (D[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n472), .A1 (n_0_0), .A2 (D[21]));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n545), .A1 (n_0_0), .A2 (D[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n448), .A1 (n_0_0), .A2 (D[19]));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n466), .A1 (n_0_0), .A2 (D[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n460), .A1 (n_0_0), .A2 (D[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n454), .A1 (n_0_0), .A2 (D[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n486), .A1 (n_0_0), .A2 (D[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n442), .A1 (n_0_0), .A2 (D[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n524), .A1 (n_0_0), .A2 (D[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n542), .A1 (n_0_0), .A2 (D[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n518), .A1 (n_0_0), .A2 (D[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n500), .A1 (n_0_0), .A2 (D[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n506), .A1 (n_0_0), .A2 (D[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n551), .A1 (n_0_0), .A2 (D[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n424), .A1 (n_0_0), .A2 (D[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n382), .A1 (n_0_0), .A2 (D[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n430), .A1 (n_0_0), .A2 (D[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n394), .A1 (n_0_0), .A2 (D[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n376), .A1 (n_0_0), .A2 (D[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n388), .A1 (n_0_0), .A2 (D[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n512), .A1 (n_0_0), .A2 (D[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n539), .A1 (n_0_0), .A2 (D[0]));
INV_X2 i_0_1 (.ZN (n_0_0), .A (rst));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (rst));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (CTS_n_tid0_2), .D (n_2));
DFF_X1 \Q_reg[1]  (.Q (Q[1]), .CK (CTS_n_tid0_2), .D (n_3));
DFF_X1 \Q_reg[2]  (.Q (Q[2]), .CK (CTS_n_tid0_2), .D (n_4));
DFF_X1 \Q_reg[3]  (.Q (Q[3]), .CK (CTS_n_tid0_2), .D (n_5));
DFF_X1 \Q_reg[4]  (.Q (Q[4]), .CK (CTS_n_tid0_2), .D (n_6));
DFF_X1 \Q_reg[5]  (.Q (Q[5]), .CK (CTS_n_tid0_2), .D (n_7));
DFF_X1 \Q_reg[6]  (.Q (Q[6]), .CK (CTS_n_tid0_2), .D (n_8));
DFF_X1 \Q_reg[7]  (.Q (Q[7]), .CK (CTS_n_tid0_2), .D (n_9));
DFF_X1 \Q_reg[8]  (.Q (Q[8]), .CK (CTS_n_tid0_2), .D (n_10));
DFF_X1 \Q_reg[9]  (.Q (Q[9]), .CK (CTS_n_tid0_2), .D (n_11));
DFF_X1 \Q_reg[10]  (.Q (Q[10]), .CK (CTS_n_tid0_2), .D (n_12));
DFF_X1 \Q_reg[11]  (.Q (Q[11]), .CK (CTS_n_tid0_2), .D (n_13));
DFF_X1 \Q_reg[12]  (.Q (Q[12]), .CK (CTS_n_tid0_2), .D (n_14));
DFF_X1 \Q_reg[13]  (.Q (Q[13]), .CK (CTS_n_tid0_2), .D (n_15));
DFF_X1 \Q_reg[14]  (.Q (Q[14]), .CK (CTS_n_tid0_2), .D (n_16));
DFF_X1 \Q_reg[15]  (.Q (Q[15]), .CK (CTS_n_tid0_2), .D (n_17));
DFF_X1 \Q_reg[16]  (.Q (Q[16]), .CK (CTS_n_tid0_2), .D (n_18));
DFF_X1 \Q_reg[17]  (.Q (Q[17]), .CK (CTS_n_tid0_2), .D (n_19));
DFF_X1 \Q_reg[18]  (.Q (Q[18]), .CK (CTS_n_tid0_2), .D (n_20));
DFF_X1 \Q_reg[19]  (.Q (Q[19]), .CK (CTS_n_tid0_2), .D (n_21));
DFF_X1 \Q_reg[20]  (.Q (Q[20]), .CK (CTS_n_tid0_2), .D (n_22));
DFF_X1 \Q_reg[21]  (.Q (Q[21]), .CK (CTS_n_tid0_2), .D (n_23));
DFF_X1 \Q_reg[22]  (.Q (Q[22]), .CK (CTS_n_tid0_2), .D (n_24));
DFF_X1 \Q_reg[23]  (.Q (Q[23]), .CK (CTS_n_tid0_2), .D (n_25));
DFF_X1 \Q_reg[24]  (.Q (Q[24]), .CK (CTS_n_tid0_2), .D (n_26));
DFF_X1 \Q_reg[25]  (.Q (Q[25]), .CK (CTS_n_tid0_2), .D (n_27));
DFF_X1 \Q_reg[26]  (.Q (Q[26]), .CK (CTS_n_tid0_2), .D (n_28));
DFF_X1 \Q_reg[27]  (.Q (Q[27]), .CK (CTS_n_tid0_2), .D (n_29));
DFF_X1 \Q_reg[28]  (.Q (Q[28]), .CK (CTS_n_tid0_2), .D (n_30));
DFF_X1 \Q_reg[29]  (.Q (Q[29]), .CK (CTS_n_tid0_2), .D (n_31));
DFF_X1 \Q_reg[30]  (.Q (Q[30]), .CK (CTS_n_tid0_2), .D (n_32));
DFF_X1 \Q_reg[31]  (.Q (Q[31]), .CK (CTS_n_tid0_2), .D (n_33));
CLKGATETST_X8 clk_gate_Q_reg (.GCK (CTS_n_tid0_3), .CK (clk_CTS_0_PP_0), .E (n_1), .SE (1'b0 ));
CLKBUF_X3 CTS_L4_c_tid0_3 (.Z (CTS_n_tid0_2), .A (CTS_n_tid0_3));
CLKBUF_X1 CLOCK_slh__c326 (.Z (CLOCK_slh__n378), .A (CLOCK_slh__n377));
CLKBUF_X1 CLOCK_slh__c325 (.Z (CLOCK_slh__n377), .A (CLOCK_slh__n376));
CLKBUF_X1 CLOCK_slh__c327 (.Z (n_5), .A (CLOCK_slh__n378));
CLKBUF_X1 CLOCK_slh__c331 (.Z (CLOCK_slh__n383), .A (CLOCK_slh__n382));
CLKBUF_X1 CLOCK_slh__c332 (.Z (CLOCK_slh__n384), .A (CLOCK_slh__n383));
CLKBUF_X1 CLOCK_slh__c333 (.Z (n_8), .A (CLOCK_slh__n384));
CLKBUF_X1 CLOCK_slh__c337 (.Z (CLOCK_slh__n389), .A (CLOCK_slh__n388));
CLKBUF_X1 CLOCK_slh__c338 (.Z (CLOCK_slh__n390), .A (CLOCK_slh__n389));
CLKBUF_X1 CLOCK_slh__c339 (.Z (n_4), .A (CLOCK_slh__n390));
CLKBUF_X1 CLOCK_slh__c343 (.Z (CLOCK_slh__n395), .A (CLOCK_slh__n394));
CLKBUF_X1 CLOCK_slh__c344 (.Z (CLOCK_slh__n396), .A (CLOCK_slh__n395));
CLKBUF_X1 CLOCK_slh__c345 (.Z (n_6), .A (CLOCK_slh__n396));
CLKBUF_X1 CLOCK_slh__c349 (.Z (CLOCK_slh__n401), .A (CLOCK_slh__n400));
CLKBUF_X1 CLOCK_slh__c350 (.Z (CLOCK_slh__n402), .A (CLOCK_slh__n401));
CLKBUF_X1 CLOCK_slh__c351 (.Z (n_30), .A (CLOCK_slh__n402));
CLKBUF_X1 CLOCK_slh__c355 (.Z (CLOCK_slh__n407), .A (CLOCK_slh__n406));
CLKBUF_X1 CLOCK_slh__c356 (.Z (CLOCK_slh__n408), .A (CLOCK_slh__n407));
CLKBUF_X1 CLOCK_slh__c357 (.Z (n_32), .A (CLOCK_slh__n408));
CLKBUF_X1 CLOCK_slh__c361 (.Z (CLOCK_slh__n413), .A (CLOCK_slh__n412));
CLKBUF_X1 CLOCK_slh__c362 (.Z (CLOCK_slh__n414), .A (CLOCK_slh__n413));
CLKBUF_X1 CLOCK_slh__c363 (.Z (n_33), .A (CLOCK_slh__n414));
CLKBUF_X1 CLOCK_slh__c367 (.Z (CLOCK_slh__n418), .A (D[30]));
CLKBUF_X1 CLOCK_slh__c369 (.Z (CLOCK_slh__n420), .A (D[28]));
CLKBUF_X1 CLOCK_slh__c371 (.Z (CLOCK_slh__n422), .A (D[31]));
CLKBUF_X1 CLOCK_slh__c373 (.Z (CLOCK_slh__n425), .A (CLOCK_slh__n424));
CLKBUF_X1 CLOCK_slh__c374 (.Z (CLOCK_slh__n426), .A (CLOCK_slh__n425));
CLKBUF_X1 CLOCK_slh__c375 (.Z (n_9), .A (CLOCK_slh__n426));
CLKBUF_X1 CLOCK_slh__c379 (.Z (CLOCK_slh__n431), .A (CLOCK_slh__n430));
CLKBUF_X1 CLOCK_slh__c380 (.Z (CLOCK_slh__n432), .A (CLOCK_slh__n431));
CLKBUF_X1 CLOCK_slh__c381 (.Z (n_7), .A (CLOCK_slh__n432));
CLKBUF_X1 CLOCK_slh__c385 (.Z (CLOCK_slh__n437), .A (CLOCK_slh__n436));
CLKBUF_X1 CLOCK_slh__c386 (.Z (CLOCK_slh__n438), .A (CLOCK_slh__n437));
CLKBUF_X1 CLOCK_slh__c387 (.Z (n_28), .A (CLOCK_slh__n438));
CLKBUF_X1 CLOCK_slh__c391 (.Z (CLOCK_slh__n443), .A (CLOCK_slh__n442));
CLKBUF_X1 CLOCK_slh__c392 (.Z (CLOCK_slh__n444), .A (CLOCK_slh__n443));
CLKBUF_X1 CLOCK_slh__c393 (.Z (n_16), .A (CLOCK_slh__n444));
CLKBUF_X1 CLOCK_slh__c397 (.Z (CLOCK_slh__n449), .A (CLOCK_slh__n448));
CLKBUF_X1 CLOCK_slh__c398 (.Z (CLOCK_slh__n450), .A (CLOCK_slh__n449));
CLKBUF_X1 CLOCK_slh__c399 (.Z (n_21), .A (CLOCK_slh__n450));
CLKBUF_X1 CLOCK_slh__c403 (.Z (CLOCK_slh__n455), .A (CLOCK_slh__n454));
CLKBUF_X1 CLOCK_slh__c404 (.Z (CLOCK_slh__n456), .A (CLOCK_slh__n455));
CLKBUF_X1 CLOCK_slh__c405 (.Z (n_18), .A (CLOCK_slh__n456));
CLKBUF_X1 CLOCK_slh__c409 (.Z (CLOCK_slh__n461), .A (CLOCK_slh__n460));
CLKBUF_X1 CLOCK_slh__c410 (.Z (CLOCK_slh__n462), .A (CLOCK_slh__n461));
CLKBUF_X1 CLOCK_slh__c411 (.Z (n_19), .A (CLOCK_slh__n462));
CLKBUF_X1 CLOCK_slh__c415 (.Z (CLOCK_slh__n467), .A (CLOCK_slh__n466));
CLKBUF_X1 CLOCK_slh__c416 (.Z (CLOCK_slh__n468), .A (CLOCK_slh__n467));
CLKBUF_X1 CLOCK_slh__c417 (.Z (n_20), .A (CLOCK_slh__n468));
CLKBUF_X1 CLOCK_slh__c421 (.Z (CLOCK_slh__n473), .A (CLOCK_slh__n472));
CLKBUF_X1 CLOCK_slh__c422 (.Z (CLOCK_slh__n474), .A (CLOCK_slh__n473));
CLKBUF_X1 CLOCK_slh__c423 (.Z (n_23), .A (CLOCK_slh__n474));
CLKBUF_X1 CLOCK_slh__c427 (.Z (CLOCK_slh__n478), .A (D[26]));
CLKBUF_X1 CLOCK_slh__c429 (.Z (CLOCK_slh__n481), .A (CLOCK_slh__n480));
CLKBUF_X1 CLOCK_slh__c430 (.Z (CLOCK_slh__n482), .A (CLOCK_slh__n481));
CLKBUF_X1 CLOCK_slh__c431 (.Z (n_31), .A (CLOCK_slh__n482));
CLKBUF_X1 CLOCK_slh__c435 (.Z (CLOCK_slh__n487), .A (CLOCK_slh__n486));
CLKBUF_X1 CLOCK_slh__c436 (.Z (CLOCK_slh__n488), .A (CLOCK_slh__n487));
CLKBUF_X1 CLOCK_slh__c437 (.Z (n_17), .A (CLOCK_slh__n488));
CLKBUF_X1 CLOCK_slh__c441 (.Z (CLOCK_slh__n492), .A (D[29]));
CLKBUF_X1 CLOCK_slh__c443 (.Z (CLOCK_slh__n495), .A (CLOCK_slh__n494));
CLKBUF_X1 CLOCK_slh__c444 (.Z (CLOCK_slh__n496), .A (CLOCK_slh__n495));
CLKBUF_X1 CLOCK_slh__c445 (.Z (n_29), .A (CLOCK_slh__n496));
CLKBUF_X1 CLOCK_slh__c449 (.Z (CLOCK_slh__n501), .A (CLOCK_slh__n500));
CLKBUF_X1 CLOCK_slh__c450 (.Z (CLOCK_slh__n502), .A (CLOCK_slh__n501));
CLKBUF_X1 CLOCK_slh__c451 (.Z (n_12), .A (CLOCK_slh__n502));
CLKBUF_X1 CLOCK_slh__c455 (.Z (CLOCK_slh__n507), .A (CLOCK_slh__n506));
CLKBUF_X1 CLOCK_slh__c456 (.Z (CLOCK_slh__n508), .A (CLOCK_slh__n507));
CLKBUF_X1 CLOCK_slh__c457 (.Z (n_11), .A (CLOCK_slh__n508));
CLKBUF_X1 CLOCK_slh__c461 (.Z (CLOCK_slh__n513), .A (CLOCK_slh__n512));
CLKBUF_X1 CLOCK_slh__c462 (.Z (CLOCK_slh__n514), .A (CLOCK_slh__n513));
CLKBUF_X1 CLOCK_slh__c463 (.Z (n_3), .A (CLOCK_slh__n514));
CLKBUF_X1 CLOCK_slh__c467 (.Z (CLOCK_slh__n519), .A (CLOCK_slh__n518));
CLKBUF_X1 CLOCK_slh__c468 (.Z (CLOCK_slh__n520), .A (CLOCK_slh__n519));
CLKBUF_X1 CLOCK_slh__c469 (.Z (n_13), .A (CLOCK_slh__n520));
CLKBUF_X1 CLOCK_slh__c473 (.Z (CLOCK_slh__n525), .A (CLOCK_slh__n524));
CLKBUF_X1 CLOCK_slh__c474 (.Z (CLOCK_slh__n526), .A (CLOCK_slh__n525));
CLKBUF_X1 CLOCK_slh__c475 (.Z (n_15), .A (CLOCK_slh__n526));
CLKBUF_X1 CLOCK_slh__c479 (.Z (CLOCK_slh__n531), .A (CLOCK_slh__n530));
CLKBUF_X1 CLOCK_slh__c480 (.Z (CLOCK_slh__n532), .A (CLOCK_slh__n531));
CLKBUF_X1 CLOCK_slh__c481 (.Z (n_26), .A (CLOCK_slh__n532));
CLKBUF_X1 CLOCK_slh__c482 (.Z (CLOCK_slh__n534), .A (CLOCK_slh__n533));
CLKBUF_X1 CLOCK_slh__c483 (.Z (CLOCK_slh__n535), .A (CLOCK_slh__n534));
CLKBUF_X1 CLOCK_slh__c484 (.Z (n_25), .A (CLOCK_slh__n535));
CLKBUF_X1 CLOCK_slh__c485 (.Z (CLOCK_slh__n537), .A (CLOCK_slh__n536));
CLKBUF_X1 CLOCK_slh__c486 (.Z (CLOCK_slh__n538), .A (CLOCK_slh__n537));
CLKBUF_X1 CLOCK_slh__c487 (.Z (n_27), .A (CLOCK_slh__n538));
CLKBUF_X1 CLOCK_slh__c488 (.Z (CLOCK_slh__n540), .A (CLOCK_slh__n539));
CLKBUF_X1 CLOCK_slh__c489 (.Z (CLOCK_slh__n541), .A (CLOCK_slh__n540));
CLKBUF_X1 CLOCK_slh__c490 (.Z (n_2), .A (CLOCK_slh__n541));
CLKBUF_X1 CLOCK_slh__c491 (.Z (CLOCK_slh__n543), .A (CLOCK_slh__n542));
CLKBUF_X1 CLOCK_slh__c492 (.Z (CLOCK_slh__n544), .A (CLOCK_slh__n543));
CLKBUF_X1 CLOCK_slh__c493 (.Z (n_14), .A (CLOCK_slh__n544));
CLKBUF_X1 CLOCK_slh__c494 (.Z (CLOCK_slh__n546), .A (CLOCK_slh__n545));
CLKBUF_X1 CLOCK_slh__c495 (.Z (CLOCK_slh__n547), .A (CLOCK_slh__n546));
CLKBUF_X1 CLOCK_slh__c496 (.Z (n_22), .A (CLOCK_slh__n547));
CLKBUF_X1 CLOCK_slh__c497 (.Z (CLOCK_slh__n549), .A (CLOCK_slh__n548));
CLKBUF_X1 CLOCK_slh__c498 (.Z (CLOCK_slh__n550), .A (CLOCK_slh__n549));
CLKBUF_X1 CLOCK_slh__c499 (.Z (n_24), .A (CLOCK_slh__n550));
CLKBUF_X1 CLOCK_slh__c500 (.Z (CLOCK_slh__n552), .A (CLOCK_slh__n551));
CLKBUF_X1 CLOCK_slh__c501 (.Z (CLOCK_slh__n553), .A (CLOCK_slh__n552));
CLKBUF_X1 CLOCK_slh__c502 (.Z (n_10), .A (CLOCK_slh__n553));

endmodule //buffer__0_68

module simpleMultiplier (clk, rst, en, a, b, c);

output [63:0] c;
input [31:0] a;
input [31:0] b;
input clk;
input en;
input rst;
wire CTS_n_tid0_3;
wire CLOCK_slh_n232;
wire CLOCK_slh_n247;
wire CLOCK_slh_n262;
wire CLOCK_slh_n242;
wire CLOCK_slh_n257;
wire CLOCK_slh_n280;
wire CLOCK_slh_n237;
wire CLOCK_slh_n252;
wire CLOCK_slh_n197;
wire CLOCK_slh_n271;
wire CLOCK_slh_n210;
wire CLOCK_slh_n177;
wire CLOCK_slh_n192;
wire CLOCK_slh_n132;
wire CLOCK_slh_n162;
wire CLOCK_slh_n157;
wire CLOCK_slh_n172;
wire CLOCK_slh_n167;
wire CLOCK_slh_n142;
wire CLOCK_slh_n127;
wire CLOCK_slh_n137;
wire CLOCK_slh_n182;
wire CLOCK_slh_n227;
wire CLOCK_slh_n285;
wire CLOCK_slh_n295;
wire CLOCK_slh_n290;
wire CLOCK_slh_n187;
wire CLOCK_slh_n152;
wire CLOCK_slh_n122;
wire CLOCK_slh_n147;
wire CLOCK_slh_n112;
wire CLOCK_slh_n117;
wire \a_out[31] ;
wire \a_out[30] ;
wire \a_out[29] ;
wire \a_out[28] ;
wire \a_out[27] ;
wire \a_out[26] ;
wire \a_out[25] ;
wire \a_out[24] ;
wire \a_out[23] ;
wire \a_out[22] ;
wire \a_out[21] ;
wire \a_out[20] ;
wire \a_out[19] ;
wire \a_out[18] ;
wire \a_out[17] ;
wire \a_out[16] ;
wire \a_out[15] ;
wire \a_out[14] ;
wire \a_out[13] ;
wire \a_out[12] ;
wire \a_out[11] ;
wire \a_out[10] ;
wire \a_out[9] ;
wire \a_out[8] ;
wire \a_out[7] ;
wire \a_out[6] ;
wire \a_out[5] ;
wire \a_out[4] ;
wire \a_out[3] ;
wire \a_out[2] ;
wire \a_out[1] ;
wire \a_out[0] ;
wire \b_out[31] ;
wire \b_out[30] ;
wire \b_out[29] ;
wire \b_out[28] ;
wire \b_out[27] ;
wire \b_out[26] ;
wire \b_out[25] ;
wire \b_out[24] ;
wire \b_out[23] ;
wire \b_out[22] ;
wire \b_out[21] ;
wire \b_out[20] ;
wire \b_out[19] ;
wire \b_out[18] ;
wire \b_out[17] ;
wire \b_out[16] ;
wire \b_out[15] ;
wire \b_out[14] ;
wire \b_out[13] ;
wire \b_out[12] ;
wire \b_out[11] ;
wire \b_out[10] ;
wire \b_out[9] ;
wire \b_out[8] ;
wire \b_out[7] ;
wire \b_out[6] ;
wire \b_out[5] ;
wire \b_out[4] ;
wire \b_out[3] ;
wire \b_out[2] ;
wire \b_out[1] ;
wire \b_out[0] ;
wire \c_out[63] ;
wire \c_out[62] ;
wire \c_out[61] ;
wire \c_out[60] ;
wire \c_out[59] ;
wire \c_out[58] ;
wire \c_out[57] ;
wire \c_out[56] ;
wire \c_out[55] ;
wire \c_out[54] ;
wire \c_out[53] ;
wire \c_out[52] ;
wire \c_out[51] ;
wire \c_out[50] ;
wire \c_out[49] ;
wire \c_out[48] ;
wire \c_out[47] ;
wire \c_out[46] ;
wire \c_out[45] ;
wire \c_out[44] ;
wire \c_out[43] ;
wire \c_out[42] ;
wire \c_out[41] ;
wire \c_out[40] ;
wire \c_out[39] ;
wire \c_out[38] ;
wire \c_out[37] ;
wire \c_out[36] ;
wire \c_out[35] ;
wire \c_out[34] ;
wire \c_out[33] ;
wire \c_out[32] ;
wire \c_out[31] ;
wire \c_out[30] ;
wire \c_out[29] ;
wire \c_out[28] ;
wire \c_out[27] ;
wire \c_out[26] ;
wire \c_out[25] ;
wire \c_out[24] ;
wire \c_out[23] ;
wire \c_out[22] ;
wire \c_out[21] ;
wire \c_out[20] ;
wire \c_out[19] ;
wire \c_out[18] ;
wire \c_out[17] ;
wire \c_out[16] ;
wire \c_out[15] ;
wire \c_out[14] ;
wire \c_out[13] ;
wire \c_out[12] ;
wire \c_out[11] ;
wire \c_out[10] ;
wire \c_out[9] ;
wire \c_out[8] ;
wire \c_out[7] ;
wire \c_out[6] ;
wire \c_out[5] ;
wire \c_out[4] ;
wire \c_out[3] ;
wire \c_out[2] ;
wire \c_out[1] ;
wire \c_out[0] ;
wire CTS_n_tid0_24;


buffer__parameterized0 outReg (.Q ({c[63], c[62], c[61], c[60], c[59], c[58], c[57], 
    c[56], c[55], c[54], c[53], c[52], c[51], c[50], c[49], c[48], c[47], c[46], 
    c[45], c[44], c[43], c[42], c[41], c[40], c[39], c[38], c[37], c[36], c[35], 
    c[34], c[33], c[32], c[31], c[30], c[29], c[28], c[27], c[26], c[25], c[24], 
    c[23], c[22], c[21], c[20], c[19], c[18], c[17], c[16], c[15], c[14], c[13], 
    c[12], c[11], c[10], c[9], c[8], c[7], c[6], c[5], c[4], c[3], c[2], c[1], c[0]})
    , .D ({\c_out[63] , \c_out[62] , \c_out[61] , \c_out[60] , \c_out[59] , \c_out[58] , 
    \c_out[57] , \c_out[56] , \c_out[55] , \c_out[54] , \c_out[53] , \c_out[52] , 
    \c_out[51] , \c_out[50] , \c_out[49] , \c_out[48] , \c_out[47] , \c_out[46] , 
    \c_out[45] , \c_out[44] , \c_out[43] , \c_out[42] , \c_out[41] , \c_out[40] , 
    \c_out[39] , \c_out[38] , \c_out[37] , \c_out[36] , \c_out[35] , \c_out[34] , 
    \c_out[33] , \c_out[32] , \c_out[31] , \c_out[30] , \c_out[29] , \c_out[28] , 
    \c_out[27] , \c_out[26] , \c_out[25] , \c_out[24] , \c_out[23] , \c_out[22] , 
    \c_out[21] , \c_out[20] , \c_out[19] , \c_out[18] , \c_out[17] , \c_out[16] , 
    \c_out[15] , \c_out[14] , \c_out[13] , \c_out[12] , \c_out[11] , \c_out[10] , 
    \c_out[9] , \c_out[8] , \c_out[7] , \c_out[6] , \c_out[5] , \c_out[4] , \c_out[3] , 
    \c_out[2] , \c_out[1] , \c_out[0] }), .en (en), .rst (rst), .clk_CTS_0_PP_0 (CTS_n_tid0_24));
multOperator M64 (.c ({\c_out[63] , \c_out[62] , \c_out[61] , \c_out[60] , \c_out[59] , 
    \c_out[58] , \c_out[57] , \c_out[56] , \c_out[55] , \c_out[54] , \c_out[53] , 
    \c_out[52] , \c_out[51] , \c_out[50] , \c_out[49] , \c_out[48] , \c_out[47] , 
    \c_out[46] , \c_out[45] , \c_out[44] , \c_out[43] , \c_out[42] , \c_out[41] , 
    \c_out[40] , \c_out[39] , \c_out[38] , \c_out[37] , \c_out[36] , \c_out[35] , 
    \c_out[34] , \c_out[33] , \c_out[32] , \c_out[31] , \c_out[30] , \c_out[29] , 
    \c_out[28] , \c_out[27] , \c_out[26] , \c_out[25] , \c_out[24] , \c_out[23] , 
    \c_out[22] , \c_out[21] , \c_out[20] , \c_out[19] , \c_out[18] , \c_out[17] , 
    \c_out[16] , \c_out[15] , \c_out[14] , \c_out[13] , \c_out[12] , \c_out[11] , 
    \c_out[10] , \c_out[9] , \c_out[8] , \c_out[7] , \c_out[6] , \c_out[5] , \c_out[4] , 
    \c_out[3] , \c_out[2] , \c_out[1] , \c_out[0] }), .clk_CTS_0_PP_0 (CTS_n_tid0_3)
    , .clk_CTS_0_PP_9 (CTS_n_tid0_24), .a ({\a_out[31] , \a_out[30] , \a_out[29] , 
    \a_out[28] , \a_out[27] , \a_out[26] , \a_out[25] , \a_out[24] , \a_out[23] , 
    \a_out[22] , \a_out[21] , \a_out[20] , \a_out[19] , \a_out[18] , \a_out[17] , 
    \a_out[16] , \a_out[15] , \a_out[14] , \a_out[13] , \a_out[12] , \a_out[11] , 
    \a_out[10] , \a_out[9] , \a_out[8] , \a_out[7] , \a_out[6] , \a_out[5] , \a_out[4] , 
    \a_out[3] , \a_out[2] , \a_out[1] , \a_out[0] }), .b ({\b_out[31] , \b_out[30] , 
    \b_out[29] , \b_out[28] , \b_out[27] , \b_out[26] , \b_out[25] , \b_out[24] , 
    \b_out[23] , \b_out[22] , \b_out[21] , \b_out[20] , \b_out[19] , \b_out[18] , 
    \b_out[17] , \b_out[16] , \b_out[15] , \b_out[14] , \b_out[13] , \b_out[12] , 
    \b_out[11] , \b_out[10] , \b_out[9] , \b_out[8] , \b_out[7] , \b_out[6] , \b_out[5] , 
    \b_out[4] , \b_out[3] , \b_out[2] , \b_out[1] , \b_out[0] }), .rst (rst), .clk_CTS_0_PP_10 (clk));
buffer inRegB (.Q ({\b_out[31] , \b_out[30] , \b_out[29] , \b_out[28] , \b_out[27] , 
    \b_out[26] , \b_out[25] , \b_out[24] , \b_out[23] , \b_out[22] , \b_out[21] , 
    \b_out[20] , \b_out[19] , \b_out[18] , \b_out[17] , \b_out[16] , \b_out[15] , 
    \b_out[14] , \b_out[13] , \b_out[12] , \b_out[11] , \b_out[10] , \b_out[9] , 
    \b_out[8] , \b_out[7] , \b_out[6] , \b_out[5] , \b_out[4] , \b_out[3] , \b_out[2] , 
    \b_out[1] , \b_out[0] }), .D ({CLOCK_slh_n132, CLOCK_slh_n162, CLOCK_slh_n157, 
    CLOCK_slh_n172, CLOCK_slh_n167, b[26], CLOCK_slh_n142, CLOCK_slh_n127, CLOCK_slh_n137, 
    CLOCK_slh_n182, b[21], CLOCK_slh_n227, b[19], CLOCK_slh_n285, CLOCK_slh_n295, 
    CLOCK_slh_n290, CLOCK_slh_n187, b[14], b[13], b[12], b[11], b[10], b[9], b[8], 
    b[7], b[6], b[5], CLOCK_slh_n152, CLOCK_slh_n122, CLOCK_slh_n147, CLOCK_slh_n112, 
    CLOCK_slh_n117}), .en (en), .rst (rst), .clk_CTS_0_PP_0 (CTS_n_tid0_3));
buffer__0_68 inRegA (.Q ({\a_out[31] , \a_out[30] , \a_out[29] , \a_out[28] , \a_out[27] , 
    \a_out[26] , \a_out[25] , \a_out[24] , \a_out[23] , \a_out[22] , \a_out[21] , 
    \a_out[20] , \a_out[19] , \a_out[18] , \a_out[17] , \a_out[16] , \a_out[15] , 
    \a_out[14] , \a_out[13] , \a_out[12] , \a_out[11] , \a_out[10] , \a_out[9] , 
    \a_out[8] , \a_out[7] , \a_out[6] , \a_out[5] , \a_out[4] , \a_out[3] , \a_out[2] , 
    \a_out[1] , \a_out[0] }), .D ({a[31], a[30], a[29], a[28], a[27], a[26], a[25], 
    a[24], a[23], a[22], CLOCK_slh_n232, a[20], CLOCK_slh_n247, CLOCK_slh_n262, CLOCK_slh_n242, 
    CLOCK_slh_n257, CLOCK_slh_n280, CLOCK_slh_n237, a[13], a[12], a[11], a[10], a[9], 
    a[8], CLOCK_slh_n252, CLOCK_slh_n197, CLOCK_slh_n271, CLOCK_slh_n210, CLOCK_slh_n177, 
    CLOCK_slh_n192, a[1], a[0]}), .en (en), .rst (rst), .clk_CTS_0_PP_0 (CTS_n_tid0_3));
CLKBUF_X1 CLOCK_slh__c30 (.Z (CLOCK_slh_n112), .A (b[1]));
CLKBUF_X1 CLOCK_slh__c32 (.Z (CLOCK_slh_n117), .A (b[0]));
CLKBUF_X1 CLOCK_slh__c34 (.Z (CLOCK_slh_n122), .A (b[3]));
CLKBUF_X1 CLOCK_slh__c36 (.Z (CLOCK_slh_n127), .A (b[24]));
CLKBUF_X1 CLOCK_slh__c38 (.Z (CLOCK_slh_n132), .A (b[31]));
CLKBUF_X1 CLOCK_slh__c40 (.Z (CLOCK_slh_n137), .A (b[23]));
CLKBUF_X1 CLOCK_slh__c42 (.Z (CLOCK_slh_n142), .A (b[25]));
CLKBUF_X1 CLOCK_slh__c44 (.Z (CLOCK_slh_n147), .A (b[2]));
CLKBUF_X1 CLOCK_slh__c46 (.Z (CLOCK_slh_n152), .A (b[4]));
CLKBUF_X1 CLOCK_slh__c48 (.Z (CLOCK_slh_n157), .A (b[29]));
CLKBUF_X1 CLOCK_slh__c50 (.Z (CLOCK_slh_n162), .A (b[30]));
CLKBUF_X1 CLOCK_slh__c52 (.Z (CLOCK_slh_n167), .A (b[27]));
CLKBUF_X1 CLOCK_slh__c54 (.Z (CLOCK_slh_n172), .A (b[28]));
CLKBUF_X1 CLOCK_slh__c56 (.Z (CLOCK_slh_n177), .A (a[3]));
CLKBUF_X1 CLOCK_slh__c58 (.Z (CLOCK_slh_n182), .A (b[22]));
CLKBUF_X1 CLOCK_slh__c60 (.Z (CLOCK_slh_n187), .A (b[15]));
CLKBUF_X1 CLOCK_slh__c62 (.Z (CLOCK_slh_n192), .A (a[2]));
CLKBUF_X1 CLOCK_slh__c64 (.Z (CLOCK_slh_n197), .A (a[6]));
CLKBUF_X1 CLOCK_slh__c70 (.Z (CLOCK_slh_n210), .A (a[4]));
CLKBUF_X1 CLOCK_slh__c78 (.Z (CLOCK_slh_n227), .A (b[20]));
CLKBUF_X1 CLOCK_slh__c80 (.Z (CLOCK_slh_n232), .A (a[21]));
CLKBUF_X1 CLOCK_slh__c82 (.Z (CLOCK_slh_n237), .A (a[14]));
CLKBUF_X1 CLOCK_slh__c84 (.Z (CLOCK_slh_n242), .A (a[17]));
CLKBUF_X1 CLOCK_slh__c86 (.Z (CLOCK_slh_n247), .A (a[19]));
CLKBUF_X1 CLOCK_slh__c88 (.Z (CLOCK_slh_n252), .A (a[7]));
CLKBUF_X1 CLOCK_slh__c90 (.Z (CLOCK_slh_n257), .A (a[16]));
CLKBUF_X1 CLOCK_slh__c92 (.Z (CLOCK_slh_n262), .A (a[18]));
CLKBUF_X1 CLOCK_slh__c96 (.Z (CLOCK_slh_n271), .A (a[5]));
CLKBUF_X1 CLOCK_slh__c100 (.Z (CLOCK_slh_n280), .A (a[15]));
CLKBUF_X1 CLOCK_slh__c102 (.Z (CLOCK_slh_n285), .A (b[18]));
CLKBUF_X1 CLOCK_slh__c104 (.Z (CLOCK_slh_n290), .A (b[16]));
CLKBUF_X1 CLOCK_slh__c106 (.Z (CLOCK_slh_n295), .A (b[17]));

endmodule //simpleMultiplier


