/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Dec 27 13:40:25 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3548166540 */

module CSA__1_2(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;

   AND2_X1 i_0_0 (.A1(in2[1]), .A2(in1[1]), .ZN(c[2]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[3]));
   OAI21_X1 i_0_2 (.A(in2[2]), .B1(in3[2]), .B2(in1[2]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[2]), .A2(in1[2]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[4]));
   OAI21_X1 i_0_5 (.A(in2[3]), .B1(in3[3]), .B2(in1[3]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[3]), .A2(in1[3]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[5]));
   OAI21_X1 i_0_8 (.A(in2[4]), .B1(in3[4]), .B2(in1[4]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[4]), .A2(in1[4]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[6]));
   OAI21_X1 i_0_11 (.A(in2[5]), .B1(in3[5]), .B2(in1[5]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[5]), .A2(in1[5]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[7]));
   OAI21_X1 i_0_14 (.A(in2[6]), .B1(in3[6]), .B2(in1[6]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[6]), .A2(in1[6]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[8]));
   OAI21_X1 i_0_17 (.A(in2[7]), .B1(in3[7]), .B2(in1[7]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[7]), .A2(in1[7]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[9]));
   OAI21_X1 i_0_20 (.A(in2[8]), .B1(in3[8]), .B2(in1[8]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[8]), .A2(in1[8]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[10]));
   OAI21_X1 i_0_23 (.A(in2[9]), .B1(in3[9]), .B2(in1[9]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[9]), .A2(in1[9]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[11]));
   OAI21_X1 i_0_26 (.A(in2[10]), .B1(in3[10]), .B2(in1[10]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[10]), .A2(in1[10]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[12]));
   OAI21_X1 i_0_29 (.A(in2[11]), .B1(in3[11]), .B2(in1[11]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[11]), .A2(in1[11]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[13]));
   OAI21_X1 i_0_32 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[14]));
   OAI21_X1 i_0_35 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[15]));
   OAI21_X1 i_0_38 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[16]));
   OAI21_X1 i_0_41 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[17]));
   OAI21_X1 i_0_44 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[18]));
   OAI21_X1 i_0_47 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[19]));
   OAI21_X1 i_0_50 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[20]));
   OAI21_X1 i_0_53 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[21]));
   OAI21_X1 i_0_56 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[22]));
   OAI21_X1 i_0_59 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[23]));
   OAI21_X1 i_0_62 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[24]));
   OAI21_X1 i_0_65 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[25]));
   OAI21_X1 i_0_68 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[26]));
   OAI21_X1 i_0_71 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[27]));
   OAI21_X1 i_0_74 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[28]));
   OAI21_X1 i_0_77 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[29]));
   OAI21_X1 i_0_80 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[30]));
   OAI21_X1 i_0_83 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[31]));
   OAI21_X1 i_0_86 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[32]));
   OAI21_X1 i_0_89 (.A(in2[31]), .B1(in3[31]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[31]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_62), .A2(n_0_60), .ZN(c[33]));
   OAI21_X1 i_0_92 (.A(in3[32]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(c[63]));
   OAI21_X1 i_0_94 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   XOR2_X1 i_0_96 (.A(in2[1]), .B(in1[1]), .Z(sum[1]));
   XNOR2_X1 i_0_97 (.A(in2[2]), .B(n_0_63), .ZN(sum[2]));
   XNOR2_X1 i_0_98 (.A(in3[2]), .B(in1[2]), .ZN(n_0_63));
   XNOR2_X1 i_0_99 (.A(in2[3]), .B(n_0_64), .ZN(sum[3]));
   XNOR2_X1 i_0_100 (.A(in3[3]), .B(in1[3]), .ZN(n_0_64));
   XNOR2_X1 i_0_101 (.A(in2[4]), .B(n_0_65), .ZN(sum[4]));
   XNOR2_X1 i_0_102 (.A(in3[4]), .B(in1[4]), .ZN(n_0_65));
   XNOR2_X1 i_0_103 (.A(in2[5]), .B(n_0_66), .ZN(sum[5]));
   XNOR2_X1 i_0_104 (.A(in3[5]), .B(in1[5]), .ZN(n_0_66));
   XNOR2_X1 i_0_105 (.A(in2[6]), .B(n_0_67), .ZN(sum[6]));
   XNOR2_X1 i_0_106 (.A(in3[6]), .B(in1[6]), .ZN(n_0_67));
   XNOR2_X1 i_0_107 (.A(in2[7]), .B(n_0_68), .ZN(sum[7]));
   XNOR2_X1 i_0_108 (.A(in3[7]), .B(in1[7]), .ZN(n_0_68));
   XNOR2_X1 i_0_109 (.A(in2[8]), .B(n_0_69), .ZN(sum[8]));
   XNOR2_X1 i_0_110 (.A(in3[8]), .B(in1[8]), .ZN(n_0_69));
   XNOR2_X1 i_0_111 (.A(in2[9]), .B(n_0_70), .ZN(sum[9]));
   XNOR2_X1 i_0_112 (.A(in3[9]), .B(in1[9]), .ZN(n_0_70));
   XNOR2_X1 i_0_113 (.A(in2[10]), .B(n_0_71), .ZN(sum[10]));
   XNOR2_X1 i_0_114 (.A(in3[10]), .B(in1[10]), .ZN(n_0_71));
   XNOR2_X1 i_0_115 (.A(in2[11]), .B(n_0_72), .ZN(sum[11]));
   XNOR2_X1 i_0_116 (.A(in3[11]), .B(in1[11]), .ZN(n_0_72));
   XNOR2_X1 i_0_117 (.A(in2[12]), .B(n_0_73), .ZN(sum[12]));
   XNOR2_X1 i_0_118 (.A(in3[12]), .B(in1[12]), .ZN(n_0_73));
   XNOR2_X1 i_0_119 (.A(in2[13]), .B(n_0_74), .ZN(sum[13]));
   XNOR2_X1 i_0_120 (.A(in3[13]), .B(in1[13]), .ZN(n_0_74));
   XNOR2_X1 i_0_121 (.A(in2[14]), .B(n_0_75), .ZN(sum[14]));
   XNOR2_X1 i_0_122 (.A(in3[14]), .B(in1[14]), .ZN(n_0_75));
   XNOR2_X1 i_0_123 (.A(in2[15]), .B(n_0_76), .ZN(sum[15]));
   XNOR2_X1 i_0_124 (.A(in3[15]), .B(in1[15]), .ZN(n_0_76));
   XNOR2_X1 i_0_125 (.A(in2[16]), .B(n_0_77), .ZN(sum[16]));
   XNOR2_X1 i_0_126 (.A(in3[16]), .B(in1[16]), .ZN(n_0_77));
   XNOR2_X1 i_0_127 (.A(in2[17]), .B(n_0_78), .ZN(sum[17]));
   XNOR2_X1 i_0_128 (.A(in3[17]), .B(in1[17]), .ZN(n_0_78));
   XNOR2_X1 i_0_129 (.A(in2[18]), .B(n_0_79), .ZN(sum[18]));
   XNOR2_X1 i_0_130 (.A(in3[18]), .B(in1[18]), .ZN(n_0_79));
   XNOR2_X1 i_0_131 (.A(in2[19]), .B(n_0_80), .ZN(sum[19]));
   XNOR2_X1 i_0_132 (.A(in3[19]), .B(in1[19]), .ZN(n_0_80));
   XNOR2_X1 i_0_133 (.A(in2[20]), .B(n_0_81), .ZN(sum[20]));
   XNOR2_X1 i_0_134 (.A(in3[20]), .B(in1[20]), .ZN(n_0_81));
   XNOR2_X1 i_0_135 (.A(in2[21]), .B(n_0_82), .ZN(sum[21]));
   XNOR2_X1 i_0_136 (.A(in3[21]), .B(in1[21]), .ZN(n_0_82));
   XNOR2_X1 i_0_137 (.A(in2[22]), .B(n_0_83), .ZN(sum[22]));
   XNOR2_X1 i_0_138 (.A(in3[22]), .B(in1[22]), .ZN(n_0_83));
   XNOR2_X1 i_0_139 (.A(in2[23]), .B(n_0_84), .ZN(sum[23]));
   XNOR2_X1 i_0_140 (.A(in3[23]), .B(in1[23]), .ZN(n_0_84));
   XNOR2_X1 i_0_141 (.A(in2[24]), .B(n_0_85), .ZN(sum[24]));
   XNOR2_X1 i_0_142 (.A(in3[24]), .B(in1[24]), .ZN(n_0_85));
   XNOR2_X1 i_0_143 (.A(in2[25]), .B(n_0_86), .ZN(sum[25]));
   XNOR2_X1 i_0_144 (.A(in3[25]), .B(in1[25]), .ZN(n_0_86));
   XNOR2_X1 i_0_145 (.A(in2[26]), .B(n_0_87), .ZN(sum[26]));
   XNOR2_X1 i_0_146 (.A(in3[26]), .B(in1[26]), .ZN(n_0_87));
   XNOR2_X1 i_0_147 (.A(in2[27]), .B(n_0_88), .ZN(sum[27]));
   XNOR2_X1 i_0_148 (.A(in3[27]), .B(in1[27]), .ZN(n_0_88));
   XNOR2_X1 i_0_149 (.A(in2[28]), .B(n_0_89), .ZN(sum[28]));
   XNOR2_X1 i_0_150 (.A(in3[28]), .B(in1[28]), .ZN(n_0_89));
   XNOR2_X1 i_0_151 (.A(in2[29]), .B(n_0_90), .ZN(sum[29]));
   XNOR2_X1 i_0_152 (.A(in3[29]), .B(in1[29]), .ZN(n_0_90));
   XNOR2_X1 i_0_153 (.A(in2[30]), .B(n_0_91), .ZN(sum[30]));
   XNOR2_X1 i_0_154 (.A(in3[30]), .B(in1[30]), .ZN(n_0_91));
   XNOR2_X1 i_0_155 (.A(in2[31]), .B(n_0_92), .ZN(sum[31]));
   XNOR2_X1 i_0_156 (.A(in3[31]), .B(in1[63]), .ZN(n_0_92));
   XOR2_X1 i_0_157 (.A(in3[32]), .B(n_0_93), .Z(sum[32]));
   INV_X1 i_0_158 (.A(n_0_94), .ZN(n_0_93));
   NAND2_X1 i_0_159 (.A1(n_0_99), .A2(n_0_98), .ZN(n_0_94));
   NOR2_X1 i_0_160 (.A1(n_0_95), .A2(n_0_97), .ZN(sum[63]));
   INV_X1 i_0_161 (.A(n_0_96), .ZN(n_0_95));
   NAND3_X1 i_0_162 (.A1(n_0_99), .A2(in3[63]), .A3(n_0_98), .ZN(n_0_96));
   AOI21_X1 i_0_163 (.A(in3[63]), .B1(n_0_99), .B2(n_0_98), .ZN(n_0_97));
   NAND2_X1 i_0_164 (.A1(in1[63]), .A2(in2[63]), .ZN(n_0_98));
   NAND2_X1 i_0_165 (.A1(n_0_100), .A2(n_0_101), .ZN(n_0_99));
   INV_X1 i_0_166 (.A(in1[63]), .ZN(n_0_100));
   INV_X1 i_0_167 (.A(in2[63]), .ZN(n_0_101));
endmodule

module CSA__1_5(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;

   AND2_X1 i_0_0 (.A1(in2[4]), .A2(in1[4]), .ZN(c[5]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[6]));
   OAI21_X1 i_0_2 (.A(in2[5]), .B1(in3[5]), .B2(in1[5]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[5]), .A2(in1[5]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[7]));
   OAI21_X1 i_0_5 (.A(in2[6]), .B1(in3[6]), .B2(in1[6]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[6]), .A2(in1[6]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[8]));
   OAI21_X1 i_0_8 (.A(in2[7]), .B1(in3[7]), .B2(in1[7]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[7]), .A2(in1[7]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[9]));
   OAI21_X1 i_0_11 (.A(in2[8]), .B1(in3[8]), .B2(in1[8]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[8]), .A2(in1[8]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[10]));
   OAI21_X1 i_0_14 (.A(in2[9]), .B1(in3[9]), .B2(in1[9]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[9]), .A2(in1[9]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[11]));
   OAI21_X1 i_0_17 (.A(in2[10]), .B1(in3[10]), .B2(in1[10]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[10]), .A2(in1[10]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[12]));
   OAI21_X1 i_0_20 (.A(in2[11]), .B1(in3[11]), .B2(in1[11]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[11]), .A2(in1[11]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[13]));
   OAI21_X1 i_0_23 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[14]));
   OAI21_X1 i_0_26 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[15]));
   OAI21_X1 i_0_29 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[16]));
   OAI21_X1 i_0_32 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[17]));
   OAI21_X1 i_0_35 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[18]));
   OAI21_X1 i_0_38 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[19]));
   OAI21_X1 i_0_41 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[20]));
   OAI21_X1 i_0_44 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[21]));
   OAI21_X1 i_0_47 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[22]));
   OAI21_X1 i_0_50 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[23]));
   OAI21_X1 i_0_53 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[24]));
   OAI21_X1 i_0_56 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[25]));
   OAI21_X1 i_0_59 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[26]));
   OAI21_X1 i_0_62 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[27]));
   OAI21_X1 i_0_65 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[28]));
   OAI21_X1 i_0_68 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[29]));
   OAI21_X1 i_0_71 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[30]));
   OAI21_X1 i_0_74 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[31]));
   OAI21_X1 i_0_77 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[32]));
   OAI21_X1 i_0_80 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[33]));
   OAI21_X1 i_0_83 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[34]));
   OAI21_X1 i_0_86 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[35]));
   OAI21_X1 i_0_89 (.A(in2[34]), .B1(in3[34]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[34]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_62), .A2(n_0_60), .ZN(c[36]));
   OAI21_X1 i_0_92 (.A(in3[35]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(c[63]));
   OAI21_X1 i_0_94 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   XOR2_X1 i_0_96 (.A(in2[4]), .B(in1[4]), .Z(sum[4]));
   XNOR2_X1 i_0_97 (.A(in2[5]), .B(n_0_63), .ZN(sum[5]));
   XNOR2_X1 i_0_98 (.A(in3[5]), .B(in1[5]), .ZN(n_0_63));
   XNOR2_X1 i_0_99 (.A(in2[6]), .B(n_0_64), .ZN(sum[6]));
   XNOR2_X1 i_0_100 (.A(in3[6]), .B(in1[6]), .ZN(n_0_64));
   XNOR2_X1 i_0_101 (.A(in2[7]), .B(n_0_65), .ZN(sum[7]));
   XNOR2_X1 i_0_102 (.A(in3[7]), .B(in1[7]), .ZN(n_0_65));
   XNOR2_X1 i_0_103 (.A(in2[8]), .B(n_0_66), .ZN(sum[8]));
   XNOR2_X1 i_0_104 (.A(in3[8]), .B(in1[8]), .ZN(n_0_66));
   XNOR2_X1 i_0_105 (.A(in2[9]), .B(n_0_67), .ZN(sum[9]));
   XNOR2_X1 i_0_106 (.A(in3[9]), .B(in1[9]), .ZN(n_0_67));
   XNOR2_X1 i_0_107 (.A(in2[10]), .B(n_0_68), .ZN(sum[10]));
   XNOR2_X1 i_0_108 (.A(in3[10]), .B(in1[10]), .ZN(n_0_68));
   XNOR2_X1 i_0_109 (.A(in2[11]), .B(n_0_69), .ZN(sum[11]));
   XNOR2_X1 i_0_110 (.A(in3[11]), .B(in1[11]), .ZN(n_0_69));
   XNOR2_X1 i_0_111 (.A(in2[12]), .B(n_0_70), .ZN(sum[12]));
   XNOR2_X1 i_0_112 (.A(in3[12]), .B(in1[12]), .ZN(n_0_70));
   XNOR2_X1 i_0_113 (.A(in2[13]), .B(n_0_71), .ZN(sum[13]));
   XNOR2_X1 i_0_114 (.A(in3[13]), .B(in1[13]), .ZN(n_0_71));
   XNOR2_X1 i_0_115 (.A(in2[14]), .B(n_0_72), .ZN(sum[14]));
   XNOR2_X1 i_0_116 (.A(in3[14]), .B(in1[14]), .ZN(n_0_72));
   XNOR2_X1 i_0_117 (.A(in2[15]), .B(n_0_73), .ZN(sum[15]));
   XNOR2_X1 i_0_118 (.A(in3[15]), .B(in1[15]), .ZN(n_0_73));
   XNOR2_X1 i_0_119 (.A(in2[16]), .B(n_0_74), .ZN(sum[16]));
   XNOR2_X1 i_0_120 (.A(in3[16]), .B(in1[16]), .ZN(n_0_74));
   XNOR2_X1 i_0_121 (.A(in2[17]), .B(n_0_75), .ZN(sum[17]));
   XNOR2_X1 i_0_122 (.A(in3[17]), .B(in1[17]), .ZN(n_0_75));
   XNOR2_X1 i_0_123 (.A(in2[18]), .B(n_0_76), .ZN(sum[18]));
   XNOR2_X1 i_0_124 (.A(in3[18]), .B(in1[18]), .ZN(n_0_76));
   XNOR2_X1 i_0_125 (.A(in2[19]), .B(n_0_77), .ZN(sum[19]));
   XNOR2_X1 i_0_126 (.A(in3[19]), .B(in1[19]), .ZN(n_0_77));
   XNOR2_X1 i_0_127 (.A(in2[20]), .B(n_0_78), .ZN(sum[20]));
   XNOR2_X1 i_0_128 (.A(in3[20]), .B(in1[20]), .ZN(n_0_78));
   XNOR2_X1 i_0_129 (.A(in2[21]), .B(n_0_79), .ZN(sum[21]));
   XNOR2_X1 i_0_130 (.A(in3[21]), .B(in1[21]), .ZN(n_0_79));
   XNOR2_X1 i_0_131 (.A(in2[22]), .B(n_0_80), .ZN(sum[22]));
   XNOR2_X1 i_0_132 (.A(in3[22]), .B(in1[22]), .ZN(n_0_80));
   XNOR2_X1 i_0_133 (.A(in2[23]), .B(n_0_81), .ZN(sum[23]));
   XNOR2_X1 i_0_134 (.A(in3[23]), .B(in1[23]), .ZN(n_0_81));
   XNOR2_X1 i_0_135 (.A(in2[24]), .B(n_0_82), .ZN(sum[24]));
   XNOR2_X1 i_0_136 (.A(in3[24]), .B(in1[24]), .ZN(n_0_82));
   XNOR2_X1 i_0_137 (.A(in2[25]), .B(n_0_83), .ZN(sum[25]));
   XNOR2_X1 i_0_138 (.A(in3[25]), .B(in1[25]), .ZN(n_0_83));
   XNOR2_X1 i_0_139 (.A(in2[26]), .B(n_0_84), .ZN(sum[26]));
   XNOR2_X1 i_0_140 (.A(in3[26]), .B(in1[26]), .ZN(n_0_84));
   XNOR2_X1 i_0_141 (.A(in2[27]), .B(n_0_85), .ZN(sum[27]));
   XNOR2_X1 i_0_142 (.A(in3[27]), .B(in1[27]), .ZN(n_0_85));
   XNOR2_X1 i_0_143 (.A(in2[28]), .B(n_0_86), .ZN(sum[28]));
   XNOR2_X1 i_0_144 (.A(in3[28]), .B(in1[28]), .ZN(n_0_86));
   XNOR2_X1 i_0_145 (.A(in2[29]), .B(n_0_87), .ZN(sum[29]));
   XNOR2_X1 i_0_146 (.A(in3[29]), .B(in1[29]), .ZN(n_0_87));
   XNOR2_X1 i_0_147 (.A(in2[30]), .B(n_0_88), .ZN(sum[30]));
   XNOR2_X1 i_0_148 (.A(in3[30]), .B(in1[30]), .ZN(n_0_88));
   XNOR2_X1 i_0_149 (.A(in2[31]), .B(n_0_89), .ZN(sum[31]));
   XNOR2_X1 i_0_150 (.A(in3[31]), .B(in1[31]), .ZN(n_0_89));
   XNOR2_X1 i_0_151 (.A(in2[32]), .B(n_0_90), .ZN(sum[32]));
   XNOR2_X1 i_0_152 (.A(in3[32]), .B(in1[32]), .ZN(n_0_90));
   XNOR2_X1 i_0_153 (.A(in2[33]), .B(n_0_91), .ZN(sum[33]));
   XNOR2_X1 i_0_154 (.A(in3[33]), .B(in1[33]), .ZN(n_0_91));
   XNOR2_X1 i_0_155 (.A(in2[34]), .B(n_0_92), .ZN(sum[34]));
   XNOR2_X1 i_0_156 (.A(in3[34]), .B(in1[63]), .ZN(n_0_92));
   XOR2_X1 i_0_157 (.A(in3[35]), .B(n_0_93), .Z(sum[35]));
   INV_X1 i_0_158 (.A(n_0_94), .ZN(n_0_93));
   NAND2_X1 i_0_159 (.A1(n_0_99), .A2(n_0_98), .ZN(n_0_94));
   NOR2_X1 i_0_160 (.A1(n_0_95), .A2(n_0_97), .ZN(sum[63]));
   INV_X1 i_0_161 (.A(n_0_96), .ZN(n_0_95));
   NAND3_X1 i_0_162 (.A1(n_0_99), .A2(in3[63]), .A3(n_0_98), .ZN(n_0_96));
   AOI21_X1 i_0_163 (.A(in3[63]), .B1(n_0_99), .B2(n_0_98), .ZN(n_0_97));
   NAND2_X1 i_0_164 (.A1(in1[63]), .A2(in2[63]), .ZN(n_0_98));
   NAND2_X1 i_0_165 (.A1(n_0_100), .A2(n_0_101), .ZN(n_0_99));
   INV_X1 i_0_166 (.A(in1[63]), .ZN(n_0_100));
   INV_X1 i_0_167 (.A(in2[63]), .ZN(n_0_101));
endmodule

module CSA__1_8(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;

   AND2_X1 i_0_0 (.A1(in2[2]), .A2(in1[2]), .ZN(c[3]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[4]));
   OAI21_X1 i_0_2 (.A(in2[3]), .B1(in3[3]), .B2(in1[3]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[3]), .A2(in1[3]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[5]));
   OAI21_X1 i_0_5 (.A(in2[4]), .B1(in3[4]), .B2(in1[4]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[4]), .A2(in1[4]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[6]));
   OAI21_X1 i_0_8 (.A(in2[5]), .B1(in3[5]), .B2(in1[5]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[5]), .A2(in1[5]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[7]));
   OAI21_X1 i_0_11 (.A(in2[6]), .B1(in3[6]), .B2(in1[6]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[6]), .A2(in1[6]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[8]));
   OAI21_X1 i_0_14 (.A(in2[7]), .B1(in3[7]), .B2(in1[7]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[7]), .A2(in1[7]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[9]));
   OAI21_X1 i_0_17 (.A(in2[8]), .B1(in3[8]), .B2(in1[8]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[8]), .A2(in1[8]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[10]));
   OAI21_X1 i_0_20 (.A(in2[9]), .B1(in3[9]), .B2(in1[9]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[9]), .A2(in1[9]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[11]));
   OAI21_X1 i_0_23 (.A(in2[10]), .B1(in3[10]), .B2(in1[10]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[10]), .A2(in1[10]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[12]));
   OAI21_X1 i_0_26 (.A(in2[11]), .B1(in3[11]), .B2(in1[11]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[11]), .A2(in1[11]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[13]));
   OAI21_X1 i_0_29 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[14]));
   OAI21_X1 i_0_32 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[15]));
   OAI21_X1 i_0_35 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[16]));
   OAI21_X1 i_0_38 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[17]));
   OAI21_X1 i_0_41 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[18]));
   OAI21_X1 i_0_44 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[19]));
   OAI21_X1 i_0_47 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[20]));
   OAI21_X1 i_0_50 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[21]));
   OAI21_X1 i_0_53 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[22]));
   OAI21_X1 i_0_56 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[23]));
   OAI21_X1 i_0_59 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[24]));
   OAI21_X1 i_0_62 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[25]));
   OAI21_X1 i_0_65 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[26]));
   OAI21_X1 i_0_68 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[27]));
   OAI21_X1 i_0_71 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[28]));
   OAI21_X1 i_0_74 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[29]));
   OAI21_X1 i_0_77 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[30]));
   OAI21_X1 i_0_80 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[31]));
   OAI21_X1 i_0_83 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[32]));
   OAI21_X1 i_0_86 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[33]));
   OAI21_X1 i_0_89 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_61), .A2(n_0_60), .ZN(c[34]));
   OAI21_X1 i_0_92 (.A(in2[33]), .B1(in3[33]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(in3[33]), .A2(in1[63]), .ZN(n_0_61));
   AOI21_X1 i_0_94 (.A(n_0_63), .B1(n_0_62), .B2(n_0_96), .ZN(c[35]));
   AOI21_X1 i_0_95 (.A(n_0_63), .B1(n_0_62), .B2(n_0_97), .ZN(c[36]));
   AOI21_X1 i_0_96 (.A(n_0_63), .B1(n_0_62), .B2(n_0_98), .ZN(c[63]));
   NAND2_X1 i_0_97 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   NOR2_X1 i_0_98 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_63));
   XOR2_X1 i_0_99 (.A(in2[2]), .B(in1[2]), .Z(sum[2]));
   XNOR2_X1 i_0_100 (.A(in2[3]), .B(n_0_64), .ZN(sum[3]));
   XNOR2_X1 i_0_101 (.A(in3[3]), .B(in1[3]), .ZN(n_0_64));
   XNOR2_X1 i_0_102 (.A(in2[4]), .B(n_0_65), .ZN(sum[4]));
   XNOR2_X1 i_0_103 (.A(in3[4]), .B(in1[4]), .ZN(n_0_65));
   XNOR2_X1 i_0_104 (.A(in2[5]), .B(n_0_66), .ZN(sum[5]));
   XNOR2_X1 i_0_105 (.A(in3[5]), .B(in1[5]), .ZN(n_0_66));
   XNOR2_X1 i_0_106 (.A(in2[6]), .B(n_0_67), .ZN(sum[6]));
   XNOR2_X1 i_0_107 (.A(in3[6]), .B(in1[6]), .ZN(n_0_67));
   XNOR2_X1 i_0_108 (.A(in2[7]), .B(n_0_68), .ZN(sum[7]));
   XNOR2_X1 i_0_109 (.A(in3[7]), .B(in1[7]), .ZN(n_0_68));
   XNOR2_X1 i_0_110 (.A(in2[8]), .B(n_0_69), .ZN(sum[8]));
   XNOR2_X1 i_0_111 (.A(in3[8]), .B(in1[8]), .ZN(n_0_69));
   XNOR2_X1 i_0_112 (.A(in2[9]), .B(n_0_70), .ZN(sum[9]));
   XNOR2_X1 i_0_113 (.A(in3[9]), .B(in1[9]), .ZN(n_0_70));
   XNOR2_X1 i_0_114 (.A(in2[10]), .B(n_0_71), .ZN(sum[10]));
   XNOR2_X1 i_0_115 (.A(in3[10]), .B(in1[10]), .ZN(n_0_71));
   XNOR2_X1 i_0_116 (.A(in2[11]), .B(n_0_72), .ZN(sum[11]));
   XNOR2_X1 i_0_117 (.A(in3[11]), .B(in1[11]), .ZN(n_0_72));
   XNOR2_X1 i_0_118 (.A(in2[12]), .B(n_0_73), .ZN(sum[12]));
   XNOR2_X1 i_0_119 (.A(in3[12]), .B(in1[12]), .ZN(n_0_73));
   XNOR2_X1 i_0_120 (.A(in2[13]), .B(n_0_74), .ZN(sum[13]));
   XNOR2_X1 i_0_121 (.A(in3[13]), .B(in1[13]), .ZN(n_0_74));
   XNOR2_X1 i_0_122 (.A(in2[14]), .B(n_0_75), .ZN(sum[14]));
   XNOR2_X1 i_0_123 (.A(in3[14]), .B(in1[14]), .ZN(n_0_75));
   XNOR2_X1 i_0_124 (.A(in2[15]), .B(n_0_76), .ZN(sum[15]));
   XNOR2_X1 i_0_125 (.A(in3[15]), .B(in1[15]), .ZN(n_0_76));
   XNOR2_X1 i_0_126 (.A(in2[16]), .B(n_0_77), .ZN(sum[16]));
   XNOR2_X1 i_0_127 (.A(in3[16]), .B(in1[16]), .ZN(n_0_77));
   XNOR2_X1 i_0_128 (.A(in2[17]), .B(n_0_78), .ZN(sum[17]));
   XNOR2_X1 i_0_129 (.A(in3[17]), .B(in1[17]), .ZN(n_0_78));
   XNOR2_X1 i_0_130 (.A(in2[18]), .B(n_0_79), .ZN(sum[18]));
   XNOR2_X1 i_0_131 (.A(in3[18]), .B(in1[18]), .ZN(n_0_79));
   XNOR2_X1 i_0_132 (.A(in2[19]), .B(n_0_80), .ZN(sum[19]));
   XNOR2_X1 i_0_133 (.A(in3[19]), .B(in1[19]), .ZN(n_0_80));
   XNOR2_X1 i_0_134 (.A(in2[20]), .B(n_0_81), .ZN(sum[20]));
   XNOR2_X1 i_0_135 (.A(in3[20]), .B(in1[20]), .ZN(n_0_81));
   XNOR2_X1 i_0_136 (.A(in2[21]), .B(n_0_82), .ZN(sum[21]));
   XNOR2_X1 i_0_137 (.A(in3[21]), .B(in1[21]), .ZN(n_0_82));
   XNOR2_X1 i_0_138 (.A(in2[22]), .B(n_0_83), .ZN(sum[22]));
   XNOR2_X1 i_0_139 (.A(in3[22]), .B(in1[22]), .ZN(n_0_83));
   XNOR2_X1 i_0_140 (.A(in2[23]), .B(n_0_84), .ZN(sum[23]));
   XNOR2_X1 i_0_141 (.A(in3[23]), .B(in1[23]), .ZN(n_0_84));
   XNOR2_X1 i_0_142 (.A(in2[24]), .B(n_0_85), .ZN(sum[24]));
   XNOR2_X1 i_0_143 (.A(in3[24]), .B(in1[24]), .ZN(n_0_85));
   XNOR2_X1 i_0_144 (.A(in2[25]), .B(n_0_86), .ZN(sum[25]));
   XNOR2_X1 i_0_145 (.A(in3[25]), .B(in1[25]), .ZN(n_0_86));
   XNOR2_X1 i_0_146 (.A(in2[26]), .B(n_0_87), .ZN(sum[26]));
   XNOR2_X1 i_0_147 (.A(in3[26]), .B(in1[26]), .ZN(n_0_87));
   XNOR2_X1 i_0_148 (.A(in2[27]), .B(n_0_88), .ZN(sum[27]));
   XNOR2_X1 i_0_149 (.A(in3[27]), .B(in1[27]), .ZN(n_0_88));
   XNOR2_X1 i_0_150 (.A(in2[28]), .B(n_0_89), .ZN(sum[28]));
   XNOR2_X1 i_0_151 (.A(in3[28]), .B(in1[28]), .ZN(n_0_89));
   XNOR2_X1 i_0_152 (.A(in2[29]), .B(n_0_90), .ZN(sum[29]));
   XNOR2_X1 i_0_153 (.A(in3[29]), .B(in1[29]), .ZN(n_0_90));
   XNOR2_X1 i_0_154 (.A(in2[30]), .B(n_0_91), .ZN(sum[30]));
   XNOR2_X1 i_0_155 (.A(in3[30]), .B(in1[30]), .ZN(n_0_91));
   XNOR2_X1 i_0_156 (.A(in2[31]), .B(n_0_92), .ZN(sum[31]));
   XNOR2_X1 i_0_157 (.A(in3[31]), .B(in1[31]), .ZN(n_0_92));
   XNOR2_X1 i_0_158 (.A(in2[32]), .B(n_0_93), .ZN(sum[32]));
   XNOR2_X1 i_0_159 (.A(in3[32]), .B(in1[32]), .ZN(n_0_93));
   XNOR2_X1 i_0_160 (.A(in2[33]), .B(n_0_94), .ZN(sum[33]));
   XNOR2_X1 i_0_161 (.A(in3[33]), .B(in1[63]), .ZN(n_0_94));
   XNOR2_X1 i_0_162 (.A(n_0_96), .B(n_0_95), .ZN(sum[34]));
   XNOR2_X1 i_0_163 (.A(n_0_97), .B(n_0_95), .ZN(sum[35]));
   XNOR2_X1 i_0_164 (.A(n_0_98), .B(n_0_95), .ZN(sum[63]));
   XOR2_X1 i_0_165 (.A(in2[63]), .B(in1[63]), .Z(n_0_95));
   INV_X1 i_0_166 (.A(in3[34]), .ZN(n_0_96));
   INV_X1 i_0_167 (.A(in3[35]), .ZN(n_0_97));
   INV_X1 i_0_168 (.A(in3[63]), .ZN(n_0_98));
endmodule

module CSA__1_11(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;

   AND2_X1 i_0_0 (.A1(in2[7]), .A2(in1[7]), .ZN(c[8]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[9]));
   OAI21_X1 i_0_2 (.A(in2[8]), .B1(in3[8]), .B2(in1[8]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[8]), .A2(in1[8]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[10]));
   OAI21_X1 i_0_5 (.A(in2[9]), .B1(in3[9]), .B2(in1[9]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[9]), .A2(in1[9]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[11]));
   OAI21_X1 i_0_8 (.A(in2[10]), .B1(in3[10]), .B2(in1[10]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[10]), .A2(in1[10]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[12]));
   OAI21_X1 i_0_11 (.A(in2[11]), .B1(in3[11]), .B2(in1[11]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[11]), .A2(in1[11]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[13]));
   OAI21_X1 i_0_14 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[14]));
   OAI21_X1 i_0_17 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[15]));
   OAI21_X1 i_0_20 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[16]));
   OAI21_X1 i_0_23 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[17]));
   OAI21_X1 i_0_26 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[18]));
   OAI21_X1 i_0_29 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[19]));
   OAI21_X1 i_0_32 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[20]));
   OAI21_X1 i_0_35 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[21]));
   OAI21_X1 i_0_38 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[22]));
   OAI21_X1 i_0_41 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[23]));
   OAI21_X1 i_0_44 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[24]));
   OAI21_X1 i_0_47 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[25]));
   OAI21_X1 i_0_50 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[26]));
   OAI21_X1 i_0_53 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[27]));
   OAI21_X1 i_0_56 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[28]));
   OAI21_X1 i_0_59 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[29]));
   OAI21_X1 i_0_62 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[30]));
   OAI21_X1 i_0_65 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[31]));
   OAI21_X1 i_0_68 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[32]));
   OAI21_X1 i_0_71 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[33]));
   OAI21_X1 i_0_74 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[34]));
   OAI21_X1 i_0_77 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[35]));
   OAI21_X1 i_0_80 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[36]));
   OAI21_X1 i_0_83 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[37]));
   OAI21_X1 i_0_86 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[38]));
   OAI21_X1 i_0_89 (.A(in2[37]), .B1(in3[37]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[37]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_62), .A2(n_0_60), .ZN(c[39]));
   OAI21_X1 i_0_92 (.A(in3[38]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(c[63]));
   OAI21_X1 i_0_94 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   XOR2_X1 i_0_96 (.A(in2[7]), .B(in1[7]), .Z(sum[7]));
   XNOR2_X1 i_0_97 (.A(in2[8]), .B(n_0_63), .ZN(sum[8]));
   XNOR2_X1 i_0_98 (.A(in3[8]), .B(in1[8]), .ZN(n_0_63));
   XNOR2_X1 i_0_99 (.A(in2[9]), .B(n_0_64), .ZN(sum[9]));
   XNOR2_X1 i_0_100 (.A(in3[9]), .B(in1[9]), .ZN(n_0_64));
   XNOR2_X1 i_0_101 (.A(in2[10]), .B(n_0_65), .ZN(sum[10]));
   XNOR2_X1 i_0_102 (.A(in3[10]), .B(in1[10]), .ZN(n_0_65));
   XNOR2_X1 i_0_103 (.A(in2[11]), .B(n_0_66), .ZN(sum[11]));
   XNOR2_X1 i_0_104 (.A(in3[11]), .B(in1[11]), .ZN(n_0_66));
   XNOR2_X1 i_0_105 (.A(in2[12]), .B(n_0_67), .ZN(sum[12]));
   XNOR2_X1 i_0_106 (.A(in3[12]), .B(in1[12]), .ZN(n_0_67));
   XNOR2_X1 i_0_107 (.A(in2[13]), .B(n_0_68), .ZN(sum[13]));
   XNOR2_X1 i_0_108 (.A(in3[13]), .B(in1[13]), .ZN(n_0_68));
   XNOR2_X1 i_0_109 (.A(in2[14]), .B(n_0_69), .ZN(sum[14]));
   XNOR2_X1 i_0_110 (.A(in3[14]), .B(in1[14]), .ZN(n_0_69));
   XNOR2_X1 i_0_111 (.A(in2[15]), .B(n_0_70), .ZN(sum[15]));
   XNOR2_X1 i_0_112 (.A(in3[15]), .B(in1[15]), .ZN(n_0_70));
   XNOR2_X1 i_0_113 (.A(in2[16]), .B(n_0_71), .ZN(sum[16]));
   XNOR2_X1 i_0_114 (.A(in3[16]), .B(in1[16]), .ZN(n_0_71));
   XNOR2_X1 i_0_115 (.A(in2[17]), .B(n_0_72), .ZN(sum[17]));
   XNOR2_X1 i_0_116 (.A(in3[17]), .B(in1[17]), .ZN(n_0_72));
   XNOR2_X1 i_0_117 (.A(in2[18]), .B(n_0_73), .ZN(sum[18]));
   XNOR2_X1 i_0_118 (.A(in3[18]), .B(in1[18]), .ZN(n_0_73));
   XNOR2_X1 i_0_119 (.A(in2[19]), .B(n_0_74), .ZN(sum[19]));
   XNOR2_X1 i_0_120 (.A(in3[19]), .B(in1[19]), .ZN(n_0_74));
   XNOR2_X1 i_0_121 (.A(in2[20]), .B(n_0_75), .ZN(sum[20]));
   XNOR2_X1 i_0_122 (.A(in3[20]), .B(in1[20]), .ZN(n_0_75));
   XNOR2_X1 i_0_123 (.A(in2[21]), .B(n_0_76), .ZN(sum[21]));
   XNOR2_X1 i_0_124 (.A(in3[21]), .B(in1[21]), .ZN(n_0_76));
   XNOR2_X1 i_0_125 (.A(in2[22]), .B(n_0_77), .ZN(sum[22]));
   XNOR2_X1 i_0_126 (.A(in3[22]), .B(in1[22]), .ZN(n_0_77));
   XNOR2_X1 i_0_127 (.A(in2[23]), .B(n_0_78), .ZN(sum[23]));
   XNOR2_X1 i_0_128 (.A(in3[23]), .B(in1[23]), .ZN(n_0_78));
   XNOR2_X1 i_0_129 (.A(in2[24]), .B(n_0_79), .ZN(sum[24]));
   XNOR2_X1 i_0_130 (.A(in3[24]), .B(in1[24]), .ZN(n_0_79));
   XNOR2_X1 i_0_131 (.A(in2[25]), .B(n_0_80), .ZN(sum[25]));
   XNOR2_X1 i_0_132 (.A(in3[25]), .B(in1[25]), .ZN(n_0_80));
   XNOR2_X1 i_0_133 (.A(in2[26]), .B(n_0_81), .ZN(sum[26]));
   XNOR2_X1 i_0_134 (.A(in3[26]), .B(in1[26]), .ZN(n_0_81));
   XNOR2_X1 i_0_135 (.A(in2[27]), .B(n_0_82), .ZN(sum[27]));
   XNOR2_X1 i_0_136 (.A(in3[27]), .B(in1[27]), .ZN(n_0_82));
   XNOR2_X1 i_0_137 (.A(in2[28]), .B(n_0_83), .ZN(sum[28]));
   XNOR2_X1 i_0_138 (.A(in3[28]), .B(in1[28]), .ZN(n_0_83));
   XNOR2_X1 i_0_139 (.A(in2[29]), .B(n_0_84), .ZN(sum[29]));
   XNOR2_X1 i_0_140 (.A(in3[29]), .B(in1[29]), .ZN(n_0_84));
   XNOR2_X1 i_0_141 (.A(in2[30]), .B(n_0_85), .ZN(sum[30]));
   XNOR2_X1 i_0_142 (.A(in3[30]), .B(in1[30]), .ZN(n_0_85));
   XNOR2_X1 i_0_143 (.A(in2[31]), .B(n_0_86), .ZN(sum[31]));
   XNOR2_X1 i_0_144 (.A(in3[31]), .B(in1[31]), .ZN(n_0_86));
   XNOR2_X1 i_0_145 (.A(in2[32]), .B(n_0_87), .ZN(sum[32]));
   XNOR2_X1 i_0_146 (.A(in3[32]), .B(in1[32]), .ZN(n_0_87));
   XNOR2_X1 i_0_147 (.A(in2[33]), .B(n_0_88), .ZN(sum[33]));
   XNOR2_X1 i_0_148 (.A(in3[33]), .B(in1[33]), .ZN(n_0_88));
   XNOR2_X1 i_0_149 (.A(in2[34]), .B(n_0_89), .ZN(sum[34]));
   XNOR2_X1 i_0_150 (.A(in3[34]), .B(in1[34]), .ZN(n_0_89));
   XNOR2_X1 i_0_151 (.A(in2[35]), .B(n_0_90), .ZN(sum[35]));
   XNOR2_X1 i_0_152 (.A(in3[35]), .B(in1[35]), .ZN(n_0_90));
   XNOR2_X1 i_0_153 (.A(in2[36]), .B(n_0_91), .ZN(sum[36]));
   XNOR2_X1 i_0_154 (.A(in3[36]), .B(in1[36]), .ZN(n_0_91));
   XNOR2_X1 i_0_155 (.A(in2[37]), .B(n_0_92), .ZN(sum[37]));
   XNOR2_X1 i_0_156 (.A(in3[37]), .B(in1[63]), .ZN(n_0_92));
   XOR2_X1 i_0_157 (.A(in3[38]), .B(n_0_93), .Z(sum[38]));
   XOR2_X1 i_0_158 (.A(in3[63]), .B(n_0_93), .Z(sum[63]));
   XOR2_X1 i_0_159 (.A(in2[63]), .B(in1[63]), .Z(n_0_93));
endmodule

module CSA__1_14(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;

   AND2_X1 i_0_0 (.A1(in2[6]), .A2(in1[6]), .ZN(c[7]));
   AND2_X1 i_0_1 (.A1(in2[7]), .A2(in1[7]), .ZN(c[8]));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_0), .ZN(c[9]));
   OAI21_X1 i_0_3 (.A(in2[8]), .B1(in3[8]), .B2(in1[8]), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(in3[8]), .A2(in1[8]), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .ZN(c[10]));
   OAI21_X1 i_0_6 (.A(in2[9]), .B1(in3[9]), .B2(in1[9]), .ZN(n_0_2));
   NAND2_X1 i_0_7 (.A1(in3[9]), .A2(in1[9]), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_4), .ZN(c[11]));
   OAI21_X1 i_0_9 (.A(in2[10]), .B1(in3[10]), .B2(in1[10]), .ZN(n_0_4));
   NAND2_X1 i_0_10 (.A1(in3[10]), .A2(in1[10]), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(n_0_7), .A2(n_0_6), .ZN(c[12]));
   OAI21_X1 i_0_12 (.A(in2[11]), .B1(in3[11]), .B2(in1[11]), .ZN(n_0_6));
   NAND2_X1 i_0_13 (.A1(in3[11]), .A2(in1[11]), .ZN(n_0_7));
   NAND2_X1 i_0_14 (.A1(n_0_9), .A2(n_0_8), .ZN(c[13]));
   OAI21_X1 i_0_15 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_8));
   NAND2_X1 i_0_16 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_9));
   NAND2_X1 i_0_17 (.A1(n_0_11), .A2(n_0_10), .ZN(c[14]));
   OAI21_X1 i_0_18 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_10));
   NAND2_X1 i_0_19 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_11));
   NAND2_X1 i_0_20 (.A1(n_0_13), .A2(n_0_12), .ZN(c[15]));
   OAI21_X1 i_0_21 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_12));
   NAND2_X1 i_0_22 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_13));
   NAND2_X1 i_0_23 (.A1(n_0_15), .A2(n_0_14), .ZN(c[16]));
   OAI21_X1 i_0_24 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_14));
   NAND2_X1 i_0_25 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_15));
   NAND2_X1 i_0_26 (.A1(n_0_17), .A2(n_0_16), .ZN(c[17]));
   OAI21_X1 i_0_27 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_16));
   NAND2_X1 i_0_28 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_17));
   NAND2_X1 i_0_29 (.A1(n_0_19), .A2(n_0_18), .ZN(c[18]));
   OAI21_X1 i_0_30 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_18));
   NAND2_X1 i_0_31 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_19));
   NAND2_X1 i_0_32 (.A1(n_0_21), .A2(n_0_20), .ZN(c[19]));
   OAI21_X1 i_0_33 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_20));
   NAND2_X1 i_0_34 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_21));
   NAND2_X1 i_0_35 (.A1(n_0_23), .A2(n_0_22), .ZN(c[20]));
   OAI21_X1 i_0_36 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_22));
   NAND2_X1 i_0_37 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_23));
   NAND2_X1 i_0_38 (.A1(n_0_25), .A2(n_0_24), .ZN(c[21]));
   OAI21_X1 i_0_39 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_24));
   NAND2_X1 i_0_40 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_25));
   NAND2_X1 i_0_41 (.A1(n_0_27), .A2(n_0_26), .ZN(c[22]));
   OAI21_X1 i_0_42 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_26));
   NAND2_X1 i_0_43 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_27));
   NAND2_X1 i_0_44 (.A1(n_0_29), .A2(n_0_28), .ZN(c[23]));
   OAI21_X1 i_0_45 (.A(in1[22]), .B1(in3[22]), .B2(in2[22]), .ZN(n_0_28));
   NAND2_X1 i_0_46 (.A1(in2[22]), .A2(in3[22]), .ZN(n_0_29));
   NAND2_X1 i_0_47 (.A1(n_0_31), .A2(n_0_30), .ZN(c[24]));
   OAI21_X1 i_0_48 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_30));
   NAND2_X1 i_0_49 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_31));
   NAND2_X1 i_0_50 (.A1(n_0_33), .A2(n_0_32), .ZN(c[25]));
   OAI21_X1 i_0_51 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_32));
   NAND2_X1 i_0_52 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_33));
   NAND2_X1 i_0_53 (.A1(n_0_35), .A2(n_0_34), .ZN(c[26]));
   OAI21_X1 i_0_54 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_34));
   NAND2_X1 i_0_55 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_35));
   NAND2_X1 i_0_56 (.A1(n_0_37), .A2(n_0_36), .ZN(c[27]));
   OAI21_X1 i_0_57 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_36));
   NAND2_X1 i_0_58 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_37));
   NAND2_X1 i_0_59 (.A1(n_0_39), .A2(n_0_38), .ZN(c[28]));
   OAI21_X1 i_0_60 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_38));
   NAND2_X1 i_0_61 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_39));
   NAND2_X1 i_0_62 (.A1(n_0_41), .A2(n_0_40), .ZN(c[29]));
   OAI21_X1 i_0_63 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_40));
   NAND2_X1 i_0_64 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_41));
   NAND2_X1 i_0_65 (.A1(n_0_43), .A2(n_0_42), .ZN(c[30]));
   OAI21_X1 i_0_66 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_42));
   NAND2_X1 i_0_67 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_43));
   NAND2_X1 i_0_68 (.A1(n_0_45), .A2(n_0_44), .ZN(c[31]));
   OAI21_X1 i_0_69 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_44));
   NAND2_X1 i_0_70 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_45));
   NAND2_X1 i_0_71 (.A1(n_0_47), .A2(n_0_46), .ZN(c[32]));
   OAI21_X1 i_0_72 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_46));
   NAND2_X1 i_0_73 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_47));
   NAND2_X1 i_0_74 (.A1(n_0_49), .A2(n_0_48), .ZN(c[33]));
   OAI21_X1 i_0_75 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_48));
   NAND2_X1 i_0_76 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_49));
   NAND2_X1 i_0_77 (.A1(n_0_51), .A2(n_0_50), .ZN(c[34]));
   OAI21_X1 i_0_78 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_50));
   NAND2_X1 i_0_79 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_51));
   NAND2_X1 i_0_80 (.A1(n_0_53), .A2(n_0_52), .ZN(c[35]));
   OAI21_X1 i_0_81 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_52));
   NAND2_X1 i_0_82 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_53));
   NAND2_X1 i_0_83 (.A1(n_0_55), .A2(n_0_54), .ZN(c[36]));
   OAI21_X1 i_0_84 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_54));
   NAND2_X1 i_0_85 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_55));
   NAND2_X1 i_0_86 (.A1(n_0_57), .A2(n_0_56), .ZN(c[37]));
   OAI21_X1 i_0_87 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_56));
   NAND2_X1 i_0_88 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_57));
   NAND2_X1 i_0_89 (.A1(n_0_59), .A2(n_0_58), .ZN(c[38]));
   OAI21_X1 i_0_90 (.A(in2[37]), .B1(in3[37]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_91 (.A1(in3[37]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_92 (.A1(n_0_61), .A2(n_0_60), .ZN(c[39]));
   OAI21_X1 i_0_93 (.A(in2[38]), .B1(in3[38]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_94 (.A1(in3[38]), .A2(in1[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(n_0_64), .A2(n_0_62), .ZN(c[40]));
   OAI21_X1 i_0_96 (.A(in3[39]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_62));
   NAND2_X1 i_0_97 (.A1(n_0_64), .A2(n_0_63), .ZN(c[63]));
   OAI21_X1 i_0_98 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_63));
   NAND2_X1 i_0_99 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_64));
   XOR2_X1 i_0_100 (.A(in2[6]), .B(in1[6]), .Z(sum[6]));
   XOR2_X1 i_0_101 (.A(in2[7]), .B(in1[7]), .Z(sum[7]));
   XNOR2_X1 i_0_102 (.A(in2[8]), .B(n_0_65), .ZN(sum[8]));
   XNOR2_X1 i_0_103 (.A(in3[8]), .B(in1[8]), .ZN(n_0_65));
   XNOR2_X1 i_0_104 (.A(in2[9]), .B(n_0_66), .ZN(sum[9]));
   XNOR2_X1 i_0_105 (.A(in3[9]), .B(in1[9]), .ZN(n_0_66));
   XNOR2_X1 i_0_106 (.A(in2[10]), .B(n_0_67), .ZN(sum[10]));
   XNOR2_X1 i_0_107 (.A(in3[10]), .B(in1[10]), .ZN(n_0_67));
   XNOR2_X1 i_0_108 (.A(in2[11]), .B(n_0_68), .ZN(sum[11]));
   XNOR2_X1 i_0_109 (.A(in3[11]), .B(in1[11]), .ZN(n_0_68));
   XNOR2_X1 i_0_110 (.A(in2[12]), .B(n_0_69), .ZN(sum[12]));
   XNOR2_X1 i_0_111 (.A(in3[12]), .B(in1[12]), .ZN(n_0_69));
   XNOR2_X1 i_0_112 (.A(in2[13]), .B(n_0_70), .ZN(sum[13]));
   XNOR2_X1 i_0_113 (.A(in3[13]), .B(in1[13]), .ZN(n_0_70));
   XNOR2_X1 i_0_114 (.A(in2[14]), .B(n_0_71), .ZN(sum[14]));
   XNOR2_X1 i_0_115 (.A(in3[14]), .B(in1[14]), .ZN(n_0_71));
   XNOR2_X1 i_0_116 (.A(in2[15]), .B(n_0_72), .ZN(sum[15]));
   XNOR2_X1 i_0_117 (.A(in3[15]), .B(in1[15]), .ZN(n_0_72));
   XNOR2_X1 i_0_118 (.A(in2[16]), .B(n_0_73), .ZN(sum[16]));
   XNOR2_X1 i_0_119 (.A(in3[16]), .B(in1[16]), .ZN(n_0_73));
   XNOR2_X1 i_0_120 (.A(in2[17]), .B(n_0_74), .ZN(sum[17]));
   XNOR2_X1 i_0_121 (.A(in3[17]), .B(in1[17]), .ZN(n_0_74));
   XNOR2_X1 i_0_122 (.A(in2[18]), .B(n_0_75), .ZN(sum[18]));
   XNOR2_X1 i_0_123 (.A(in3[18]), .B(in1[18]), .ZN(n_0_75));
   XNOR2_X1 i_0_124 (.A(in2[19]), .B(n_0_76), .ZN(sum[19]));
   XNOR2_X1 i_0_125 (.A(in3[19]), .B(in1[19]), .ZN(n_0_76));
   XNOR2_X1 i_0_126 (.A(in2[20]), .B(n_0_77), .ZN(sum[20]));
   XNOR2_X1 i_0_127 (.A(in3[20]), .B(in1[20]), .ZN(n_0_77));
   XNOR2_X1 i_0_128 (.A(in2[21]), .B(n_0_78), .ZN(sum[21]));
   XNOR2_X1 i_0_129 (.A(in3[21]), .B(in1[21]), .ZN(n_0_78));
   XNOR2_X1 i_0_130 (.A(in2[22]), .B(n_0_79), .ZN(sum[22]));
   XNOR2_X1 i_0_131 (.A(in3[22]), .B(in1[22]), .ZN(n_0_79));
   XNOR2_X1 i_0_132 (.A(in2[23]), .B(n_0_80), .ZN(sum[23]));
   XNOR2_X1 i_0_133 (.A(in3[23]), .B(in1[23]), .ZN(n_0_80));
   XNOR2_X1 i_0_134 (.A(in2[24]), .B(n_0_81), .ZN(sum[24]));
   XNOR2_X1 i_0_135 (.A(in3[24]), .B(in1[24]), .ZN(n_0_81));
   XNOR2_X1 i_0_136 (.A(in2[25]), .B(n_0_82), .ZN(sum[25]));
   XNOR2_X1 i_0_137 (.A(in3[25]), .B(in1[25]), .ZN(n_0_82));
   XNOR2_X1 i_0_138 (.A(in2[26]), .B(n_0_83), .ZN(sum[26]));
   XNOR2_X1 i_0_139 (.A(in3[26]), .B(in1[26]), .ZN(n_0_83));
   XNOR2_X1 i_0_140 (.A(in2[27]), .B(n_0_84), .ZN(sum[27]));
   XNOR2_X1 i_0_141 (.A(in3[27]), .B(in1[27]), .ZN(n_0_84));
   XNOR2_X1 i_0_142 (.A(in2[28]), .B(n_0_85), .ZN(sum[28]));
   XNOR2_X1 i_0_143 (.A(in3[28]), .B(in1[28]), .ZN(n_0_85));
   XNOR2_X1 i_0_144 (.A(in2[29]), .B(n_0_86), .ZN(sum[29]));
   XNOR2_X1 i_0_145 (.A(in3[29]), .B(in1[29]), .ZN(n_0_86));
   XNOR2_X1 i_0_146 (.A(in2[30]), .B(n_0_87), .ZN(sum[30]));
   XNOR2_X1 i_0_147 (.A(in3[30]), .B(in1[30]), .ZN(n_0_87));
   XNOR2_X1 i_0_148 (.A(in2[31]), .B(n_0_88), .ZN(sum[31]));
   XNOR2_X1 i_0_149 (.A(in3[31]), .B(in1[31]), .ZN(n_0_88));
   XNOR2_X1 i_0_150 (.A(in2[32]), .B(n_0_89), .ZN(sum[32]));
   XNOR2_X1 i_0_151 (.A(in3[32]), .B(in1[32]), .ZN(n_0_89));
   XNOR2_X1 i_0_152 (.A(in2[33]), .B(n_0_90), .ZN(sum[33]));
   XNOR2_X1 i_0_153 (.A(in3[33]), .B(in1[33]), .ZN(n_0_90));
   XNOR2_X1 i_0_154 (.A(in2[34]), .B(n_0_91), .ZN(sum[34]));
   XNOR2_X1 i_0_155 (.A(in3[34]), .B(in1[34]), .ZN(n_0_91));
   XNOR2_X1 i_0_156 (.A(in2[35]), .B(n_0_92), .ZN(sum[35]));
   XNOR2_X1 i_0_157 (.A(in3[35]), .B(in1[35]), .ZN(n_0_92));
   XNOR2_X1 i_0_158 (.A(in2[36]), .B(n_0_93), .ZN(sum[36]));
   XNOR2_X1 i_0_159 (.A(in3[36]), .B(in1[36]), .ZN(n_0_93));
   XNOR2_X1 i_0_160 (.A(in2[37]), .B(n_0_94), .ZN(sum[37]));
   XNOR2_X1 i_0_161 (.A(in3[37]), .B(in1[63]), .ZN(n_0_94));
   XNOR2_X1 i_0_162 (.A(in2[38]), .B(n_0_95), .ZN(sum[38]));
   XNOR2_X1 i_0_163 (.A(in3[38]), .B(in1[63]), .ZN(n_0_95));
   XOR2_X1 i_0_164 (.A(in3[39]), .B(n_0_96), .Z(sum[39]));
   INV_X1 i_0_165 (.A(n_0_97), .ZN(n_0_96));
   NAND2_X1 i_0_166 (.A1(n_0_102), .A2(n_0_101), .ZN(n_0_97));
   NOR2_X1 i_0_167 (.A1(n_0_98), .A2(n_0_100), .ZN(sum[63]));
   INV_X1 i_0_168 (.A(n_0_99), .ZN(n_0_98));
   NAND3_X1 i_0_169 (.A1(n_0_102), .A2(in3[63]), .A3(n_0_101), .ZN(n_0_99));
   AOI21_X1 i_0_170 (.A(in3[63]), .B1(n_0_102), .B2(n_0_101), .ZN(n_0_100));
   NAND2_X1 i_0_171 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_101));
   NAND2_X1 i_0_172 (.A1(n_0_104), .A2(n_0_103), .ZN(n_0_102));
   INV_X1 i_0_173 (.A(in1[63]), .ZN(n_0_103));
   INV_X1 i_0_174 (.A(in2[63]), .ZN(n_0_104));
endmodule

module CSA__1_17(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;

   AND2_X1 i_0_0 (.A1(in2[3]), .A2(in1[3]), .ZN(c[4]));
   AND2_X1 i_0_1 (.A1(in2[4]), .A2(in1[4]), .ZN(c[5]));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_0), .ZN(c[6]));
   OAI21_X1 i_0_3 (.A(in2[5]), .B1(in3[5]), .B2(in1[5]), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(in3[5]), .A2(in1[5]), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .ZN(c[7]));
   OAI21_X1 i_0_6 (.A(in2[6]), .B1(in3[6]), .B2(in1[6]), .ZN(n_0_2));
   NAND2_X1 i_0_7 (.A1(in3[6]), .A2(in1[6]), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_4), .ZN(c[8]));
   OAI21_X1 i_0_9 (.A(in2[7]), .B1(in3[7]), .B2(in1[7]), .ZN(n_0_4));
   NAND2_X1 i_0_10 (.A1(in3[7]), .A2(in1[7]), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(n_0_7), .A2(n_0_6), .ZN(c[9]));
   OAI21_X1 i_0_12 (.A(in2[8]), .B1(in3[8]), .B2(in1[8]), .ZN(n_0_6));
   NAND2_X1 i_0_13 (.A1(in3[8]), .A2(in1[8]), .ZN(n_0_7));
   NAND2_X1 i_0_14 (.A1(n_0_9), .A2(n_0_8), .ZN(c[10]));
   OAI21_X1 i_0_15 (.A(in2[9]), .B1(in3[9]), .B2(in1[9]), .ZN(n_0_8));
   NAND2_X1 i_0_16 (.A1(in3[9]), .A2(in1[9]), .ZN(n_0_9));
   NAND2_X1 i_0_17 (.A1(n_0_11), .A2(n_0_10), .ZN(c[11]));
   OAI21_X1 i_0_18 (.A(in2[10]), .B1(in3[10]), .B2(in1[10]), .ZN(n_0_10));
   NAND2_X1 i_0_19 (.A1(in3[10]), .A2(in1[10]), .ZN(n_0_11));
   NAND2_X1 i_0_20 (.A1(n_0_13), .A2(n_0_12), .ZN(c[12]));
   OAI21_X1 i_0_21 (.A(in2[11]), .B1(in3[11]), .B2(in1[11]), .ZN(n_0_12));
   NAND2_X1 i_0_22 (.A1(in3[11]), .A2(in1[11]), .ZN(n_0_13));
   NAND2_X1 i_0_23 (.A1(n_0_15), .A2(n_0_14), .ZN(c[13]));
   OAI21_X1 i_0_24 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_14));
   NAND2_X1 i_0_25 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_15));
   NAND2_X1 i_0_26 (.A1(n_0_17), .A2(n_0_16), .ZN(c[14]));
   OAI21_X1 i_0_27 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_16));
   NAND2_X1 i_0_28 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_17));
   NAND2_X1 i_0_29 (.A1(n_0_19), .A2(n_0_18), .ZN(c[15]));
   OAI21_X1 i_0_30 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_18));
   NAND2_X1 i_0_31 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_19));
   NAND2_X1 i_0_32 (.A1(n_0_21), .A2(n_0_20), .ZN(c[16]));
   OAI21_X1 i_0_33 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_20));
   NAND2_X1 i_0_34 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_21));
   NAND2_X1 i_0_35 (.A1(n_0_23), .A2(n_0_22), .ZN(c[17]));
   OAI21_X1 i_0_36 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_22));
   NAND2_X1 i_0_37 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_23));
   NAND2_X1 i_0_38 (.A1(n_0_25), .A2(n_0_24), .ZN(c[18]));
   OAI21_X1 i_0_39 (.A(in1[17]), .B1(in3[17]), .B2(in2[17]), .ZN(n_0_24));
   NAND2_X1 i_0_40 (.A1(in2[17]), .A2(in3[17]), .ZN(n_0_25));
   NAND2_X1 i_0_41 (.A1(n_0_27), .A2(n_0_26), .ZN(c[19]));
   OAI21_X1 i_0_42 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_26));
   NAND2_X1 i_0_43 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_27));
   NAND2_X1 i_0_44 (.A1(n_0_29), .A2(n_0_28), .ZN(c[20]));
   OAI21_X1 i_0_45 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_28));
   NAND2_X1 i_0_46 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_29));
   NAND2_X1 i_0_47 (.A1(n_0_31), .A2(n_0_30), .ZN(c[21]));
   OAI21_X1 i_0_48 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_30));
   NAND2_X1 i_0_49 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_31));
   NAND2_X1 i_0_50 (.A1(n_0_33), .A2(n_0_32), .ZN(c[22]));
   OAI21_X1 i_0_51 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_32));
   NAND2_X1 i_0_52 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_33));
   NAND2_X1 i_0_53 (.A1(n_0_35), .A2(n_0_34), .ZN(c[23]));
   OAI21_X1 i_0_54 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_34));
   NAND2_X1 i_0_55 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_35));
   NAND2_X1 i_0_56 (.A1(n_0_37), .A2(n_0_36), .ZN(c[24]));
   OAI21_X1 i_0_57 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_36));
   NAND2_X1 i_0_58 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_37));
   NAND2_X1 i_0_59 (.A1(n_0_39), .A2(n_0_38), .ZN(c[25]));
   OAI21_X1 i_0_60 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_38));
   NAND2_X1 i_0_61 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_39));
   NAND2_X1 i_0_62 (.A1(n_0_41), .A2(n_0_40), .ZN(c[26]));
   OAI21_X1 i_0_63 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_40));
   NAND2_X1 i_0_64 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_41));
   NAND2_X1 i_0_65 (.A1(n_0_43), .A2(n_0_42), .ZN(c[27]));
   OAI21_X1 i_0_66 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_42));
   NAND2_X1 i_0_67 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_43));
   NAND2_X1 i_0_68 (.A1(n_0_45), .A2(n_0_44), .ZN(c[28]));
   OAI21_X1 i_0_69 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_44));
   NAND2_X1 i_0_70 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_45));
   NAND2_X1 i_0_71 (.A1(n_0_47), .A2(n_0_46), .ZN(c[29]));
   OAI21_X1 i_0_72 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_46));
   NAND2_X1 i_0_73 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_47));
   NAND2_X1 i_0_74 (.A1(n_0_49), .A2(n_0_48), .ZN(c[30]));
   OAI21_X1 i_0_75 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_48));
   NAND2_X1 i_0_76 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_49));
   NAND2_X1 i_0_77 (.A1(n_0_51), .A2(n_0_50), .ZN(c[31]));
   OAI21_X1 i_0_78 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_50));
   NAND2_X1 i_0_79 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_51));
   NAND2_X1 i_0_80 (.A1(n_0_53), .A2(n_0_52), .ZN(c[32]));
   OAI21_X1 i_0_81 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_52));
   NAND2_X1 i_0_82 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_53));
   NAND2_X1 i_0_83 (.A1(n_0_55), .A2(n_0_54), .ZN(c[33]));
   OAI21_X1 i_0_84 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_54));
   NAND2_X1 i_0_85 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_55));
   NAND2_X1 i_0_86 (.A1(n_0_57), .A2(n_0_56), .ZN(c[34]));
   OAI21_X1 i_0_87 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_56));
   NAND2_X1 i_0_88 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_57));
   NAND2_X1 i_0_89 (.A1(n_0_59), .A2(n_0_58), .ZN(c[35]));
   OAI21_X1 i_0_90 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_58));
   NAND2_X1 i_0_91 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_59));
   NAND2_X1 i_0_92 (.A1(n_0_61), .A2(n_0_60), .ZN(c[36]));
   OAI21_X1 i_0_93 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_60));
   NAND2_X1 i_0_94 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(n_0_63), .A2(n_0_62), .ZN(c[37]));
   OAI21_X1 i_0_96 (.A(in2[36]), .B1(in3[36]), .B2(in1[63]), .ZN(n_0_62));
   NAND2_X1 i_0_97 (.A1(in3[36]), .A2(in1[63]), .ZN(n_0_63));
   AOI21_X1 i_0_98 (.A(n_0_65), .B1(n_0_64), .B2(n_0_99), .ZN(c[38]));
   AOI21_X1 i_0_99 (.A(n_0_65), .B1(n_0_64), .B2(n_0_100), .ZN(c[39]));
   AOI21_X1 i_0_100 (.A(n_0_65), .B1(n_0_64), .B2(n_0_101), .ZN(c[40]));
   AOI21_X1 i_0_101 (.A(n_0_65), .B1(n_0_64), .B2(n_0_102), .ZN(c[63]));
   NAND2_X1 i_0_102 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_64));
   NOR2_X1 i_0_103 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_65));
   XOR2_X1 i_0_104 (.A(in2[3]), .B(in1[3]), .Z(sum[3]));
   XOR2_X1 i_0_105 (.A(in2[4]), .B(in1[4]), .Z(sum[4]));
   XNOR2_X1 i_0_106 (.A(in2[5]), .B(n_0_66), .ZN(sum[5]));
   XNOR2_X1 i_0_107 (.A(in3[5]), .B(in1[5]), .ZN(n_0_66));
   XNOR2_X1 i_0_108 (.A(in2[6]), .B(n_0_67), .ZN(sum[6]));
   XNOR2_X1 i_0_109 (.A(in3[6]), .B(in1[6]), .ZN(n_0_67));
   XNOR2_X1 i_0_110 (.A(in2[7]), .B(n_0_68), .ZN(sum[7]));
   XNOR2_X1 i_0_111 (.A(in3[7]), .B(in1[7]), .ZN(n_0_68));
   XNOR2_X1 i_0_112 (.A(in2[8]), .B(n_0_69), .ZN(sum[8]));
   XNOR2_X1 i_0_113 (.A(in3[8]), .B(in1[8]), .ZN(n_0_69));
   XNOR2_X1 i_0_114 (.A(in2[9]), .B(n_0_70), .ZN(sum[9]));
   XNOR2_X1 i_0_115 (.A(in3[9]), .B(in1[9]), .ZN(n_0_70));
   XNOR2_X1 i_0_116 (.A(in2[10]), .B(n_0_71), .ZN(sum[10]));
   XNOR2_X1 i_0_117 (.A(in3[10]), .B(in1[10]), .ZN(n_0_71));
   XNOR2_X1 i_0_118 (.A(in2[11]), .B(n_0_72), .ZN(sum[11]));
   XNOR2_X1 i_0_119 (.A(in3[11]), .B(in1[11]), .ZN(n_0_72));
   XNOR2_X1 i_0_120 (.A(in2[12]), .B(n_0_73), .ZN(sum[12]));
   XNOR2_X1 i_0_121 (.A(in3[12]), .B(in1[12]), .ZN(n_0_73));
   XNOR2_X1 i_0_122 (.A(in2[13]), .B(n_0_74), .ZN(sum[13]));
   XNOR2_X1 i_0_123 (.A(in3[13]), .B(in1[13]), .ZN(n_0_74));
   XNOR2_X1 i_0_124 (.A(in2[14]), .B(n_0_75), .ZN(sum[14]));
   XNOR2_X1 i_0_125 (.A(in3[14]), .B(in1[14]), .ZN(n_0_75));
   XNOR2_X1 i_0_126 (.A(in2[15]), .B(n_0_76), .ZN(sum[15]));
   XNOR2_X1 i_0_127 (.A(in3[15]), .B(in1[15]), .ZN(n_0_76));
   XNOR2_X1 i_0_128 (.A(in2[16]), .B(n_0_77), .ZN(sum[16]));
   XNOR2_X1 i_0_129 (.A(in3[16]), .B(in1[16]), .ZN(n_0_77));
   XNOR2_X1 i_0_130 (.A(in2[17]), .B(n_0_78), .ZN(sum[17]));
   XNOR2_X1 i_0_131 (.A(in3[17]), .B(in1[17]), .ZN(n_0_78));
   XNOR2_X1 i_0_132 (.A(in2[18]), .B(n_0_79), .ZN(sum[18]));
   XNOR2_X1 i_0_133 (.A(in3[18]), .B(in1[18]), .ZN(n_0_79));
   XNOR2_X1 i_0_134 (.A(in2[19]), .B(n_0_80), .ZN(sum[19]));
   XNOR2_X1 i_0_135 (.A(in3[19]), .B(in1[19]), .ZN(n_0_80));
   XNOR2_X1 i_0_136 (.A(in2[20]), .B(n_0_81), .ZN(sum[20]));
   XNOR2_X1 i_0_137 (.A(in3[20]), .B(in1[20]), .ZN(n_0_81));
   XNOR2_X1 i_0_138 (.A(in2[21]), .B(n_0_82), .ZN(sum[21]));
   XNOR2_X1 i_0_139 (.A(in3[21]), .B(in1[21]), .ZN(n_0_82));
   XNOR2_X1 i_0_140 (.A(in2[22]), .B(n_0_83), .ZN(sum[22]));
   XNOR2_X1 i_0_141 (.A(in3[22]), .B(in1[22]), .ZN(n_0_83));
   XNOR2_X1 i_0_142 (.A(in2[23]), .B(n_0_84), .ZN(sum[23]));
   XNOR2_X1 i_0_143 (.A(in3[23]), .B(in1[23]), .ZN(n_0_84));
   XNOR2_X1 i_0_144 (.A(in2[24]), .B(n_0_85), .ZN(sum[24]));
   XNOR2_X1 i_0_145 (.A(in3[24]), .B(in1[24]), .ZN(n_0_85));
   XNOR2_X1 i_0_146 (.A(in2[25]), .B(n_0_86), .ZN(sum[25]));
   XNOR2_X1 i_0_147 (.A(in3[25]), .B(in1[25]), .ZN(n_0_86));
   XNOR2_X1 i_0_148 (.A(in2[26]), .B(n_0_87), .ZN(sum[26]));
   XNOR2_X1 i_0_149 (.A(in3[26]), .B(in1[26]), .ZN(n_0_87));
   XNOR2_X1 i_0_150 (.A(in2[27]), .B(n_0_88), .ZN(sum[27]));
   XNOR2_X1 i_0_151 (.A(in3[27]), .B(in1[27]), .ZN(n_0_88));
   XNOR2_X1 i_0_152 (.A(in2[28]), .B(n_0_89), .ZN(sum[28]));
   XNOR2_X1 i_0_153 (.A(in3[28]), .B(in1[28]), .ZN(n_0_89));
   XNOR2_X1 i_0_154 (.A(in2[29]), .B(n_0_90), .ZN(sum[29]));
   XNOR2_X1 i_0_155 (.A(in3[29]), .B(in1[29]), .ZN(n_0_90));
   XNOR2_X1 i_0_156 (.A(in2[30]), .B(n_0_91), .ZN(sum[30]));
   XNOR2_X1 i_0_157 (.A(in3[30]), .B(in1[30]), .ZN(n_0_91));
   XNOR2_X1 i_0_158 (.A(in2[31]), .B(n_0_92), .ZN(sum[31]));
   XNOR2_X1 i_0_159 (.A(in3[31]), .B(in1[31]), .ZN(n_0_92));
   XNOR2_X1 i_0_160 (.A(in2[32]), .B(n_0_93), .ZN(sum[32]));
   XNOR2_X1 i_0_161 (.A(in3[32]), .B(in1[32]), .ZN(n_0_93));
   XNOR2_X1 i_0_162 (.A(in2[33]), .B(n_0_94), .ZN(sum[33]));
   XNOR2_X1 i_0_163 (.A(in3[33]), .B(in1[33]), .ZN(n_0_94));
   XNOR2_X1 i_0_164 (.A(in2[34]), .B(n_0_95), .ZN(sum[34]));
   XNOR2_X1 i_0_165 (.A(in3[34]), .B(in1[34]), .ZN(n_0_95));
   XNOR2_X1 i_0_166 (.A(in2[35]), .B(n_0_96), .ZN(sum[35]));
   XNOR2_X1 i_0_167 (.A(in3[35]), .B(in1[35]), .ZN(n_0_96));
   XNOR2_X1 i_0_168 (.A(in2[36]), .B(n_0_97), .ZN(sum[36]));
   XNOR2_X1 i_0_169 (.A(in3[36]), .B(in1[63]), .ZN(n_0_97));
   XNOR2_X1 i_0_170 (.A(n_0_99), .B(n_0_98), .ZN(sum[37]));
   XNOR2_X1 i_0_171 (.A(n_0_100), .B(n_0_98), .ZN(sum[38]));
   XNOR2_X1 i_0_172 (.A(n_0_101), .B(n_0_98), .ZN(sum[39]));
   XNOR2_X1 i_0_173 (.A(n_0_102), .B(n_0_98), .ZN(sum[63]));
   XOR2_X1 i_0_174 (.A(in2[63]), .B(in1[63]), .Z(n_0_98));
   INV_X1 i_0_175 (.A(in3[37]), .ZN(n_0_99));
   INV_X1 i_0_176 (.A(in3[38]), .ZN(n_0_100));
   INV_X1 i_0_177 (.A(in3[39]), .ZN(n_0_101));
   INV_X1 i_0_178 (.A(in3[63]), .ZN(n_0_102));
endmodule

module CSA__1_20(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;

   AND2_X1 i_0_0 (.A1(in2[10]), .A2(in1[10]), .ZN(c[11]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[12]));
   OAI21_X1 i_0_2 (.A(in2[11]), .B1(in3[11]), .B2(in1[11]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[11]), .A2(in1[11]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[13]));
   OAI21_X1 i_0_5 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[14]));
   OAI21_X1 i_0_8 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[15]));
   OAI21_X1 i_0_11 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[16]));
   OAI21_X1 i_0_14 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[17]));
   OAI21_X1 i_0_17 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[18]));
   OAI21_X1 i_0_20 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[19]));
   OAI21_X1 i_0_23 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[20]));
   OAI21_X1 i_0_26 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[21]));
   OAI21_X1 i_0_29 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[22]));
   OAI21_X1 i_0_32 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[23]));
   OAI21_X1 i_0_35 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[24]));
   OAI21_X1 i_0_38 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[25]));
   OAI21_X1 i_0_41 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[26]));
   OAI21_X1 i_0_44 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[27]));
   OAI21_X1 i_0_47 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[28]));
   OAI21_X1 i_0_50 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[29]));
   OAI21_X1 i_0_53 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[30]));
   OAI21_X1 i_0_56 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[31]));
   OAI21_X1 i_0_59 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[32]));
   OAI21_X1 i_0_62 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[33]));
   OAI21_X1 i_0_65 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[34]));
   OAI21_X1 i_0_68 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[35]));
   OAI21_X1 i_0_71 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[36]));
   OAI21_X1 i_0_74 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[37]));
   OAI21_X1 i_0_77 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[38]));
   OAI21_X1 i_0_80 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[39]));
   OAI21_X1 i_0_83 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[40]));
   OAI21_X1 i_0_86 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[41]));
   OAI21_X1 i_0_89 (.A(in2[40]), .B1(in3[40]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[40]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_62), .A2(n_0_60), .ZN(c[42]));
   OAI21_X1 i_0_92 (.A(in3[41]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(c[63]));
   OAI21_X1 i_0_94 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   XOR2_X1 i_0_96 (.A(in2[10]), .B(in1[10]), .Z(sum[10]));
   XNOR2_X1 i_0_97 (.A(in2[11]), .B(n_0_63), .ZN(sum[11]));
   XNOR2_X1 i_0_98 (.A(in3[11]), .B(in1[11]), .ZN(n_0_63));
   XNOR2_X1 i_0_99 (.A(in2[12]), .B(n_0_64), .ZN(sum[12]));
   XNOR2_X1 i_0_100 (.A(in3[12]), .B(in1[12]), .ZN(n_0_64));
   XNOR2_X1 i_0_101 (.A(in2[13]), .B(n_0_65), .ZN(sum[13]));
   XNOR2_X1 i_0_102 (.A(in3[13]), .B(in1[13]), .ZN(n_0_65));
   XNOR2_X1 i_0_103 (.A(in2[14]), .B(n_0_66), .ZN(sum[14]));
   XNOR2_X1 i_0_104 (.A(in3[14]), .B(in1[14]), .ZN(n_0_66));
   XNOR2_X1 i_0_105 (.A(in2[15]), .B(n_0_67), .ZN(sum[15]));
   XNOR2_X1 i_0_106 (.A(in3[15]), .B(in1[15]), .ZN(n_0_67));
   XNOR2_X1 i_0_107 (.A(in2[16]), .B(n_0_68), .ZN(sum[16]));
   XNOR2_X1 i_0_108 (.A(in3[16]), .B(in1[16]), .ZN(n_0_68));
   XNOR2_X1 i_0_109 (.A(in2[17]), .B(n_0_69), .ZN(sum[17]));
   XNOR2_X1 i_0_110 (.A(in3[17]), .B(in1[17]), .ZN(n_0_69));
   XNOR2_X1 i_0_111 (.A(in2[18]), .B(n_0_70), .ZN(sum[18]));
   XNOR2_X1 i_0_112 (.A(in3[18]), .B(in1[18]), .ZN(n_0_70));
   XNOR2_X1 i_0_113 (.A(in2[19]), .B(n_0_71), .ZN(sum[19]));
   XNOR2_X1 i_0_114 (.A(in3[19]), .B(in1[19]), .ZN(n_0_71));
   XNOR2_X1 i_0_115 (.A(in2[20]), .B(n_0_72), .ZN(sum[20]));
   XNOR2_X1 i_0_116 (.A(in3[20]), .B(in1[20]), .ZN(n_0_72));
   XNOR2_X1 i_0_117 (.A(in2[21]), .B(n_0_73), .ZN(sum[21]));
   XNOR2_X1 i_0_118 (.A(in3[21]), .B(in1[21]), .ZN(n_0_73));
   XNOR2_X1 i_0_119 (.A(in2[22]), .B(n_0_74), .ZN(sum[22]));
   XNOR2_X1 i_0_120 (.A(in3[22]), .B(in1[22]), .ZN(n_0_74));
   XNOR2_X1 i_0_121 (.A(in2[23]), .B(n_0_75), .ZN(sum[23]));
   XNOR2_X1 i_0_122 (.A(in3[23]), .B(in1[23]), .ZN(n_0_75));
   XNOR2_X1 i_0_123 (.A(in2[24]), .B(n_0_76), .ZN(sum[24]));
   XNOR2_X1 i_0_124 (.A(in3[24]), .B(in1[24]), .ZN(n_0_76));
   XNOR2_X1 i_0_125 (.A(in2[25]), .B(n_0_77), .ZN(sum[25]));
   XNOR2_X1 i_0_126 (.A(in3[25]), .B(in1[25]), .ZN(n_0_77));
   XNOR2_X1 i_0_127 (.A(in2[26]), .B(n_0_78), .ZN(sum[26]));
   XNOR2_X1 i_0_128 (.A(in3[26]), .B(in1[26]), .ZN(n_0_78));
   XNOR2_X1 i_0_129 (.A(in2[27]), .B(n_0_79), .ZN(sum[27]));
   XNOR2_X1 i_0_130 (.A(in3[27]), .B(in1[27]), .ZN(n_0_79));
   XNOR2_X1 i_0_131 (.A(in2[28]), .B(n_0_80), .ZN(sum[28]));
   XNOR2_X1 i_0_132 (.A(in3[28]), .B(in1[28]), .ZN(n_0_80));
   XNOR2_X1 i_0_133 (.A(in2[29]), .B(n_0_81), .ZN(sum[29]));
   XNOR2_X1 i_0_134 (.A(in3[29]), .B(in1[29]), .ZN(n_0_81));
   XNOR2_X1 i_0_135 (.A(in2[30]), .B(n_0_82), .ZN(sum[30]));
   XNOR2_X1 i_0_136 (.A(in3[30]), .B(in1[30]), .ZN(n_0_82));
   XNOR2_X1 i_0_137 (.A(in2[31]), .B(n_0_83), .ZN(sum[31]));
   XNOR2_X1 i_0_138 (.A(in3[31]), .B(in1[31]), .ZN(n_0_83));
   XNOR2_X1 i_0_139 (.A(in2[32]), .B(n_0_84), .ZN(sum[32]));
   XNOR2_X1 i_0_140 (.A(in3[32]), .B(in1[32]), .ZN(n_0_84));
   XNOR2_X1 i_0_141 (.A(in2[33]), .B(n_0_85), .ZN(sum[33]));
   XNOR2_X1 i_0_142 (.A(in3[33]), .B(in1[33]), .ZN(n_0_85));
   XNOR2_X1 i_0_143 (.A(in2[34]), .B(n_0_86), .ZN(sum[34]));
   XNOR2_X1 i_0_144 (.A(in3[34]), .B(in1[34]), .ZN(n_0_86));
   XNOR2_X1 i_0_145 (.A(in2[35]), .B(n_0_87), .ZN(sum[35]));
   XNOR2_X1 i_0_146 (.A(in3[35]), .B(in1[35]), .ZN(n_0_87));
   XNOR2_X1 i_0_147 (.A(in2[36]), .B(n_0_88), .ZN(sum[36]));
   XNOR2_X1 i_0_148 (.A(in3[36]), .B(in1[36]), .ZN(n_0_88));
   XNOR2_X1 i_0_149 (.A(in2[37]), .B(n_0_89), .ZN(sum[37]));
   XNOR2_X1 i_0_150 (.A(in3[37]), .B(in1[37]), .ZN(n_0_89));
   XNOR2_X1 i_0_151 (.A(in2[38]), .B(n_0_90), .ZN(sum[38]));
   XNOR2_X1 i_0_152 (.A(in3[38]), .B(in1[38]), .ZN(n_0_90));
   XNOR2_X1 i_0_153 (.A(in2[39]), .B(n_0_91), .ZN(sum[39]));
   XNOR2_X1 i_0_154 (.A(in3[39]), .B(in1[39]), .ZN(n_0_91));
   XNOR2_X1 i_0_155 (.A(in2[40]), .B(n_0_92), .ZN(sum[40]));
   XNOR2_X1 i_0_156 (.A(in3[40]), .B(in1[63]), .ZN(n_0_92));
   XOR2_X1 i_0_157 (.A(in3[41]), .B(n_0_93), .Z(sum[41]));
   XOR2_X1 i_0_158 (.A(in3[63]), .B(n_0_93), .Z(sum[63]));
   XOR2_X1 i_0_159 (.A(in2[63]), .B(in1[63]), .Z(n_0_93));
endmodule

module CSA__1_23(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;

   AND2_X1 i_0_0 (.A1(in2[25]), .A2(in1[25]), .ZN(c[26]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[27]));
   OAI21_X1 i_0_2 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[28]));
   OAI21_X1 i_0_5 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[29]));
   OAI21_X1 i_0_8 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[30]));
   OAI21_X1 i_0_11 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[31]));
   OAI21_X1 i_0_14 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[32]));
   OAI21_X1 i_0_17 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[33]));
   OAI21_X1 i_0_20 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[34]));
   OAI21_X1 i_0_23 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[35]));
   OAI21_X1 i_0_26 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[36]));
   OAI21_X1 i_0_29 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[37]));
   OAI21_X1 i_0_32 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[38]));
   OAI21_X1 i_0_35 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[39]));
   OAI21_X1 i_0_38 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[40]));
   OAI21_X1 i_0_41 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[41]));
   OAI21_X1 i_0_44 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[42]));
   OAI21_X1 i_0_47 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[43]));
   OAI21_X1 i_0_50 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[44]));
   OAI21_X1 i_0_53 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[45]));
   OAI21_X1 i_0_56 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[46]));
   OAI21_X1 i_0_59 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[47]));
   OAI21_X1 i_0_62 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[48]));
   OAI21_X1 i_0_65 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[49]));
   OAI21_X1 i_0_68 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[50]));
   OAI21_X1 i_0_71 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[51]));
   OAI21_X1 i_0_74 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[52]));
   OAI21_X1 i_0_77 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[53]));
   OAI21_X1 i_0_80 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[54]));
   OAI21_X1 i_0_83 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[55]));
   OAI21_X1 i_0_86 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[56]));
   OAI21_X1 i_0_89 (.A(in2[55]), .B1(in3[55]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[55]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_62), .A2(n_0_60), .ZN(c[57]));
   OAI21_X1 i_0_92 (.A(in3[56]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(c[63]));
   OAI21_X1 i_0_94 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   XOR2_X1 i_0_96 (.A(in2[25]), .B(in1[25]), .Z(sum[25]));
   XNOR2_X1 i_0_97 (.A(in2[26]), .B(n_0_63), .ZN(sum[26]));
   XNOR2_X1 i_0_98 (.A(in3[26]), .B(in1[26]), .ZN(n_0_63));
   XNOR2_X1 i_0_99 (.A(in2[27]), .B(n_0_64), .ZN(sum[27]));
   XNOR2_X1 i_0_100 (.A(in3[27]), .B(in1[27]), .ZN(n_0_64));
   XNOR2_X1 i_0_101 (.A(in2[28]), .B(n_0_65), .ZN(sum[28]));
   XNOR2_X1 i_0_102 (.A(in3[28]), .B(in1[28]), .ZN(n_0_65));
   XNOR2_X1 i_0_103 (.A(in2[29]), .B(n_0_66), .ZN(sum[29]));
   XNOR2_X1 i_0_104 (.A(in3[29]), .B(in1[29]), .ZN(n_0_66));
   XNOR2_X1 i_0_105 (.A(in2[30]), .B(n_0_67), .ZN(sum[30]));
   XNOR2_X1 i_0_106 (.A(in3[30]), .B(in1[30]), .ZN(n_0_67));
   XNOR2_X1 i_0_107 (.A(in2[31]), .B(n_0_68), .ZN(sum[31]));
   XNOR2_X1 i_0_108 (.A(in3[31]), .B(in1[31]), .ZN(n_0_68));
   XNOR2_X1 i_0_109 (.A(in2[32]), .B(n_0_69), .ZN(sum[32]));
   XNOR2_X1 i_0_110 (.A(in3[32]), .B(in1[32]), .ZN(n_0_69));
   XNOR2_X1 i_0_111 (.A(in2[33]), .B(n_0_70), .ZN(sum[33]));
   XNOR2_X1 i_0_112 (.A(in3[33]), .B(in1[33]), .ZN(n_0_70));
   XNOR2_X1 i_0_113 (.A(in2[34]), .B(n_0_71), .ZN(sum[34]));
   XNOR2_X1 i_0_114 (.A(in3[34]), .B(in1[34]), .ZN(n_0_71));
   XNOR2_X1 i_0_115 (.A(in2[35]), .B(n_0_72), .ZN(sum[35]));
   XNOR2_X1 i_0_116 (.A(in3[35]), .B(in1[35]), .ZN(n_0_72));
   XNOR2_X1 i_0_117 (.A(in2[36]), .B(n_0_73), .ZN(sum[36]));
   XNOR2_X1 i_0_118 (.A(in3[36]), .B(in1[36]), .ZN(n_0_73));
   XNOR2_X1 i_0_119 (.A(in2[37]), .B(n_0_74), .ZN(sum[37]));
   XNOR2_X1 i_0_120 (.A(in3[37]), .B(in1[37]), .ZN(n_0_74));
   XNOR2_X1 i_0_121 (.A(in2[38]), .B(n_0_75), .ZN(sum[38]));
   XNOR2_X1 i_0_122 (.A(in3[38]), .B(in1[38]), .ZN(n_0_75));
   XNOR2_X1 i_0_123 (.A(in2[39]), .B(n_0_76), .ZN(sum[39]));
   XNOR2_X1 i_0_124 (.A(in3[39]), .B(in1[39]), .ZN(n_0_76));
   XNOR2_X1 i_0_125 (.A(in2[40]), .B(n_0_77), .ZN(sum[40]));
   XNOR2_X1 i_0_126 (.A(in3[40]), .B(in1[40]), .ZN(n_0_77));
   XNOR2_X1 i_0_127 (.A(in2[41]), .B(n_0_78), .ZN(sum[41]));
   XNOR2_X1 i_0_128 (.A(in3[41]), .B(in1[41]), .ZN(n_0_78));
   XNOR2_X1 i_0_129 (.A(in2[42]), .B(n_0_79), .ZN(sum[42]));
   XNOR2_X1 i_0_130 (.A(in3[42]), .B(in1[42]), .ZN(n_0_79));
   XNOR2_X1 i_0_131 (.A(in2[43]), .B(n_0_80), .ZN(sum[43]));
   XNOR2_X1 i_0_132 (.A(in3[43]), .B(in1[43]), .ZN(n_0_80));
   XNOR2_X1 i_0_133 (.A(in2[44]), .B(n_0_81), .ZN(sum[44]));
   XNOR2_X1 i_0_134 (.A(in3[44]), .B(in1[44]), .ZN(n_0_81));
   XNOR2_X1 i_0_135 (.A(in2[45]), .B(n_0_82), .ZN(sum[45]));
   XNOR2_X1 i_0_136 (.A(in3[45]), .B(in1[45]), .ZN(n_0_82));
   XNOR2_X1 i_0_137 (.A(in2[46]), .B(n_0_83), .ZN(sum[46]));
   XNOR2_X1 i_0_138 (.A(in3[46]), .B(in1[46]), .ZN(n_0_83));
   XNOR2_X1 i_0_139 (.A(in2[47]), .B(n_0_84), .ZN(sum[47]));
   XNOR2_X1 i_0_140 (.A(in3[47]), .B(in1[47]), .ZN(n_0_84));
   XNOR2_X1 i_0_141 (.A(in2[48]), .B(n_0_85), .ZN(sum[48]));
   XNOR2_X1 i_0_142 (.A(in3[48]), .B(in1[48]), .ZN(n_0_85));
   XNOR2_X1 i_0_143 (.A(in2[49]), .B(n_0_86), .ZN(sum[49]));
   XNOR2_X1 i_0_144 (.A(in3[49]), .B(in1[49]), .ZN(n_0_86));
   XNOR2_X1 i_0_145 (.A(in2[50]), .B(n_0_87), .ZN(sum[50]));
   XNOR2_X1 i_0_146 (.A(in3[50]), .B(in1[50]), .ZN(n_0_87));
   XNOR2_X1 i_0_147 (.A(in2[51]), .B(n_0_88), .ZN(sum[51]));
   XNOR2_X1 i_0_148 (.A(in3[51]), .B(in1[51]), .ZN(n_0_88));
   XNOR2_X1 i_0_149 (.A(in2[52]), .B(n_0_89), .ZN(sum[52]));
   XNOR2_X1 i_0_150 (.A(in3[52]), .B(in1[52]), .ZN(n_0_89));
   XNOR2_X1 i_0_151 (.A(in2[53]), .B(n_0_90), .ZN(sum[53]));
   XNOR2_X1 i_0_152 (.A(in3[53]), .B(in1[53]), .ZN(n_0_90));
   XNOR2_X1 i_0_153 (.A(in2[54]), .B(n_0_91), .ZN(sum[54]));
   XNOR2_X1 i_0_154 (.A(in3[54]), .B(in1[54]), .ZN(n_0_91));
   XNOR2_X1 i_0_155 (.A(in2[55]), .B(n_0_92), .ZN(sum[55]));
   XNOR2_X1 i_0_156 (.A(in3[55]), .B(in1[63]), .ZN(n_0_92));
   XOR2_X1 i_0_157 (.A(in3[56]), .B(n_0_93), .Z(sum[56]));
   XOR2_X1 i_0_158 (.A(in3[63]), .B(n_0_93), .Z(sum[63]));
   XOR2_X1 i_0_159 (.A(in2[63]), .B(in1[63]), .Z(n_0_93));
endmodule

module CSA__1_26(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;

   AND2_X1 i_0_0 (.A1(in2[11]), .A2(in1[11]), .ZN(c[12]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[13]));
   OAI21_X1 i_0_2 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[14]));
   OAI21_X1 i_0_5 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[15]));
   OAI21_X1 i_0_8 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[16]));
   OAI21_X1 i_0_11 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[17]));
   OAI21_X1 i_0_14 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[18]));
   OAI21_X1 i_0_17 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[19]));
   OAI21_X1 i_0_20 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[20]));
   OAI21_X1 i_0_23 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[21]));
   OAI21_X1 i_0_26 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[22]));
   OAI21_X1 i_0_29 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[23]));
   OAI21_X1 i_0_32 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[24]));
   OAI21_X1 i_0_35 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[25]));
   OAI21_X1 i_0_38 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[26]));
   OAI21_X1 i_0_41 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[27]));
   OAI21_X1 i_0_44 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[28]));
   OAI21_X1 i_0_47 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[29]));
   OAI21_X1 i_0_50 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[30]));
   OAI21_X1 i_0_53 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[31]));
   OAI21_X1 i_0_56 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[32]));
   OAI21_X1 i_0_59 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[33]));
   OAI21_X1 i_0_62 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[34]));
   OAI21_X1 i_0_65 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[35]));
   OAI21_X1 i_0_68 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[36]));
   OAI21_X1 i_0_71 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[37]));
   OAI21_X1 i_0_74 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[38]));
   OAI21_X1 i_0_77 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[39]));
   OAI21_X1 i_0_80 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[40]));
   OAI21_X1 i_0_83 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[41]));
   OAI21_X1 i_0_86 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[42]));
   OAI21_X1 i_0_89 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_61), .A2(n_0_60), .ZN(c[43]));
   OAI21_X1 i_0_92 (.A(in2[42]), .B1(in3[42]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(in3[42]), .A2(in1[63]), .ZN(n_0_61));
   AOI21_X1 i_0_94 (.A(n_0_63), .B1(n_0_62), .B2(n_0_96), .ZN(c[44]));
   AOI21_X1 i_0_95 (.A(n_0_63), .B1(n_0_62), .B2(n_0_97), .ZN(c[45]));
   AOI21_X1 i_0_96 (.A(n_0_63), .B1(n_0_62), .B2(n_0_98), .ZN(c[63]));
   NAND2_X1 i_0_97 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   NOR2_X1 i_0_98 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_63));
   XOR2_X1 i_0_99 (.A(in2[11]), .B(in1[11]), .Z(sum[11]));
   XNOR2_X1 i_0_100 (.A(in2[12]), .B(n_0_64), .ZN(sum[12]));
   XNOR2_X1 i_0_101 (.A(in3[12]), .B(in1[12]), .ZN(n_0_64));
   XNOR2_X1 i_0_102 (.A(in2[13]), .B(n_0_65), .ZN(sum[13]));
   XNOR2_X1 i_0_103 (.A(in3[13]), .B(in1[13]), .ZN(n_0_65));
   XNOR2_X1 i_0_104 (.A(in2[14]), .B(n_0_66), .ZN(sum[14]));
   XNOR2_X1 i_0_105 (.A(in3[14]), .B(in1[14]), .ZN(n_0_66));
   XNOR2_X1 i_0_106 (.A(in2[15]), .B(n_0_67), .ZN(sum[15]));
   XNOR2_X1 i_0_107 (.A(in3[15]), .B(in1[15]), .ZN(n_0_67));
   XNOR2_X1 i_0_108 (.A(in2[16]), .B(n_0_68), .ZN(sum[16]));
   XNOR2_X1 i_0_109 (.A(in3[16]), .B(in1[16]), .ZN(n_0_68));
   XNOR2_X1 i_0_110 (.A(in2[17]), .B(n_0_69), .ZN(sum[17]));
   XNOR2_X1 i_0_111 (.A(in3[17]), .B(in1[17]), .ZN(n_0_69));
   XNOR2_X1 i_0_112 (.A(in2[18]), .B(n_0_70), .ZN(sum[18]));
   XNOR2_X1 i_0_113 (.A(in3[18]), .B(in1[18]), .ZN(n_0_70));
   XNOR2_X1 i_0_114 (.A(in2[19]), .B(n_0_71), .ZN(sum[19]));
   XNOR2_X1 i_0_115 (.A(in3[19]), .B(in1[19]), .ZN(n_0_71));
   XNOR2_X1 i_0_116 (.A(in2[20]), .B(n_0_72), .ZN(sum[20]));
   XNOR2_X1 i_0_117 (.A(in3[20]), .B(in1[20]), .ZN(n_0_72));
   XNOR2_X1 i_0_118 (.A(in2[21]), .B(n_0_73), .ZN(sum[21]));
   XNOR2_X1 i_0_119 (.A(in3[21]), .B(in1[21]), .ZN(n_0_73));
   XNOR2_X1 i_0_120 (.A(in2[22]), .B(n_0_74), .ZN(sum[22]));
   XNOR2_X1 i_0_121 (.A(in3[22]), .B(in1[22]), .ZN(n_0_74));
   XNOR2_X1 i_0_122 (.A(in2[23]), .B(n_0_75), .ZN(sum[23]));
   XNOR2_X1 i_0_123 (.A(in3[23]), .B(in1[23]), .ZN(n_0_75));
   XNOR2_X1 i_0_124 (.A(in2[24]), .B(n_0_76), .ZN(sum[24]));
   XNOR2_X1 i_0_125 (.A(in3[24]), .B(in1[24]), .ZN(n_0_76));
   XNOR2_X1 i_0_126 (.A(in2[25]), .B(n_0_77), .ZN(sum[25]));
   XNOR2_X1 i_0_127 (.A(in3[25]), .B(in1[25]), .ZN(n_0_77));
   XNOR2_X1 i_0_128 (.A(in2[26]), .B(n_0_78), .ZN(sum[26]));
   XNOR2_X1 i_0_129 (.A(in3[26]), .B(in1[26]), .ZN(n_0_78));
   XNOR2_X1 i_0_130 (.A(in2[27]), .B(n_0_79), .ZN(sum[27]));
   XNOR2_X1 i_0_131 (.A(in3[27]), .B(in1[27]), .ZN(n_0_79));
   XNOR2_X1 i_0_132 (.A(in2[28]), .B(n_0_80), .ZN(sum[28]));
   XNOR2_X1 i_0_133 (.A(in3[28]), .B(in1[28]), .ZN(n_0_80));
   XNOR2_X1 i_0_134 (.A(in2[29]), .B(n_0_81), .ZN(sum[29]));
   XNOR2_X1 i_0_135 (.A(in3[29]), .B(in1[29]), .ZN(n_0_81));
   XNOR2_X1 i_0_136 (.A(in2[30]), .B(n_0_82), .ZN(sum[30]));
   XNOR2_X1 i_0_137 (.A(in3[30]), .B(in1[30]), .ZN(n_0_82));
   XNOR2_X1 i_0_138 (.A(in2[31]), .B(n_0_83), .ZN(sum[31]));
   XNOR2_X1 i_0_139 (.A(in3[31]), .B(in1[31]), .ZN(n_0_83));
   XNOR2_X1 i_0_140 (.A(in2[32]), .B(n_0_84), .ZN(sum[32]));
   XNOR2_X1 i_0_141 (.A(in3[32]), .B(in1[32]), .ZN(n_0_84));
   XNOR2_X1 i_0_142 (.A(in2[33]), .B(n_0_85), .ZN(sum[33]));
   XNOR2_X1 i_0_143 (.A(in3[33]), .B(in1[33]), .ZN(n_0_85));
   XNOR2_X1 i_0_144 (.A(in2[34]), .B(n_0_86), .ZN(sum[34]));
   XNOR2_X1 i_0_145 (.A(in3[34]), .B(in1[34]), .ZN(n_0_86));
   XNOR2_X1 i_0_146 (.A(in2[35]), .B(n_0_87), .ZN(sum[35]));
   XNOR2_X1 i_0_147 (.A(in3[35]), .B(in1[35]), .ZN(n_0_87));
   XNOR2_X1 i_0_148 (.A(in2[36]), .B(n_0_88), .ZN(sum[36]));
   XNOR2_X1 i_0_149 (.A(in3[36]), .B(in1[36]), .ZN(n_0_88));
   XNOR2_X1 i_0_150 (.A(in2[37]), .B(n_0_89), .ZN(sum[37]));
   XNOR2_X1 i_0_151 (.A(in3[37]), .B(in1[37]), .ZN(n_0_89));
   XNOR2_X1 i_0_152 (.A(in2[38]), .B(n_0_90), .ZN(sum[38]));
   XNOR2_X1 i_0_153 (.A(in3[38]), .B(in1[38]), .ZN(n_0_90));
   XNOR2_X1 i_0_154 (.A(in2[39]), .B(n_0_91), .ZN(sum[39]));
   XNOR2_X1 i_0_155 (.A(in3[39]), .B(in1[39]), .ZN(n_0_91));
   XNOR2_X1 i_0_156 (.A(in2[40]), .B(n_0_92), .ZN(sum[40]));
   XNOR2_X1 i_0_157 (.A(in3[40]), .B(in1[40]), .ZN(n_0_92));
   XNOR2_X1 i_0_158 (.A(in2[41]), .B(n_0_93), .ZN(sum[41]));
   XNOR2_X1 i_0_159 (.A(in3[41]), .B(in1[41]), .ZN(n_0_93));
   XNOR2_X1 i_0_160 (.A(in2[42]), .B(n_0_94), .ZN(sum[42]));
   XNOR2_X1 i_0_161 (.A(in3[42]), .B(in1[63]), .ZN(n_0_94));
   XNOR2_X1 i_0_162 (.A(n_0_96), .B(n_0_95), .ZN(sum[43]));
   XNOR2_X1 i_0_163 (.A(n_0_97), .B(n_0_95), .ZN(sum[44]));
   XNOR2_X1 i_0_164 (.A(n_0_98), .B(n_0_95), .ZN(sum[63]));
   XOR2_X1 i_0_165 (.A(in2[63]), .B(in1[63]), .Z(n_0_95));
   INV_X1 i_0_166 (.A(in3[43]), .ZN(n_0_96));
   INV_X1 i_0_167 (.A(in3[44]), .ZN(n_0_97));
   INV_X1 i_0_168 (.A(in3[63]), .ZN(n_0_98));
endmodule

module CSA__1_29(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;

   AND2_X1 i_0_0 (.A1(in2[9]), .A2(in1[9]), .ZN(c[10]));
   AND2_X1 i_0_1 (.A1(in2[10]), .A2(in1[10]), .ZN(c[11]));
   AND2_X1 i_0_2 (.A1(in2[11]), .A2(in1[11]), .ZN(c[12]));
   NAND2_X1 i_0_3 (.A1(n_0_1), .A2(n_0_0), .ZN(c[13]));
   OAI21_X1 i_0_4 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_0));
   NAND2_X1 i_0_5 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_1));
   NAND2_X1 i_0_6 (.A1(n_0_3), .A2(n_0_2), .ZN(c[14]));
   OAI21_X1 i_0_7 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_2));
   NAND2_X1 i_0_8 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_3));
   NAND2_X1 i_0_9 (.A1(n_0_5), .A2(n_0_4), .ZN(c[15]));
   OAI21_X1 i_0_10 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_4));
   NAND2_X1 i_0_11 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_5));
   NAND2_X1 i_0_12 (.A1(n_0_7), .A2(n_0_6), .ZN(c[16]));
   OAI21_X1 i_0_13 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_6));
   NAND2_X1 i_0_14 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_7));
   NAND2_X1 i_0_15 (.A1(n_0_9), .A2(n_0_8), .ZN(c[17]));
   OAI21_X1 i_0_16 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_8));
   NAND2_X1 i_0_17 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_9));
   NAND2_X1 i_0_18 (.A1(n_0_11), .A2(n_0_10), .ZN(c[18]));
   OAI21_X1 i_0_19 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_10));
   NAND2_X1 i_0_20 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_11));
   NAND2_X1 i_0_21 (.A1(n_0_13), .A2(n_0_12), .ZN(c[19]));
   OAI21_X1 i_0_22 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_12));
   NAND2_X1 i_0_23 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_13));
   NAND2_X1 i_0_24 (.A1(n_0_15), .A2(n_0_14), .ZN(c[20]));
   OAI21_X1 i_0_25 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_14));
   NAND2_X1 i_0_26 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_15));
   NAND2_X1 i_0_27 (.A1(n_0_17), .A2(n_0_16), .ZN(c[21]));
   OAI21_X1 i_0_28 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_16));
   NAND2_X1 i_0_29 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_17));
   NAND2_X1 i_0_30 (.A1(n_0_19), .A2(n_0_18), .ZN(c[22]));
   OAI21_X1 i_0_31 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_18));
   NAND2_X1 i_0_32 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_19));
   NAND2_X1 i_0_33 (.A1(n_0_21), .A2(n_0_20), .ZN(c[23]));
   OAI21_X1 i_0_34 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_20));
   NAND2_X1 i_0_35 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_21));
   NAND2_X1 i_0_36 (.A1(n_0_23), .A2(n_0_22), .ZN(c[24]));
   OAI21_X1 i_0_37 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_22));
   NAND2_X1 i_0_38 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_23));
   NAND2_X1 i_0_39 (.A1(n_0_25), .A2(n_0_24), .ZN(c[25]));
   OAI21_X1 i_0_40 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_24));
   NAND2_X1 i_0_41 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_25));
   NAND2_X1 i_0_42 (.A1(n_0_27), .A2(n_0_26), .ZN(c[26]));
   OAI21_X1 i_0_43 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_26));
   NAND2_X1 i_0_44 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_27));
   NAND2_X1 i_0_45 (.A1(n_0_29), .A2(n_0_28), .ZN(c[27]));
   OAI21_X1 i_0_46 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_28));
   NAND2_X1 i_0_47 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_29));
   NAND2_X1 i_0_48 (.A1(n_0_31), .A2(n_0_30), .ZN(c[28]));
   OAI21_X1 i_0_49 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_30));
   NAND2_X1 i_0_50 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_31));
   NAND2_X1 i_0_51 (.A1(n_0_33), .A2(n_0_32), .ZN(c[29]));
   OAI21_X1 i_0_52 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_32));
   NAND2_X1 i_0_53 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_33));
   NAND2_X1 i_0_54 (.A1(n_0_35), .A2(n_0_34), .ZN(c[30]));
   OAI21_X1 i_0_55 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_34));
   NAND2_X1 i_0_56 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_35));
   NAND2_X1 i_0_57 (.A1(n_0_37), .A2(n_0_36), .ZN(c[31]));
   OAI21_X1 i_0_58 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_36));
   NAND2_X1 i_0_59 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_37));
   NAND2_X1 i_0_60 (.A1(n_0_39), .A2(n_0_38), .ZN(c[32]));
   OAI21_X1 i_0_61 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_38));
   NAND2_X1 i_0_62 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_39));
   NAND2_X1 i_0_63 (.A1(n_0_41), .A2(n_0_40), .ZN(c[33]));
   OAI21_X1 i_0_64 (.A(in3[32]), .B1(in1[32]), .B2(in2[32]), .ZN(n_0_40));
   NAND2_X1 i_0_65 (.A1(in2[32]), .A2(in1[32]), .ZN(n_0_41));
   NAND2_X1 i_0_66 (.A1(n_0_43), .A2(n_0_42), .ZN(c[34]));
   OAI21_X1 i_0_67 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_42));
   NAND2_X1 i_0_68 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_43));
   NAND2_X1 i_0_69 (.A1(n_0_45), .A2(n_0_44), .ZN(c[35]));
   OAI21_X1 i_0_70 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_44));
   NAND2_X1 i_0_71 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_45));
   NAND2_X1 i_0_72 (.A1(n_0_47), .A2(n_0_46), .ZN(c[36]));
   OAI21_X1 i_0_73 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_46));
   NAND2_X1 i_0_74 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_47));
   NAND2_X1 i_0_75 (.A1(n_0_49), .A2(n_0_48), .ZN(c[37]));
   OAI21_X1 i_0_76 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_48));
   NAND2_X1 i_0_77 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_49));
   NAND2_X1 i_0_78 (.A1(n_0_51), .A2(n_0_50), .ZN(c[38]));
   OAI21_X1 i_0_79 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_50));
   NAND2_X1 i_0_80 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_51));
   NAND2_X1 i_0_81 (.A1(n_0_53), .A2(n_0_52), .ZN(c[39]));
   OAI21_X1 i_0_82 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_52));
   NAND2_X1 i_0_83 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_53));
   NAND2_X1 i_0_84 (.A1(n_0_55), .A2(n_0_54), .ZN(c[40]));
   OAI21_X1 i_0_85 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_54));
   NAND2_X1 i_0_86 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_55));
   NAND2_X1 i_0_87 (.A1(n_0_57), .A2(n_0_56), .ZN(c[41]));
   OAI21_X1 i_0_88 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_56));
   NAND2_X1 i_0_89 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_57));
   NAND2_X1 i_0_90 (.A1(n_0_59), .A2(n_0_58), .ZN(c[42]));
   OAI21_X1 i_0_91 (.A(in2[41]), .B1(in3[41]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_92 (.A1(in3[41]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_93 (.A1(n_0_61), .A2(n_0_60), .ZN(c[43]));
   OAI21_X1 i_0_94 (.A(in2[42]), .B1(in3[42]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_95 (.A1(in3[42]), .A2(in1[63]), .ZN(n_0_61));
   NAND2_X1 i_0_96 (.A1(n_0_63), .A2(n_0_62), .ZN(c[44]));
   OAI21_X1 i_0_97 (.A(in2[43]), .B1(in3[43]), .B2(in1[63]), .ZN(n_0_62));
   NAND2_X1 i_0_98 (.A1(in3[43]), .A2(in1[63]), .ZN(n_0_63));
   NAND2_X1 i_0_99 (.A1(n_0_65), .A2(n_0_64), .ZN(c[45]));
   OAI21_X1 i_0_100 (.A(in2[44]), .B1(in3[44]), .B2(in1[63]), .ZN(n_0_64));
   NAND2_X1 i_0_101 (.A1(in3[44]), .A2(in1[63]), .ZN(n_0_65));
   NAND2_X1 i_0_102 (.A1(n_0_68), .A2(n_0_66), .ZN(c[46]));
   OAI21_X1 i_0_103 (.A(in3[45]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_66));
   NAND2_X1 i_0_104 (.A1(n_0_68), .A2(n_0_67), .ZN(c[63]));
   OAI21_X1 i_0_105 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_67));
   NAND2_X1 i_0_106 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_68));
   XOR2_X1 i_0_107 (.A(in2[9]), .B(in1[9]), .Z(sum[9]));
   XOR2_X1 i_0_108 (.A(in2[10]), .B(in1[10]), .Z(sum[10]));
   XOR2_X1 i_0_109 (.A(in2[11]), .B(in1[11]), .Z(sum[11]));
   XNOR2_X1 i_0_110 (.A(in2[12]), .B(n_0_69), .ZN(sum[12]));
   XNOR2_X1 i_0_111 (.A(in3[12]), .B(in1[12]), .ZN(n_0_69));
   XNOR2_X1 i_0_112 (.A(in2[13]), .B(n_0_70), .ZN(sum[13]));
   XNOR2_X1 i_0_113 (.A(in3[13]), .B(in1[13]), .ZN(n_0_70));
   XNOR2_X1 i_0_114 (.A(in2[14]), .B(n_0_71), .ZN(sum[14]));
   XNOR2_X1 i_0_115 (.A(in3[14]), .B(in1[14]), .ZN(n_0_71));
   XNOR2_X1 i_0_116 (.A(in2[15]), .B(n_0_72), .ZN(sum[15]));
   XNOR2_X1 i_0_117 (.A(in3[15]), .B(in1[15]), .ZN(n_0_72));
   XNOR2_X1 i_0_118 (.A(in2[16]), .B(n_0_73), .ZN(sum[16]));
   XNOR2_X1 i_0_119 (.A(in3[16]), .B(in1[16]), .ZN(n_0_73));
   XNOR2_X1 i_0_120 (.A(in2[17]), .B(n_0_74), .ZN(sum[17]));
   XNOR2_X1 i_0_121 (.A(in3[17]), .B(in1[17]), .ZN(n_0_74));
   XNOR2_X1 i_0_122 (.A(in2[18]), .B(n_0_75), .ZN(sum[18]));
   XNOR2_X1 i_0_123 (.A(in3[18]), .B(in1[18]), .ZN(n_0_75));
   XNOR2_X1 i_0_124 (.A(in2[19]), .B(n_0_76), .ZN(sum[19]));
   XNOR2_X1 i_0_125 (.A(in3[19]), .B(in1[19]), .ZN(n_0_76));
   XNOR2_X1 i_0_126 (.A(in2[20]), .B(n_0_77), .ZN(sum[20]));
   XNOR2_X1 i_0_127 (.A(in3[20]), .B(in1[20]), .ZN(n_0_77));
   XNOR2_X1 i_0_128 (.A(in2[21]), .B(n_0_78), .ZN(sum[21]));
   XNOR2_X1 i_0_129 (.A(in3[21]), .B(in1[21]), .ZN(n_0_78));
   XNOR2_X1 i_0_130 (.A(in2[22]), .B(n_0_79), .ZN(sum[22]));
   XNOR2_X1 i_0_131 (.A(in3[22]), .B(in1[22]), .ZN(n_0_79));
   XNOR2_X1 i_0_132 (.A(in2[23]), .B(n_0_80), .ZN(sum[23]));
   XNOR2_X1 i_0_133 (.A(in3[23]), .B(in1[23]), .ZN(n_0_80));
   XNOR2_X1 i_0_134 (.A(in2[24]), .B(n_0_81), .ZN(sum[24]));
   XNOR2_X1 i_0_135 (.A(in3[24]), .B(in1[24]), .ZN(n_0_81));
   XNOR2_X1 i_0_136 (.A(in2[25]), .B(n_0_82), .ZN(sum[25]));
   XNOR2_X1 i_0_137 (.A(in3[25]), .B(in1[25]), .ZN(n_0_82));
   XNOR2_X1 i_0_138 (.A(in2[26]), .B(n_0_83), .ZN(sum[26]));
   XNOR2_X1 i_0_139 (.A(in3[26]), .B(in1[26]), .ZN(n_0_83));
   XNOR2_X1 i_0_140 (.A(in2[27]), .B(n_0_84), .ZN(sum[27]));
   XNOR2_X1 i_0_141 (.A(in3[27]), .B(in1[27]), .ZN(n_0_84));
   XNOR2_X1 i_0_142 (.A(in2[28]), .B(n_0_85), .ZN(sum[28]));
   XNOR2_X1 i_0_143 (.A(in3[28]), .B(in1[28]), .ZN(n_0_85));
   XNOR2_X1 i_0_144 (.A(in2[29]), .B(n_0_86), .ZN(sum[29]));
   XNOR2_X1 i_0_145 (.A(in3[29]), .B(in1[29]), .ZN(n_0_86));
   XNOR2_X1 i_0_146 (.A(in2[30]), .B(n_0_87), .ZN(sum[30]));
   XNOR2_X1 i_0_147 (.A(in3[30]), .B(in1[30]), .ZN(n_0_87));
   XNOR2_X1 i_0_148 (.A(in2[31]), .B(n_0_88), .ZN(sum[31]));
   XNOR2_X1 i_0_149 (.A(in3[31]), .B(in1[31]), .ZN(n_0_88));
   XNOR2_X1 i_0_150 (.A(in2[32]), .B(n_0_89), .ZN(sum[32]));
   XNOR2_X1 i_0_151 (.A(in3[32]), .B(in1[32]), .ZN(n_0_89));
   XNOR2_X1 i_0_152 (.A(in2[33]), .B(n_0_90), .ZN(sum[33]));
   XNOR2_X1 i_0_153 (.A(in3[33]), .B(in1[33]), .ZN(n_0_90));
   XNOR2_X1 i_0_154 (.A(in2[34]), .B(n_0_91), .ZN(sum[34]));
   XNOR2_X1 i_0_155 (.A(in3[34]), .B(in1[34]), .ZN(n_0_91));
   XNOR2_X1 i_0_156 (.A(in2[35]), .B(n_0_92), .ZN(sum[35]));
   XNOR2_X1 i_0_157 (.A(in3[35]), .B(in1[35]), .ZN(n_0_92));
   XNOR2_X1 i_0_158 (.A(in2[36]), .B(n_0_93), .ZN(sum[36]));
   XNOR2_X1 i_0_159 (.A(in3[36]), .B(in1[36]), .ZN(n_0_93));
   XNOR2_X1 i_0_160 (.A(in2[37]), .B(n_0_94), .ZN(sum[37]));
   XNOR2_X1 i_0_161 (.A(in3[37]), .B(in1[37]), .ZN(n_0_94));
   XNOR2_X1 i_0_162 (.A(in2[38]), .B(n_0_95), .ZN(sum[38]));
   XNOR2_X1 i_0_163 (.A(in3[38]), .B(in1[38]), .ZN(n_0_95));
   XNOR2_X1 i_0_164 (.A(in2[39]), .B(n_0_96), .ZN(sum[39]));
   XNOR2_X1 i_0_165 (.A(in3[39]), .B(in1[39]), .ZN(n_0_96));
   XNOR2_X1 i_0_166 (.A(in2[40]), .B(n_0_97), .ZN(sum[40]));
   XNOR2_X1 i_0_167 (.A(in3[40]), .B(in1[40]), .ZN(n_0_97));
   XNOR2_X1 i_0_168 (.A(in2[41]), .B(n_0_98), .ZN(sum[41]));
   XNOR2_X1 i_0_169 (.A(in3[41]), .B(in1[63]), .ZN(n_0_98));
   XNOR2_X1 i_0_170 (.A(in2[42]), .B(n_0_99), .ZN(sum[42]));
   XNOR2_X1 i_0_171 (.A(in3[42]), .B(in1[63]), .ZN(n_0_99));
   XNOR2_X1 i_0_172 (.A(in2[43]), .B(n_0_100), .ZN(sum[43]));
   XNOR2_X1 i_0_173 (.A(in3[43]), .B(in1[63]), .ZN(n_0_100));
   XNOR2_X1 i_0_174 (.A(in2[44]), .B(n_0_101), .ZN(sum[44]));
   XNOR2_X1 i_0_175 (.A(in3[44]), .B(in1[63]), .ZN(n_0_101));
   XOR2_X1 i_0_176 (.A(in3[45]), .B(n_0_102), .Z(sum[45]));
   XOR2_X1 i_0_177 (.A(in3[63]), .B(n_0_102), .Z(sum[63]));
   XOR2_X1 i_0_178 (.A(in2[63]), .B(in1[63]), .Z(n_0_102));
endmodule

module CSA__1_32(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;

   AND2_X1 i_0_0 (.A1(in2[4]), .A2(in1[4]), .ZN(c[5]));
   AND2_X1 i_0_1 (.A1(in2[5]), .A2(in1[5]), .ZN(c[6]));
   AND2_X1 i_0_2 (.A1(in2[6]), .A2(in1[6]), .ZN(c[7]));
   NAND2_X1 i_0_3 (.A1(n_0_1), .A2(n_0_0), .ZN(c[8]));
   OAI21_X1 i_0_4 (.A(in2[7]), .B1(in3[7]), .B2(in1[7]), .ZN(n_0_0));
   NAND2_X1 i_0_5 (.A1(in3[7]), .A2(in1[7]), .ZN(n_0_1));
   NAND2_X1 i_0_6 (.A1(n_0_3), .A2(n_0_2), .ZN(c[9]));
   OAI21_X1 i_0_7 (.A(in2[8]), .B1(in3[8]), .B2(in1[8]), .ZN(n_0_2));
   NAND2_X1 i_0_8 (.A1(in3[8]), .A2(in1[8]), .ZN(n_0_3));
   NAND2_X1 i_0_9 (.A1(n_0_5), .A2(n_0_4), .ZN(c[10]));
   OAI21_X1 i_0_10 (.A(in2[9]), .B1(in3[9]), .B2(in1[9]), .ZN(n_0_4));
   NAND2_X1 i_0_11 (.A1(in3[9]), .A2(in1[9]), .ZN(n_0_5));
   NAND2_X1 i_0_12 (.A1(n_0_7), .A2(n_0_6), .ZN(c[11]));
   OAI21_X1 i_0_13 (.A(in2[10]), .B1(in3[10]), .B2(in1[10]), .ZN(n_0_6));
   NAND2_X1 i_0_14 (.A1(in3[10]), .A2(in1[10]), .ZN(n_0_7));
   NAND2_X1 i_0_15 (.A1(n_0_9), .A2(n_0_8), .ZN(c[12]));
   OAI21_X1 i_0_16 (.A(in2[11]), .B1(in3[11]), .B2(in1[11]), .ZN(n_0_8));
   NAND2_X1 i_0_17 (.A1(in3[11]), .A2(in1[11]), .ZN(n_0_9));
   NAND2_X1 i_0_18 (.A1(n_0_11), .A2(n_0_10), .ZN(c[13]));
   OAI21_X1 i_0_19 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_10));
   NAND2_X1 i_0_20 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_11));
   NAND2_X1 i_0_21 (.A1(n_0_13), .A2(n_0_12), .ZN(c[14]));
   OAI21_X1 i_0_22 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_12));
   NAND2_X1 i_0_23 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_13));
   NAND2_X1 i_0_24 (.A1(n_0_15), .A2(n_0_14), .ZN(c[15]));
   OAI21_X1 i_0_25 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_14));
   NAND2_X1 i_0_26 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_15));
   NAND2_X1 i_0_27 (.A1(n_0_17), .A2(n_0_16), .ZN(c[16]));
   OAI21_X1 i_0_28 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_16));
   NAND2_X1 i_0_29 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_17));
   NAND2_X1 i_0_30 (.A1(n_0_19), .A2(n_0_18), .ZN(c[17]));
   OAI21_X1 i_0_31 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_18));
   NAND2_X1 i_0_32 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_19));
   NAND2_X1 i_0_33 (.A1(n_0_21), .A2(n_0_20), .ZN(c[18]));
   OAI21_X1 i_0_34 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_20));
   NAND2_X1 i_0_35 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_21));
   NAND2_X1 i_0_36 (.A1(n_0_23), .A2(n_0_22), .ZN(c[19]));
   OAI21_X1 i_0_37 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_22));
   NAND2_X1 i_0_38 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_23));
   NAND2_X1 i_0_39 (.A1(n_0_25), .A2(n_0_24), .ZN(c[20]));
   OAI21_X1 i_0_40 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_24));
   NAND2_X1 i_0_41 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_25));
   NAND2_X1 i_0_42 (.A1(n_0_27), .A2(n_0_26), .ZN(c[21]));
   OAI21_X1 i_0_43 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_26));
   NAND2_X1 i_0_44 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_27));
   NAND2_X1 i_0_45 (.A1(n_0_29), .A2(n_0_28), .ZN(c[22]));
   OAI21_X1 i_0_46 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_28));
   NAND2_X1 i_0_47 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_29));
   NAND2_X1 i_0_48 (.A1(n_0_31), .A2(n_0_30), .ZN(c[23]));
   OAI21_X1 i_0_49 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_30));
   NAND2_X1 i_0_50 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_31));
   NAND2_X1 i_0_51 (.A1(n_0_33), .A2(n_0_32), .ZN(c[24]));
   OAI21_X1 i_0_52 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_32));
   NAND2_X1 i_0_53 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_33));
   NAND2_X1 i_0_54 (.A1(n_0_35), .A2(n_0_34), .ZN(c[25]));
   OAI21_X1 i_0_55 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_34));
   NAND2_X1 i_0_56 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_35));
   NAND2_X1 i_0_57 (.A1(n_0_37), .A2(n_0_36), .ZN(c[26]));
   OAI21_X1 i_0_58 (.A(in3[25]), .B1(in1[25]), .B2(in2[25]), .ZN(n_0_36));
   NAND2_X1 i_0_59 (.A1(in2[25]), .A2(in1[25]), .ZN(n_0_37));
   NAND2_X1 i_0_60 (.A1(n_0_39), .A2(n_0_38), .ZN(c[27]));
   OAI21_X1 i_0_61 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_38));
   NAND2_X1 i_0_62 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_39));
   NAND2_X1 i_0_63 (.A1(n_0_41), .A2(n_0_40), .ZN(c[28]));
   OAI21_X1 i_0_64 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_40));
   NAND2_X1 i_0_65 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_41));
   NAND2_X1 i_0_66 (.A1(n_0_43), .A2(n_0_42), .ZN(c[29]));
   OAI21_X1 i_0_67 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_42));
   NAND2_X1 i_0_68 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_43));
   NAND2_X1 i_0_69 (.A1(n_0_45), .A2(n_0_44), .ZN(c[30]));
   OAI21_X1 i_0_70 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_44));
   NAND2_X1 i_0_71 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_45));
   NAND2_X1 i_0_72 (.A1(n_0_47), .A2(n_0_46), .ZN(c[31]));
   OAI21_X1 i_0_73 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_46));
   NAND2_X1 i_0_74 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_47));
   NAND2_X1 i_0_75 (.A1(n_0_49), .A2(n_0_48), .ZN(c[32]));
   OAI21_X1 i_0_76 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_48));
   NAND2_X1 i_0_77 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_49));
   NAND2_X1 i_0_78 (.A1(n_0_51), .A2(n_0_50), .ZN(c[33]));
   OAI21_X1 i_0_79 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_50));
   NAND2_X1 i_0_80 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_51));
   NAND2_X1 i_0_81 (.A1(n_0_53), .A2(n_0_52), .ZN(c[34]));
   OAI21_X1 i_0_82 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_52));
   NAND2_X1 i_0_83 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_53));
   NAND2_X1 i_0_84 (.A1(n_0_55), .A2(n_0_54), .ZN(c[35]));
   OAI21_X1 i_0_85 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_54));
   NAND2_X1 i_0_86 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_55));
   NAND2_X1 i_0_87 (.A1(n_0_57), .A2(n_0_56), .ZN(c[36]));
   OAI21_X1 i_0_88 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_56));
   NAND2_X1 i_0_89 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_57));
   NAND2_X1 i_0_90 (.A1(n_0_59), .A2(n_0_58), .ZN(c[37]));
   OAI21_X1 i_0_91 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_58));
   NAND2_X1 i_0_92 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_59));
   NAND2_X1 i_0_93 (.A1(n_0_61), .A2(n_0_60), .ZN(c[38]));
   OAI21_X1 i_0_94 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_60));
   NAND2_X1 i_0_95 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_61));
   NAND2_X1 i_0_96 (.A1(n_0_63), .A2(n_0_62), .ZN(c[39]));
   OAI21_X1 i_0_97 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_62));
   NAND2_X1 i_0_98 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_63));
   NAND2_X1 i_0_99 (.A1(n_0_65), .A2(n_0_64), .ZN(c[40]));
   OAI21_X1 i_0_100 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_64));
   NAND2_X1 i_0_101 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_65));
   NAND2_X1 i_0_102 (.A1(n_0_67), .A2(n_0_66), .ZN(c[41]));
   OAI21_X1 i_0_103 (.A(in2[40]), .B1(in3[40]), .B2(in1[63]), .ZN(n_0_66));
   NAND2_X1 i_0_104 (.A1(in3[40]), .A2(in1[63]), .ZN(n_0_67));
   AOI21_X1 i_0_105 (.A(n_0_69), .B1(n_0_68), .B2(n_0_105), .ZN(c[42]));
   AOI21_X1 i_0_106 (.A(n_0_69), .B1(n_0_68), .B2(n_0_106), .ZN(c[43]));
   AOI21_X1 i_0_107 (.A(n_0_69), .B1(n_0_68), .B2(n_0_107), .ZN(c[44]));
   AOI21_X1 i_0_108 (.A(n_0_69), .B1(n_0_68), .B2(n_0_108), .ZN(c[45]));
   AOI21_X1 i_0_109 (.A(n_0_69), .B1(n_0_68), .B2(n_0_109), .ZN(c[46]));
   AOI21_X1 i_0_110 (.A(n_0_69), .B1(n_0_68), .B2(n_0_110), .ZN(c[63]));
   NAND2_X1 i_0_111 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_68));
   NOR2_X1 i_0_112 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_69));
   XOR2_X1 i_0_113 (.A(in2[4]), .B(in1[4]), .Z(sum[4]));
   XOR2_X1 i_0_114 (.A(in2[5]), .B(in1[5]), .Z(sum[5]));
   XOR2_X1 i_0_115 (.A(in2[6]), .B(in1[6]), .Z(sum[6]));
   XNOR2_X1 i_0_116 (.A(in2[7]), .B(n_0_70), .ZN(sum[7]));
   XNOR2_X1 i_0_117 (.A(in3[7]), .B(in1[7]), .ZN(n_0_70));
   XNOR2_X1 i_0_118 (.A(in2[8]), .B(n_0_71), .ZN(sum[8]));
   XNOR2_X1 i_0_119 (.A(in3[8]), .B(in1[8]), .ZN(n_0_71));
   XNOR2_X1 i_0_120 (.A(in2[9]), .B(n_0_72), .ZN(sum[9]));
   XNOR2_X1 i_0_121 (.A(in3[9]), .B(in1[9]), .ZN(n_0_72));
   XNOR2_X1 i_0_122 (.A(in2[10]), .B(n_0_73), .ZN(sum[10]));
   XNOR2_X1 i_0_123 (.A(in3[10]), .B(in1[10]), .ZN(n_0_73));
   XNOR2_X1 i_0_124 (.A(in2[11]), .B(n_0_74), .ZN(sum[11]));
   XNOR2_X1 i_0_125 (.A(in3[11]), .B(in1[11]), .ZN(n_0_74));
   XNOR2_X1 i_0_126 (.A(in2[12]), .B(n_0_75), .ZN(sum[12]));
   XNOR2_X1 i_0_127 (.A(in3[12]), .B(in1[12]), .ZN(n_0_75));
   XNOR2_X1 i_0_128 (.A(in2[13]), .B(n_0_76), .ZN(sum[13]));
   XNOR2_X1 i_0_129 (.A(in3[13]), .B(in1[13]), .ZN(n_0_76));
   XNOR2_X1 i_0_130 (.A(in2[14]), .B(n_0_77), .ZN(sum[14]));
   XNOR2_X1 i_0_131 (.A(in3[14]), .B(in1[14]), .ZN(n_0_77));
   XNOR2_X1 i_0_132 (.A(in2[15]), .B(n_0_78), .ZN(sum[15]));
   XNOR2_X1 i_0_133 (.A(in3[15]), .B(in1[15]), .ZN(n_0_78));
   XNOR2_X1 i_0_134 (.A(in2[16]), .B(n_0_79), .ZN(sum[16]));
   XNOR2_X1 i_0_135 (.A(in3[16]), .B(in1[16]), .ZN(n_0_79));
   XNOR2_X1 i_0_136 (.A(in2[17]), .B(n_0_80), .ZN(sum[17]));
   XNOR2_X1 i_0_137 (.A(in3[17]), .B(in1[17]), .ZN(n_0_80));
   XNOR2_X1 i_0_138 (.A(in2[18]), .B(n_0_81), .ZN(sum[18]));
   XNOR2_X1 i_0_139 (.A(in3[18]), .B(in1[18]), .ZN(n_0_81));
   XNOR2_X1 i_0_140 (.A(in2[19]), .B(n_0_82), .ZN(sum[19]));
   XNOR2_X1 i_0_141 (.A(in3[19]), .B(in1[19]), .ZN(n_0_82));
   XNOR2_X1 i_0_142 (.A(in2[20]), .B(n_0_83), .ZN(sum[20]));
   XNOR2_X1 i_0_143 (.A(in3[20]), .B(in1[20]), .ZN(n_0_83));
   XNOR2_X1 i_0_144 (.A(in2[21]), .B(n_0_84), .ZN(sum[21]));
   XNOR2_X1 i_0_145 (.A(in3[21]), .B(in1[21]), .ZN(n_0_84));
   XNOR2_X1 i_0_146 (.A(in2[22]), .B(n_0_85), .ZN(sum[22]));
   XNOR2_X1 i_0_147 (.A(in3[22]), .B(in1[22]), .ZN(n_0_85));
   XNOR2_X1 i_0_148 (.A(in2[23]), .B(n_0_86), .ZN(sum[23]));
   XNOR2_X1 i_0_149 (.A(in3[23]), .B(in1[23]), .ZN(n_0_86));
   XNOR2_X1 i_0_150 (.A(in2[24]), .B(n_0_87), .ZN(sum[24]));
   XNOR2_X1 i_0_151 (.A(in3[24]), .B(in1[24]), .ZN(n_0_87));
   XNOR2_X1 i_0_152 (.A(in2[25]), .B(n_0_88), .ZN(sum[25]));
   XNOR2_X1 i_0_153 (.A(in3[25]), .B(in1[25]), .ZN(n_0_88));
   XNOR2_X1 i_0_154 (.A(in2[26]), .B(n_0_89), .ZN(sum[26]));
   XNOR2_X1 i_0_155 (.A(in3[26]), .B(in1[26]), .ZN(n_0_89));
   XNOR2_X1 i_0_156 (.A(in2[27]), .B(n_0_90), .ZN(sum[27]));
   XNOR2_X1 i_0_157 (.A(in3[27]), .B(in1[27]), .ZN(n_0_90));
   XNOR2_X1 i_0_158 (.A(in2[28]), .B(n_0_91), .ZN(sum[28]));
   XNOR2_X1 i_0_159 (.A(in3[28]), .B(in1[28]), .ZN(n_0_91));
   XNOR2_X1 i_0_160 (.A(in2[29]), .B(n_0_92), .ZN(sum[29]));
   XNOR2_X1 i_0_161 (.A(in3[29]), .B(in1[29]), .ZN(n_0_92));
   XNOR2_X1 i_0_162 (.A(in2[30]), .B(n_0_93), .ZN(sum[30]));
   XNOR2_X1 i_0_163 (.A(in3[30]), .B(in1[30]), .ZN(n_0_93));
   XNOR2_X1 i_0_164 (.A(in2[31]), .B(n_0_94), .ZN(sum[31]));
   XNOR2_X1 i_0_165 (.A(in3[31]), .B(in1[31]), .ZN(n_0_94));
   XNOR2_X1 i_0_166 (.A(in2[32]), .B(n_0_95), .ZN(sum[32]));
   XNOR2_X1 i_0_167 (.A(in3[32]), .B(in1[32]), .ZN(n_0_95));
   XNOR2_X1 i_0_168 (.A(in2[33]), .B(n_0_96), .ZN(sum[33]));
   XNOR2_X1 i_0_169 (.A(in3[33]), .B(in1[33]), .ZN(n_0_96));
   XNOR2_X1 i_0_170 (.A(in2[34]), .B(n_0_97), .ZN(sum[34]));
   XNOR2_X1 i_0_171 (.A(in3[34]), .B(in1[34]), .ZN(n_0_97));
   XNOR2_X1 i_0_172 (.A(in2[35]), .B(n_0_98), .ZN(sum[35]));
   XNOR2_X1 i_0_173 (.A(in3[35]), .B(in1[35]), .ZN(n_0_98));
   XNOR2_X1 i_0_174 (.A(in2[36]), .B(n_0_99), .ZN(sum[36]));
   XNOR2_X1 i_0_175 (.A(in3[36]), .B(in1[36]), .ZN(n_0_99));
   XNOR2_X1 i_0_176 (.A(in2[37]), .B(n_0_100), .ZN(sum[37]));
   XNOR2_X1 i_0_177 (.A(in3[37]), .B(in1[37]), .ZN(n_0_100));
   XNOR2_X1 i_0_178 (.A(in2[38]), .B(n_0_101), .ZN(sum[38]));
   XNOR2_X1 i_0_179 (.A(in3[38]), .B(in1[38]), .ZN(n_0_101));
   XNOR2_X1 i_0_180 (.A(in2[39]), .B(n_0_102), .ZN(sum[39]));
   XNOR2_X1 i_0_181 (.A(in3[39]), .B(in1[39]), .ZN(n_0_102));
   XNOR2_X1 i_0_182 (.A(in2[40]), .B(n_0_103), .ZN(sum[40]));
   XNOR2_X1 i_0_183 (.A(in3[40]), .B(in1[63]), .ZN(n_0_103));
   XNOR2_X1 i_0_184 (.A(n_0_105), .B(n_0_104), .ZN(sum[41]));
   XNOR2_X1 i_0_185 (.A(n_0_106), .B(n_0_104), .ZN(sum[42]));
   XNOR2_X1 i_0_186 (.A(n_0_107), .B(n_0_104), .ZN(sum[43]));
   XNOR2_X1 i_0_187 (.A(n_0_108), .B(n_0_104), .ZN(sum[44]));
   XNOR2_X1 i_0_188 (.A(n_0_109), .B(n_0_104), .ZN(sum[45]));
   XNOR2_X1 i_0_189 (.A(n_0_110), .B(n_0_104), .ZN(sum[63]));
   XOR2_X1 i_0_190 (.A(in2[63]), .B(in1[63]), .Z(n_0_104));
   INV_X1 i_0_191 (.A(in3[41]), .ZN(n_0_105));
   INV_X1 i_0_192 (.A(in3[42]), .ZN(n_0_106));
   INV_X1 i_0_193 (.A(in3[43]), .ZN(n_0_107));
   INV_X1 i_0_194 (.A(in3[44]), .ZN(n_0_108));
   INV_X1 i_0_195 (.A(in3[45]), .ZN(n_0_109));
   INV_X1 i_0_196 (.A(in3[63]), .ZN(n_0_110));
endmodule

module CSA__1_35(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;

   AND2_X1 i_0_0 (.A1(in2[24]), .A2(in1[24]), .ZN(c[25]));
   AND2_X1 i_0_1 (.A1(in2[25]), .A2(in1[25]), .ZN(c[26]));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_0), .ZN(c[27]));
   OAI21_X1 i_0_3 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .ZN(c[28]));
   OAI21_X1 i_0_6 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_2));
   NAND2_X1 i_0_7 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_4), .ZN(c[29]));
   OAI21_X1 i_0_9 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_4));
   NAND2_X1 i_0_10 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(n_0_7), .A2(n_0_6), .ZN(c[30]));
   OAI21_X1 i_0_12 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_6));
   NAND2_X1 i_0_13 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_7));
   NAND2_X1 i_0_14 (.A1(n_0_9), .A2(n_0_8), .ZN(c[31]));
   OAI21_X1 i_0_15 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_8));
   NAND2_X1 i_0_16 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_9));
   NAND2_X1 i_0_17 (.A1(n_0_11), .A2(n_0_10), .ZN(c[32]));
   OAI21_X1 i_0_18 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_10));
   NAND2_X1 i_0_19 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_11));
   NAND2_X1 i_0_20 (.A1(n_0_13), .A2(n_0_12), .ZN(c[33]));
   OAI21_X1 i_0_21 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_12));
   NAND2_X1 i_0_22 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_13));
   NAND2_X1 i_0_23 (.A1(n_0_15), .A2(n_0_14), .ZN(c[34]));
   OAI21_X1 i_0_24 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_14));
   NAND2_X1 i_0_25 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_15));
   NAND2_X1 i_0_26 (.A1(n_0_17), .A2(n_0_16), .ZN(c[35]));
   OAI21_X1 i_0_27 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_16));
   NAND2_X1 i_0_28 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_17));
   NAND2_X1 i_0_29 (.A1(n_0_19), .A2(n_0_18), .ZN(c[36]));
   OAI21_X1 i_0_30 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_18));
   NAND2_X1 i_0_31 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_19));
   NAND2_X1 i_0_32 (.A1(n_0_21), .A2(n_0_20), .ZN(c[37]));
   OAI21_X1 i_0_33 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_20));
   NAND2_X1 i_0_34 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_21));
   NAND2_X1 i_0_35 (.A1(n_0_23), .A2(n_0_22), .ZN(c[38]));
   OAI21_X1 i_0_36 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_22));
   NAND2_X1 i_0_37 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_23));
   NAND2_X1 i_0_38 (.A1(n_0_25), .A2(n_0_24), .ZN(c[39]));
   OAI21_X1 i_0_39 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_24));
   NAND2_X1 i_0_40 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_25));
   NAND2_X1 i_0_41 (.A1(n_0_27), .A2(n_0_26), .ZN(c[40]));
   OAI21_X1 i_0_42 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_26));
   NAND2_X1 i_0_43 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_27));
   NAND2_X1 i_0_44 (.A1(n_0_29), .A2(n_0_28), .ZN(c[41]));
   OAI21_X1 i_0_45 (.A(in1[40]), .B1(in3[40]), .B2(in2[40]), .ZN(n_0_28));
   NAND2_X1 i_0_46 (.A1(in2[40]), .A2(in3[40]), .ZN(n_0_29));
   NAND2_X1 i_0_47 (.A1(n_0_31), .A2(n_0_30), .ZN(c[42]));
   OAI21_X1 i_0_48 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_30));
   NAND2_X1 i_0_49 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_31));
   NAND2_X1 i_0_50 (.A1(n_0_33), .A2(n_0_32), .ZN(c[43]));
   OAI21_X1 i_0_51 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_32));
   NAND2_X1 i_0_52 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_33));
   NAND2_X1 i_0_53 (.A1(n_0_35), .A2(n_0_34), .ZN(c[44]));
   OAI21_X1 i_0_54 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_34));
   NAND2_X1 i_0_55 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_35));
   NAND2_X1 i_0_56 (.A1(n_0_37), .A2(n_0_36), .ZN(c[45]));
   OAI21_X1 i_0_57 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_36));
   NAND2_X1 i_0_58 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_37));
   NAND2_X1 i_0_59 (.A1(n_0_39), .A2(n_0_38), .ZN(c[46]));
   OAI21_X1 i_0_60 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_38));
   NAND2_X1 i_0_61 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_39));
   NAND2_X1 i_0_62 (.A1(n_0_41), .A2(n_0_40), .ZN(c[47]));
   OAI21_X1 i_0_63 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_40));
   NAND2_X1 i_0_64 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_41));
   NAND2_X1 i_0_65 (.A1(n_0_43), .A2(n_0_42), .ZN(c[48]));
   OAI21_X1 i_0_66 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_42));
   NAND2_X1 i_0_67 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_43));
   NAND2_X1 i_0_68 (.A1(n_0_45), .A2(n_0_44), .ZN(c[49]));
   OAI21_X1 i_0_69 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_44));
   NAND2_X1 i_0_70 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_45));
   NAND2_X1 i_0_71 (.A1(n_0_47), .A2(n_0_46), .ZN(c[50]));
   OAI21_X1 i_0_72 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_46));
   NAND2_X1 i_0_73 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_47));
   NAND2_X1 i_0_74 (.A1(n_0_49), .A2(n_0_48), .ZN(c[51]));
   OAI21_X1 i_0_75 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_48));
   NAND2_X1 i_0_76 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_49));
   NAND2_X1 i_0_77 (.A1(n_0_51), .A2(n_0_50), .ZN(c[52]));
   OAI21_X1 i_0_78 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_50));
   NAND2_X1 i_0_79 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_51));
   NAND2_X1 i_0_80 (.A1(n_0_53), .A2(n_0_52), .ZN(c[53]));
   OAI21_X1 i_0_81 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_52));
   NAND2_X1 i_0_82 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_53));
   NAND2_X1 i_0_83 (.A1(n_0_55), .A2(n_0_54), .ZN(c[54]));
   OAI21_X1 i_0_84 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_54));
   NAND2_X1 i_0_85 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_55));
   NAND2_X1 i_0_86 (.A1(n_0_57), .A2(n_0_56), .ZN(c[55]));
   OAI21_X1 i_0_87 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_56));
   NAND2_X1 i_0_88 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_57));
   NAND2_X1 i_0_89 (.A1(n_0_59), .A2(n_0_58), .ZN(c[56]));
   OAI21_X1 i_0_90 (.A(in2[55]), .B1(in3[55]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_91 (.A1(in3[55]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_92 (.A1(n_0_61), .A2(n_0_60), .ZN(c[57]));
   OAI21_X1 i_0_93 (.A(in2[56]), .B1(in3[56]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_94 (.A1(in3[56]), .A2(in1[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(n_0_64), .A2(n_0_62), .ZN(c[58]));
   OAI21_X1 i_0_96 (.A(in3[57]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_62));
   NAND2_X1 i_0_97 (.A1(n_0_64), .A2(n_0_63), .ZN(c[63]));
   OAI21_X1 i_0_98 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_63));
   NAND2_X1 i_0_99 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_64));
   XOR2_X1 i_0_100 (.A(in2[24]), .B(in1[24]), .Z(sum[24]));
   XOR2_X1 i_0_101 (.A(in2[25]), .B(in1[25]), .Z(sum[25]));
   XNOR2_X1 i_0_102 (.A(in2[26]), .B(n_0_65), .ZN(sum[26]));
   XNOR2_X1 i_0_103 (.A(in3[26]), .B(in1[26]), .ZN(n_0_65));
   XNOR2_X1 i_0_104 (.A(in2[27]), .B(n_0_66), .ZN(sum[27]));
   XNOR2_X1 i_0_105 (.A(in3[27]), .B(in1[27]), .ZN(n_0_66));
   XNOR2_X1 i_0_106 (.A(in2[28]), .B(n_0_67), .ZN(sum[28]));
   XNOR2_X1 i_0_107 (.A(in3[28]), .B(in1[28]), .ZN(n_0_67));
   XNOR2_X1 i_0_108 (.A(in2[29]), .B(n_0_68), .ZN(sum[29]));
   XNOR2_X1 i_0_109 (.A(in3[29]), .B(in1[29]), .ZN(n_0_68));
   XNOR2_X1 i_0_110 (.A(in2[30]), .B(n_0_69), .ZN(sum[30]));
   XNOR2_X1 i_0_111 (.A(in3[30]), .B(in1[30]), .ZN(n_0_69));
   XNOR2_X1 i_0_112 (.A(in2[31]), .B(n_0_70), .ZN(sum[31]));
   XNOR2_X1 i_0_113 (.A(in3[31]), .B(in1[31]), .ZN(n_0_70));
   XNOR2_X1 i_0_114 (.A(in2[32]), .B(n_0_71), .ZN(sum[32]));
   XNOR2_X1 i_0_115 (.A(in3[32]), .B(in1[32]), .ZN(n_0_71));
   XNOR2_X1 i_0_116 (.A(in2[33]), .B(n_0_72), .ZN(sum[33]));
   XNOR2_X1 i_0_117 (.A(in3[33]), .B(in1[33]), .ZN(n_0_72));
   XNOR2_X1 i_0_118 (.A(in2[34]), .B(n_0_73), .ZN(sum[34]));
   XNOR2_X1 i_0_119 (.A(in3[34]), .B(in1[34]), .ZN(n_0_73));
   XNOR2_X1 i_0_120 (.A(in2[35]), .B(n_0_74), .ZN(sum[35]));
   XNOR2_X1 i_0_121 (.A(in3[35]), .B(in1[35]), .ZN(n_0_74));
   XNOR2_X1 i_0_122 (.A(in2[36]), .B(n_0_75), .ZN(sum[36]));
   XNOR2_X1 i_0_123 (.A(in3[36]), .B(in1[36]), .ZN(n_0_75));
   XNOR2_X1 i_0_124 (.A(in2[37]), .B(n_0_76), .ZN(sum[37]));
   XNOR2_X1 i_0_125 (.A(in3[37]), .B(in1[37]), .ZN(n_0_76));
   XNOR2_X1 i_0_126 (.A(in2[38]), .B(n_0_77), .ZN(sum[38]));
   XNOR2_X1 i_0_127 (.A(in3[38]), .B(in1[38]), .ZN(n_0_77));
   XNOR2_X1 i_0_128 (.A(in2[39]), .B(n_0_78), .ZN(sum[39]));
   XNOR2_X1 i_0_129 (.A(in3[39]), .B(in1[39]), .ZN(n_0_78));
   XNOR2_X1 i_0_130 (.A(in2[40]), .B(n_0_79), .ZN(sum[40]));
   XNOR2_X1 i_0_131 (.A(in3[40]), .B(in1[40]), .ZN(n_0_79));
   XNOR2_X1 i_0_132 (.A(in2[41]), .B(n_0_80), .ZN(sum[41]));
   XNOR2_X1 i_0_133 (.A(in3[41]), .B(in1[41]), .ZN(n_0_80));
   XNOR2_X1 i_0_134 (.A(in2[42]), .B(n_0_81), .ZN(sum[42]));
   XNOR2_X1 i_0_135 (.A(in3[42]), .B(in1[42]), .ZN(n_0_81));
   XNOR2_X1 i_0_136 (.A(in2[43]), .B(n_0_82), .ZN(sum[43]));
   XNOR2_X1 i_0_137 (.A(in3[43]), .B(in1[43]), .ZN(n_0_82));
   XNOR2_X1 i_0_138 (.A(in2[44]), .B(n_0_83), .ZN(sum[44]));
   XNOR2_X1 i_0_139 (.A(in3[44]), .B(in1[44]), .ZN(n_0_83));
   XNOR2_X1 i_0_140 (.A(in2[45]), .B(n_0_84), .ZN(sum[45]));
   XNOR2_X1 i_0_141 (.A(in3[45]), .B(in1[45]), .ZN(n_0_84));
   XNOR2_X1 i_0_142 (.A(in2[46]), .B(n_0_85), .ZN(sum[46]));
   XNOR2_X1 i_0_143 (.A(in3[46]), .B(in1[46]), .ZN(n_0_85));
   XNOR2_X1 i_0_144 (.A(in2[47]), .B(n_0_86), .ZN(sum[47]));
   XNOR2_X1 i_0_145 (.A(in3[47]), .B(in1[47]), .ZN(n_0_86));
   XNOR2_X1 i_0_146 (.A(in2[48]), .B(n_0_87), .ZN(sum[48]));
   XNOR2_X1 i_0_147 (.A(in3[48]), .B(in1[48]), .ZN(n_0_87));
   XNOR2_X1 i_0_148 (.A(in2[49]), .B(n_0_88), .ZN(sum[49]));
   XNOR2_X1 i_0_149 (.A(in3[49]), .B(in1[49]), .ZN(n_0_88));
   XNOR2_X1 i_0_150 (.A(in2[50]), .B(n_0_89), .ZN(sum[50]));
   XNOR2_X1 i_0_151 (.A(in3[50]), .B(in1[50]), .ZN(n_0_89));
   XNOR2_X1 i_0_152 (.A(in2[51]), .B(n_0_90), .ZN(sum[51]));
   XNOR2_X1 i_0_153 (.A(in3[51]), .B(in1[51]), .ZN(n_0_90));
   XNOR2_X1 i_0_154 (.A(in2[52]), .B(n_0_91), .ZN(sum[52]));
   XNOR2_X1 i_0_155 (.A(in3[52]), .B(in1[52]), .ZN(n_0_91));
   XNOR2_X1 i_0_156 (.A(in2[53]), .B(n_0_92), .ZN(sum[53]));
   XNOR2_X1 i_0_157 (.A(in3[53]), .B(in1[53]), .ZN(n_0_92));
   XNOR2_X1 i_0_158 (.A(in2[54]), .B(n_0_93), .ZN(sum[54]));
   XNOR2_X1 i_0_159 (.A(in3[54]), .B(in1[54]), .ZN(n_0_93));
   XNOR2_X1 i_0_160 (.A(in2[55]), .B(n_0_94), .ZN(sum[55]));
   XNOR2_X1 i_0_161 (.A(in3[55]), .B(in1[63]), .ZN(n_0_94));
   XNOR2_X1 i_0_162 (.A(in2[56]), .B(n_0_95), .ZN(sum[56]));
   XNOR2_X1 i_0_163 (.A(in3[56]), .B(in1[63]), .ZN(n_0_95));
   XOR2_X1 i_0_164 (.A(in3[57]), .B(n_0_96), .Z(sum[57]));
   XOR2_X1 i_0_165 (.A(in3[63]), .B(n_0_96), .Z(sum[63]));
   XOR2_X1 i_0_166 (.A(in2[63]), .B(in1[63]), .Z(n_0_96));
endmodule

module CSA__1_38(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;

   AND2_X1 i_0_0 (.A1(in2[23]), .A2(in1[23]), .ZN(c[24]));
   AND2_X1 i_0_1 (.A1(in2[24]), .A2(in1[24]), .ZN(c[25]));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_0), .ZN(c[26]));
   OAI21_X1 i_0_3 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .ZN(c[27]));
   OAI21_X1 i_0_6 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_2));
   NAND2_X1 i_0_7 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_4), .ZN(c[28]));
   OAI21_X1 i_0_9 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_4));
   NAND2_X1 i_0_10 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(n_0_7), .A2(n_0_6), .ZN(c[29]));
   OAI21_X1 i_0_12 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_6));
   NAND2_X1 i_0_13 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_7));
   NAND2_X1 i_0_14 (.A1(n_0_9), .A2(n_0_8), .ZN(c[30]));
   OAI21_X1 i_0_15 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_8));
   NAND2_X1 i_0_16 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_9));
   NAND2_X1 i_0_17 (.A1(n_0_11), .A2(n_0_10), .ZN(c[31]));
   OAI21_X1 i_0_18 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_10));
   NAND2_X1 i_0_19 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_11));
   NAND2_X1 i_0_20 (.A1(n_0_13), .A2(n_0_12), .ZN(c[32]));
   OAI21_X1 i_0_21 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_12));
   NAND2_X1 i_0_22 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_13));
   NAND2_X1 i_0_23 (.A1(n_0_15), .A2(n_0_14), .ZN(c[33]));
   OAI21_X1 i_0_24 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_14));
   NAND2_X1 i_0_25 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_15));
   NAND2_X1 i_0_26 (.A1(n_0_17), .A2(n_0_16), .ZN(c[34]));
   OAI21_X1 i_0_27 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_16));
   NAND2_X1 i_0_28 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_17));
   NAND2_X1 i_0_29 (.A1(n_0_19), .A2(n_0_18), .ZN(c[35]));
   OAI21_X1 i_0_30 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_18));
   NAND2_X1 i_0_31 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_19));
   NAND2_X1 i_0_32 (.A1(n_0_21), .A2(n_0_20), .ZN(c[36]));
   OAI21_X1 i_0_33 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_20));
   NAND2_X1 i_0_34 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_21));
   NAND2_X1 i_0_35 (.A1(n_0_23), .A2(n_0_22), .ZN(c[37]));
   OAI21_X1 i_0_36 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_22));
   NAND2_X1 i_0_37 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_23));
   NAND2_X1 i_0_38 (.A1(n_0_25), .A2(n_0_24), .ZN(c[38]));
   OAI21_X1 i_0_39 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_24));
   NAND2_X1 i_0_40 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_25));
   NAND2_X1 i_0_41 (.A1(n_0_27), .A2(n_0_26), .ZN(c[39]));
   OAI21_X1 i_0_42 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_26));
   NAND2_X1 i_0_43 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_27));
   NAND2_X1 i_0_44 (.A1(n_0_29), .A2(n_0_28), .ZN(c[40]));
   OAI21_X1 i_0_45 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_28));
   NAND2_X1 i_0_46 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_29));
   NAND2_X1 i_0_47 (.A1(n_0_31), .A2(n_0_30), .ZN(c[41]));
   OAI21_X1 i_0_48 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_30));
   NAND2_X1 i_0_49 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_31));
   NAND2_X1 i_0_50 (.A1(n_0_33), .A2(n_0_32), .ZN(c[42]));
   OAI21_X1 i_0_51 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_32));
   NAND2_X1 i_0_52 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_33));
   NAND2_X1 i_0_53 (.A1(n_0_35), .A2(n_0_34), .ZN(c[43]));
   OAI21_X1 i_0_54 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_34));
   NAND2_X1 i_0_55 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_35));
   NAND2_X1 i_0_56 (.A1(n_0_37), .A2(n_0_36), .ZN(c[44]));
   OAI21_X1 i_0_57 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_36));
   NAND2_X1 i_0_58 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_37));
   NAND2_X1 i_0_59 (.A1(n_0_39), .A2(n_0_38), .ZN(c[45]));
   OAI21_X1 i_0_60 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_38));
   NAND2_X1 i_0_61 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_39));
   NAND2_X1 i_0_62 (.A1(n_0_41), .A2(n_0_40), .ZN(c[46]));
   OAI21_X1 i_0_63 (.A(in1[45]), .B1(in3[45]), .B2(in2[45]), .ZN(n_0_40));
   NAND2_X1 i_0_64 (.A1(in2[45]), .A2(in3[45]), .ZN(n_0_41));
   NAND2_X1 i_0_65 (.A1(n_0_43), .A2(n_0_42), .ZN(c[47]));
   OAI21_X1 i_0_66 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_42));
   NAND2_X1 i_0_67 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_43));
   NAND2_X1 i_0_68 (.A1(n_0_45), .A2(n_0_44), .ZN(c[48]));
   OAI21_X1 i_0_69 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_44));
   NAND2_X1 i_0_70 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_45));
   NAND2_X1 i_0_71 (.A1(n_0_47), .A2(n_0_46), .ZN(c[49]));
   OAI21_X1 i_0_72 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_46));
   NAND2_X1 i_0_73 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_47));
   NAND2_X1 i_0_74 (.A1(n_0_49), .A2(n_0_48), .ZN(c[50]));
   OAI21_X1 i_0_75 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_48));
   NAND2_X1 i_0_76 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_49));
   NAND2_X1 i_0_77 (.A1(n_0_51), .A2(n_0_50), .ZN(c[51]));
   OAI21_X1 i_0_78 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_50));
   NAND2_X1 i_0_79 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_51));
   NAND2_X1 i_0_80 (.A1(n_0_53), .A2(n_0_52), .ZN(c[52]));
   OAI21_X1 i_0_81 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_52));
   NAND2_X1 i_0_82 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_53));
   NAND2_X1 i_0_83 (.A1(n_0_55), .A2(n_0_54), .ZN(c[53]));
   OAI21_X1 i_0_84 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_54));
   NAND2_X1 i_0_85 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_55));
   NAND2_X1 i_0_86 (.A1(n_0_57), .A2(n_0_56), .ZN(c[54]));
   OAI21_X1 i_0_87 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_56));
   NAND2_X1 i_0_88 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_57));
   NAND2_X1 i_0_89 (.A1(n_0_59), .A2(n_0_58), .ZN(c[55]));
   OAI21_X1 i_0_90 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_58));
   NAND2_X1 i_0_91 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_59));
   NAND2_X1 i_0_92 (.A1(n_0_61), .A2(n_0_60), .ZN(c[56]));
   OAI21_X1 i_0_93 (.A(in2[55]), .B1(in3[55]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_94 (.A1(in3[55]), .A2(in1[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(n_0_63), .A2(n_0_62), .ZN(c[57]));
   OAI21_X1 i_0_96 (.A(in2[56]), .B1(in3[56]), .B2(in1[63]), .ZN(n_0_62));
   NAND2_X1 i_0_97 (.A1(in3[56]), .A2(in1[63]), .ZN(n_0_63));
   NAND2_X1 i_0_98 (.A1(n_0_65), .A2(n_0_64), .ZN(c[58]));
   OAI21_X1 i_0_99 (.A(in2[57]), .B1(in3[57]), .B2(in1[63]), .ZN(n_0_64));
   NAND2_X1 i_0_100 (.A1(in3[57]), .A2(in1[63]), .ZN(n_0_65));
   NAND2_X1 i_0_101 (.A1(n_0_68), .A2(n_0_66), .ZN(c[59]));
   OAI21_X1 i_0_102 (.A(in3[58]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_66));
   NAND2_X1 i_0_103 (.A1(n_0_68), .A2(n_0_67), .ZN(c[63]));
   OAI21_X1 i_0_104 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_67));
   NAND2_X1 i_0_105 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_68));
   XOR2_X1 i_0_106 (.A(in2[23]), .B(in1[23]), .Z(sum[23]));
   XOR2_X1 i_0_107 (.A(in2[24]), .B(in1[24]), .Z(sum[24]));
   XNOR2_X1 i_0_108 (.A(in2[25]), .B(n_0_69), .ZN(sum[25]));
   XNOR2_X1 i_0_109 (.A(in3[25]), .B(in1[25]), .ZN(n_0_69));
   XNOR2_X1 i_0_110 (.A(in2[26]), .B(n_0_70), .ZN(sum[26]));
   XNOR2_X1 i_0_111 (.A(in3[26]), .B(in1[26]), .ZN(n_0_70));
   XNOR2_X1 i_0_112 (.A(in2[27]), .B(n_0_71), .ZN(sum[27]));
   XNOR2_X1 i_0_113 (.A(in3[27]), .B(in1[27]), .ZN(n_0_71));
   XNOR2_X1 i_0_114 (.A(in2[28]), .B(n_0_72), .ZN(sum[28]));
   XNOR2_X1 i_0_115 (.A(in3[28]), .B(in1[28]), .ZN(n_0_72));
   XNOR2_X1 i_0_116 (.A(in2[29]), .B(n_0_73), .ZN(sum[29]));
   XNOR2_X1 i_0_117 (.A(in3[29]), .B(in1[29]), .ZN(n_0_73));
   XNOR2_X1 i_0_118 (.A(in2[30]), .B(n_0_74), .ZN(sum[30]));
   XNOR2_X1 i_0_119 (.A(in3[30]), .B(in1[30]), .ZN(n_0_74));
   XNOR2_X1 i_0_120 (.A(in2[31]), .B(n_0_75), .ZN(sum[31]));
   XNOR2_X1 i_0_121 (.A(in3[31]), .B(in1[31]), .ZN(n_0_75));
   XNOR2_X1 i_0_122 (.A(in2[32]), .B(n_0_76), .ZN(sum[32]));
   XNOR2_X1 i_0_123 (.A(in3[32]), .B(in1[32]), .ZN(n_0_76));
   XNOR2_X1 i_0_124 (.A(in2[33]), .B(n_0_77), .ZN(sum[33]));
   XNOR2_X1 i_0_125 (.A(in3[33]), .B(in1[33]), .ZN(n_0_77));
   XNOR2_X1 i_0_126 (.A(in2[34]), .B(n_0_78), .ZN(sum[34]));
   XNOR2_X1 i_0_127 (.A(in3[34]), .B(in1[34]), .ZN(n_0_78));
   XNOR2_X1 i_0_128 (.A(in2[35]), .B(n_0_79), .ZN(sum[35]));
   XNOR2_X1 i_0_129 (.A(in3[35]), .B(in1[35]), .ZN(n_0_79));
   XNOR2_X1 i_0_130 (.A(in2[36]), .B(n_0_80), .ZN(sum[36]));
   XNOR2_X1 i_0_131 (.A(in3[36]), .B(in1[36]), .ZN(n_0_80));
   XNOR2_X1 i_0_132 (.A(in2[37]), .B(n_0_81), .ZN(sum[37]));
   XNOR2_X1 i_0_133 (.A(in3[37]), .B(in1[37]), .ZN(n_0_81));
   XNOR2_X1 i_0_134 (.A(in2[38]), .B(n_0_82), .ZN(sum[38]));
   XNOR2_X1 i_0_135 (.A(in3[38]), .B(in1[38]), .ZN(n_0_82));
   XNOR2_X1 i_0_136 (.A(in2[39]), .B(n_0_83), .ZN(sum[39]));
   XNOR2_X1 i_0_137 (.A(in3[39]), .B(in1[39]), .ZN(n_0_83));
   XNOR2_X1 i_0_138 (.A(in2[40]), .B(n_0_84), .ZN(sum[40]));
   XNOR2_X1 i_0_139 (.A(in3[40]), .B(in1[40]), .ZN(n_0_84));
   XNOR2_X1 i_0_140 (.A(in2[41]), .B(n_0_85), .ZN(sum[41]));
   XNOR2_X1 i_0_141 (.A(in3[41]), .B(in1[41]), .ZN(n_0_85));
   XNOR2_X1 i_0_142 (.A(in2[42]), .B(n_0_86), .ZN(sum[42]));
   XNOR2_X1 i_0_143 (.A(in3[42]), .B(in1[42]), .ZN(n_0_86));
   XNOR2_X1 i_0_144 (.A(in2[43]), .B(n_0_87), .ZN(sum[43]));
   XNOR2_X1 i_0_145 (.A(in3[43]), .B(in1[43]), .ZN(n_0_87));
   XNOR2_X1 i_0_146 (.A(in2[44]), .B(n_0_88), .ZN(sum[44]));
   XNOR2_X1 i_0_147 (.A(in3[44]), .B(in1[44]), .ZN(n_0_88));
   XNOR2_X1 i_0_148 (.A(in2[45]), .B(n_0_89), .ZN(sum[45]));
   XNOR2_X1 i_0_149 (.A(in3[45]), .B(in1[45]), .ZN(n_0_89));
   XNOR2_X1 i_0_150 (.A(in2[46]), .B(n_0_90), .ZN(sum[46]));
   XNOR2_X1 i_0_151 (.A(in3[46]), .B(in1[46]), .ZN(n_0_90));
   XNOR2_X1 i_0_152 (.A(in2[47]), .B(n_0_91), .ZN(sum[47]));
   XNOR2_X1 i_0_153 (.A(in3[47]), .B(in1[47]), .ZN(n_0_91));
   XNOR2_X1 i_0_154 (.A(in2[48]), .B(n_0_92), .ZN(sum[48]));
   XNOR2_X1 i_0_155 (.A(in3[48]), .B(in1[48]), .ZN(n_0_92));
   XNOR2_X1 i_0_156 (.A(in2[49]), .B(n_0_93), .ZN(sum[49]));
   XNOR2_X1 i_0_157 (.A(in3[49]), .B(in1[49]), .ZN(n_0_93));
   XNOR2_X1 i_0_158 (.A(in2[50]), .B(n_0_94), .ZN(sum[50]));
   XNOR2_X1 i_0_159 (.A(in3[50]), .B(in1[50]), .ZN(n_0_94));
   XNOR2_X1 i_0_160 (.A(in2[51]), .B(n_0_95), .ZN(sum[51]));
   XNOR2_X1 i_0_161 (.A(in3[51]), .B(in1[51]), .ZN(n_0_95));
   XNOR2_X1 i_0_162 (.A(in2[52]), .B(n_0_96), .ZN(sum[52]));
   XNOR2_X1 i_0_163 (.A(in3[52]), .B(in1[52]), .ZN(n_0_96));
   XNOR2_X1 i_0_164 (.A(in2[53]), .B(n_0_97), .ZN(sum[53]));
   XNOR2_X1 i_0_165 (.A(in3[53]), .B(in1[53]), .ZN(n_0_97));
   XNOR2_X1 i_0_166 (.A(in2[54]), .B(n_0_98), .ZN(sum[54]));
   XNOR2_X1 i_0_167 (.A(in3[54]), .B(in1[54]), .ZN(n_0_98));
   XNOR2_X1 i_0_168 (.A(in2[55]), .B(n_0_99), .ZN(sum[55]));
   XNOR2_X1 i_0_169 (.A(in3[55]), .B(in1[63]), .ZN(n_0_99));
   XNOR2_X1 i_0_170 (.A(in2[56]), .B(n_0_100), .ZN(sum[56]));
   XNOR2_X1 i_0_171 (.A(in3[56]), .B(in1[63]), .ZN(n_0_100));
   XNOR2_X1 i_0_172 (.A(in2[57]), .B(n_0_101), .ZN(sum[57]));
   XNOR2_X1 i_0_173 (.A(in3[57]), .B(in1[63]), .ZN(n_0_101));
   XOR2_X1 i_0_174 (.A(in3[58]), .B(n_0_102), .Z(sum[58]));
   XOR2_X1 i_0_175 (.A(in3[63]), .B(n_0_102), .Z(sum[63]));
   XOR2_X1 i_0_176 (.A(in2[63]), .B(in1[63]), .Z(n_0_102));
endmodule

module CSA__0_68(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;

   AND2_X1 i_0_0 (.A1(in2[22]), .A2(in1[22]), .ZN(c[23]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[24]));
   OAI21_X1 i_0_2 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[25]));
   OAI21_X1 i_0_5 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[26]));
   OAI21_X1 i_0_8 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[27]));
   OAI21_X1 i_0_11 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[28]));
   OAI21_X1 i_0_14 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[29]));
   OAI21_X1 i_0_17 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[30]));
   OAI21_X1 i_0_20 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[31]));
   OAI21_X1 i_0_23 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[32]));
   OAI21_X1 i_0_26 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[33]));
   OAI21_X1 i_0_29 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[34]));
   OAI21_X1 i_0_32 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[35]));
   OAI21_X1 i_0_35 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[36]));
   OAI21_X1 i_0_38 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[37]));
   OAI21_X1 i_0_41 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[38]));
   OAI21_X1 i_0_44 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[39]));
   OAI21_X1 i_0_47 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[40]));
   OAI21_X1 i_0_50 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[41]));
   OAI21_X1 i_0_53 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[42]));
   OAI21_X1 i_0_56 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[43]));
   OAI21_X1 i_0_59 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[44]));
   OAI21_X1 i_0_62 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[45]));
   OAI21_X1 i_0_65 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[46]));
   OAI21_X1 i_0_68 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[47]));
   OAI21_X1 i_0_71 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[48]));
   OAI21_X1 i_0_74 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[49]));
   OAI21_X1 i_0_77 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[50]));
   OAI21_X1 i_0_80 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[51]));
   OAI21_X1 i_0_83 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[52]));
   OAI21_X1 i_0_86 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[53]));
   OAI21_X1 i_0_89 (.A(in2[52]), .B1(in3[52]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[52]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_62), .A2(n_0_60), .ZN(c[54]));
   OAI21_X1 i_0_92 (.A(in3[53]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(c[63]));
   OAI21_X1 i_0_94 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   XOR2_X1 i_0_96 (.A(in2[22]), .B(in1[22]), .Z(sum[22]));
   XNOR2_X1 i_0_97 (.A(in2[23]), .B(n_0_63), .ZN(sum[23]));
   XNOR2_X1 i_0_98 (.A(in3[23]), .B(in1[23]), .ZN(n_0_63));
   XNOR2_X1 i_0_99 (.A(in2[24]), .B(n_0_64), .ZN(sum[24]));
   XNOR2_X1 i_0_100 (.A(in3[24]), .B(in1[24]), .ZN(n_0_64));
   XNOR2_X1 i_0_101 (.A(in2[25]), .B(n_0_65), .ZN(sum[25]));
   XNOR2_X1 i_0_102 (.A(in3[25]), .B(in1[25]), .ZN(n_0_65));
   XNOR2_X1 i_0_103 (.A(in2[26]), .B(n_0_66), .ZN(sum[26]));
   XNOR2_X1 i_0_104 (.A(in3[26]), .B(in1[26]), .ZN(n_0_66));
   XNOR2_X1 i_0_105 (.A(in2[27]), .B(n_0_67), .ZN(sum[27]));
   XNOR2_X1 i_0_106 (.A(in3[27]), .B(in1[27]), .ZN(n_0_67));
   XNOR2_X1 i_0_107 (.A(in2[28]), .B(n_0_68), .ZN(sum[28]));
   XNOR2_X1 i_0_108 (.A(in3[28]), .B(in1[28]), .ZN(n_0_68));
   XNOR2_X1 i_0_109 (.A(in2[29]), .B(n_0_69), .ZN(sum[29]));
   XNOR2_X1 i_0_110 (.A(in3[29]), .B(in1[29]), .ZN(n_0_69));
   XNOR2_X1 i_0_111 (.A(in2[30]), .B(n_0_70), .ZN(sum[30]));
   XNOR2_X1 i_0_112 (.A(in3[30]), .B(in1[30]), .ZN(n_0_70));
   XNOR2_X1 i_0_113 (.A(in2[31]), .B(n_0_71), .ZN(sum[31]));
   XNOR2_X1 i_0_114 (.A(in3[31]), .B(in1[31]), .ZN(n_0_71));
   XNOR2_X1 i_0_115 (.A(in2[32]), .B(n_0_72), .ZN(sum[32]));
   XNOR2_X1 i_0_116 (.A(in3[32]), .B(in1[32]), .ZN(n_0_72));
   XNOR2_X1 i_0_117 (.A(in2[33]), .B(n_0_73), .ZN(sum[33]));
   XNOR2_X1 i_0_118 (.A(in3[33]), .B(in1[33]), .ZN(n_0_73));
   XNOR2_X1 i_0_119 (.A(in2[34]), .B(n_0_74), .ZN(sum[34]));
   XNOR2_X1 i_0_120 (.A(in3[34]), .B(in1[34]), .ZN(n_0_74));
   XNOR2_X1 i_0_121 (.A(in2[35]), .B(n_0_75), .ZN(sum[35]));
   XNOR2_X1 i_0_122 (.A(in3[35]), .B(in1[35]), .ZN(n_0_75));
   XNOR2_X1 i_0_123 (.A(in2[36]), .B(n_0_76), .ZN(sum[36]));
   XNOR2_X1 i_0_124 (.A(in3[36]), .B(in1[36]), .ZN(n_0_76));
   XNOR2_X1 i_0_125 (.A(in2[37]), .B(n_0_77), .ZN(sum[37]));
   XNOR2_X1 i_0_126 (.A(in3[37]), .B(in1[37]), .ZN(n_0_77));
   XNOR2_X1 i_0_127 (.A(in2[38]), .B(n_0_78), .ZN(sum[38]));
   XNOR2_X1 i_0_128 (.A(in3[38]), .B(in1[38]), .ZN(n_0_78));
   XNOR2_X1 i_0_129 (.A(in2[39]), .B(n_0_79), .ZN(sum[39]));
   XNOR2_X1 i_0_130 (.A(in3[39]), .B(in1[39]), .ZN(n_0_79));
   XNOR2_X1 i_0_131 (.A(in2[40]), .B(n_0_80), .ZN(sum[40]));
   XNOR2_X1 i_0_132 (.A(in3[40]), .B(in1[40]), .ZN(n_0_80));
   XNOR2_X1 i_0_133 (.A(in2[41]), .B(n_0_81), .ZN(sum[41]));
   XNOR2_X1 i_0_134 (.A(in3[41]), .B(in1[41]), .ZN(n_0_81));
   XNOR2_X1 i_0_135 (.A(in2[42]), .B(n_0_82), .ZN(sum[42]));
   XNOR2_X1 i_0_136 (.A(in3[42]), .B(in1[42]), .ZN(n_0_82));
   XNOR2_X1 i_0_137 (.A(in2[43]), .B(n_0_83), .ZN(sum[43]));
   XNOR2_X1 i_0_138 (.A(in3[43]), .B(in1[43]), .ZN(n_0_83));
   XNOR2_X1 i_0_139 (.A(in2[44]), .B(n_0_84), .ZN(sum[44]));
   XNOR2_X1 i_0_140 (.A(in3[44]), .B(in1[44]), .ZN(n_0_84));
   XNOR2_X1 i_0_141 (.A(in2[45]), .B(n_0_85), .ZN(sum[45]));
   XNOR2_X1 i_0_142 (.A(in3[45]), .B(in1[45]), .ZN(n_0_85));
   XNOR2_X1 i_0_143 (.A(in2[46]), .B(n_0_86), .ZN(sum[46]));
   XNOR2_X1 i_0_144 (.A(in3[46]), .B(in1[46]), .ZN(n_0_86));
   XNOR2_X1 i_0_145 (.A(in2[47]), .B(n_0_87), .ZN(sum[47]));
   XNOR2_X1 i_0_146 (.A(in3[47]), .B(in1[47]), .ZN(n_0_87));
   XNOR2_X1 i_0_147 (.A(in2[48]), .B(n_0_88), .ZN(sum[48]));
   XNOR2_X1 i_0_148 (.A(in3[48]), .B(in1[48]), .ZN(n_0_88));
   XNOR2_X1 i_0_149 (.A(in2[49]), .B(n_0_89), .ZN(sum[49]));
   XNOR2_X1 i_0_150 (.A(in3[49]), .B(in1[49]), .ZN(n_0_89));
   XNOR2_X1 i_0_151 (.A(in2[50]), .B(n_0_90), .ZN(sum[50]));
   XNOR2_X1 i_0_152 (.A(in3[50]), .B(in1[50]), .ZN(n_0_90));
   XNOR2_X1 i_0_153 (.A(in2[51]), .B(n_0_91), .ZN(sum[51]));
   XNOR2_X1 i_0_154 (.A(in3[51]), .B(in1[51]), .ZN(n_0_91));
   XNOR2_X1 i_0_155 (.A(in2[52]), .B(n_0_92), .ZN(sum[52]));
   XNOR2_X1 i_0_156 (.A(in3[52]), .B(in1[63]), .ZN(n_0_92));
   XOR2_X1 i_0_157 (.A(in3[53]), .B(n_0_93), .Z(sum[53]));
   XOR2_X1 i_0_158 (.A(in3[63]), .B(n_0_93), .Z(sum[63]));
   XOR2_X1 i_0_159 (.A(in2[63]), .B(in1[63]), .Z(n_0_93));
endmodule

module CSA__2_2(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;

   AND2_X1 i_0_0 (.A1(in2[15]), .A2(in1[15]), .ZN(c[16]));
   AND2_X1 i_0_1 (.A1(in2[16]), .A2(in1[16]), .ZN(c[17]));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_0), .ZN(c[18]));
   OAI21_X1 i_0_3 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .ZN(c[19]));
   OAI21_X1 i_0_6 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_2));
   NAND2_X1 i_0_7 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_4), .ZN(c[20]));
   OAI21_X1 i_0_9 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_4));
   NAND2_X1 i_0_10 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(n_0_7), .A2(n_0_6), .ZN(c[21]));
   OAI21_X1 i_0_12 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_6));
   NAND2_X1 i_0_13 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_7));
   NAND2_X1 i_0_14 (.A1(n_0_9), .A2(n_0_8), .ZN(c[22]));
   OAI21_X1 i_0_15 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_8));
   NAND2_X1 i_0_16 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_9));
   NAND2_X1 i_0_17 (.A1(n_0_11), .A2(n_0_10), .ZN(c[23]));
   OAI21_X1 i_0_18 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_10));
   NAND2_X1 i_0_19 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_11));
   NAND2_X1 i_0_20 (.A1(n_0_13), .A2(n_0_12), .ZN(c[24]));
   OAI21_X1 i_0_21 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_12));
   NAND2_X1 i_0_22 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_13));
   NAND2_X1 i_0_23 (.A1(n_0_15), .A2(n_0_14), .ZN(c[25]));
   OAI21_X1 i_0_24 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_14));
   NAND2_X1 i_0_25 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_15));
   NAND2_X1 i_0_26 (.A1(n_0_17), .A2(n_0_16), .ZN(c[26]));
   OAI21_X1 i_0_27 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_16));
   NAND2_X1 i_0_28 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_17));
   NAND2_X1 i_0_29 (.A1(n_0_19), .A2(n_0_18), .ZN(c[27]));
   OAI21_X1 i_0_30 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_18));
   NAND2_X1 i_0_31 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_19));
   NAND2_X1 i_0_32 (.A1(n_0_21), .A2(n_0_20), .ZN(c[28]));
   OAI21_X1 i_0_33 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_20));
   NAND2_X1 i_0_34 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_21));
   NAND2_X1 i_0_35 (.A1(n_0_23), .A2(n_0_22), .ZN(c[29]));
   OAI21_X1 i_0_36 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_22));
   NAND2_X1 i_0_37 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_23));
   NAND2_X1 i_0_38 (.A1(n_0_25), .A2(n_0_24), .ZN(c[30]));
   OAI21_X1 i_0_39 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_24));
   NAND2_X1 i_0_40 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_25));
   NAND2_X1 i_0_41 (.A1(n_0_27), .A2(n_0_26), .ZN(c[31]));
   OAI21_X1 i_0_42 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_26));
   NAND2_X1 i_0_43 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_27));
   NAND2_X1 i_0_44 (.A1(n_0_29), .A2(n_0_28), .ZN(c[32]));
   OAI21_X1 i_0_45 (.A(in1[31]), .B1(in3[31]), .B2(in2[31]), .ZN(n_0_28));
   NAND2_X1 i_0_46 (.A1(in2[31]), .A2(in3[31]), .ZN(n_0_29));
   NAND2_X1 i_0_47 (.A1(n_0_31), .A2(n_0_30), .ZN(c[33]));
   OAI21_X1 i_0_48 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_30));
   NAND2_X1 i_0_49 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_31));
   NAND2_X1 i_0_50 (.A1(n_0_33), .A2(n_0_32), .ZN(c[34]));
   OAI21_X1 i_0_51 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_32));
   NAND2_X1 i_0_52 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_33));
   NAND2_X1 i_0_53 (.A1(n_0_35), .A2(n_0_34), .ZN(c[35]));
   OAI21_X1 i_0_54 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_34));
   NAND2_X1 i_0_55 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_35));
   NAND2_X1 i_0_56 (.A1(n_0_37), .A2(n_0_36), .ZN(c[36]));
   OAI21_X1 i_0_57 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_36));
   NAND2_X1 i_0_58 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_37));
   NAND2_X1 i_0_59 (.A1(n_0_39), .A2(n_0_38), .ZN(c[37]));
   OAI21_X1 i_0_60 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_38));
   NAND2_X1 i_0_61 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_39));
   NAND2_X1 i_0_62 (.A1(n_0_41), .A2(n_0_40), .ZN(c[38]));
   OAI21_X1 i_0_63 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_40));
   NAND2_X1 i_0_64 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_41));
   NAND2_X1 i_0_65 (.A1(n_0_43), .A2(n_0_42), .ZN(c[39]));
   OAI21_X1 i_0_66 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_42));
   NAND2_X1 i_0_67 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_43));
   NAND2_X1 i_0_68 (.A1(n_0_45), .A2(n_0_44), .ZN(c[40]));
   OAI21_X1 i_0_69 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_44));
   NAND2_X1 i_0_70 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_45));
   NAND2_X1 i_0_71 (.A1(n_0_47), .A2(n_0_46), .ZN(c[41]));
   OAI21_X1 i_0_72 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_46));
   NAND2_X1 i_0_73 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_47));
   NAND2_X1 i_0_74 (.A1(n_0_49), .A2(n_0_48), .ZN(c[42]));
   OAI21_X1 i_0_75 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_48));
   NAND2_X1 i_0_76 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_49));
   NAND2_X1 i_0_77 (.A1(n_0_51), .A2(n_0_50), .ZN(c[43]));
   OAI21_X1 i_0_78 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_50));
   NAND2_X1 i_0_79 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_51));
   NAND2_X1 i_0_80 (.A1(n_0_53), .A2(n_0_52), .ZN(c[44]));
   OAI21_X1 i_0_81 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_52));
   NAND2_X1 i_0_82 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_53));
   NAND2_X1 i_0_83 (.A1(n_0_55), .A2(n_0_54), .ZN(c[45]));
   OAI21_X1 i_0_84 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_54));
   NAND2_X1 i_0_85 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_55));
   NAND2_X1 i_0_86 (.A1(n_0_57), .A2(n_0_56), .ZN(c[46]));
   OAI21_X1 i_0_87 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_56));
   NAND2_X1 i_0_88 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_57));
   NAND2_X1 i_0_89 (.A1(n_0_59), .A2(n_0_58), .ZN(c[47]));
   OAI21_X1 i_0_90 (.A(in2[46]), .B1(in3[46]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_91 (.A1(in3[46]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_92 (.A1(n_0_61), .A2(n_0_60), .ZN(c[48]));
   OAI21_X1 i_0_93 (.A(in2[47]), .B1(in3[47]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_94 (.A1(in3[47]), .A2(in1[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(n_0_64), .A2(n_0_62), .ZN(c[49]));
   OAI21_X1 i_0_96 (.A(in3[48]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_62));
   NAND2_X1 i_0_97 (.A1(n_0_64), .A2(n_0_63), .ZN(c[63]));
   OAI21_X1 i_0_98 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_63));
   NAND2_X1 i_0_99 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_64));
   XOR2_X1 i_0_100 (.A(in2[15]), .B(in1[15]), .Z(sum[15]));
   XOR2_X1 i_0_101 (.A(in2[16]), .B(in1[16]), .Z(sum[16]));
   XNOR2_X1 i_0_102 (.A(in2[17]), .B(n_0_65), .ZN(sum[17]));
   XNOR2_X1 i_0_103 (.A(in3[17]), .B(in1[17]), .ZN(n_0_65));
   XNOR2_X1 i_0_104 (.A(in2[18]), .B(n_0_66), .ZN(sum[18]));
   XNOR2_X1 i_0_105 (.A(in3[18]), .B(in1[18]), .ZN(n_0_66));
   XNOR2_X1 i_0_106 (.A(in2[19]), .B(n_0_67), .ZN(sum[19]));
   XNOR2_X1 i_0_107 (.A(in3[19]), .B(in1[19]), .ZN(n_0_67));
   XNOR2_X1 i_0_108 (.A(in2[20]), .B(n_0_68), .ZN(sum[20]));
   XNOR2_X1 i_0_109 (.A(in3[20]), .B(in1[20]), .ZN(n_0_68));
   XNOR2_X1 i_0_110 (.A(in2[21]), .B(n_0_69), .ZN(sum[21]));
   XNOR2_X1 i_0_111 (.A(in3[21]), .B(in1[21]), .ZN(n_0_69));
   XNOR2_X1 i_0_112 (.A(in2[22]), .B(n_0_70), .ZN(sum[22]));
   XNOR2_X1 i_0_113 (.A(in3[22]), .B(in1[22]), .ZN(n_0_70));
   XNOR2_X1 i_0_114 (.A(in2[23]), .B(n_0_71), .ZN(sum[23]));
   XNOR2_X1 i_0_115 (.A(in3[23]), .B(in1[23]), .ZN(n_0_71));
   XNOR2_X1 i_0_116 (.A(in2[24]), .B(n_0_72), .ZN(sum[24]));
   XNOR2_X1 i_0_117 (.A(in3[24]), .B(in1[24]), .ZN(n_0_72));
   XNOR2_X1 i_0_118 (.A(in2[25]), .B(n_0_73), .ZN(sum[25]));
   XNOR2_X1 i_0_119 (.A(in3[25]), .B(in1[25]), .ZN(n_0_73));
   XNOR2_X1 i_0_120 (.A(in2[26]), .B(n_0_74), .ZN(sum[26]));
   XNOR2_X1 i_0_121 (.A(in3[26]), .B(in1[26]), .ZN(n_0_74));
   XNOR2_X1 i_0_122 (.A(in2[27]), .B(n_0_75), .ZN(sum[27]));
   XNOR2_X1 i_0_123 (.A(in3[27]), .B(in1[27]), .ZN(n_0_75));
   XNOR2_X1 i_0_124 (.A(in2[28]), .B(n_0_76), .ZN(sum[28]));
   XNOR2_X1 i_0_125 (.A(in3[28]), .B(in1[28]), .ZN(n_0_76));
   XNOR2_X1 i_0_126 (.A(in2[29]), .B(n_0_77), .ZN(sum[29]));
   XNOR2_X1 i_0_127 (.A(in3[29]), .B(in1[29]), .ZN(n_0_77));
   XNOR2_X1 i_0_128 (.A(in2[30]), .B(n_0_78), .ZN(sum[30]));
   XNOR2_X1 i_0_129 (.A(in3[30]), .B(in1[30]), .ZN(n_0_78));
   XNOR2_X1 i_0_130 (.A(in2[31]), .B(n_0_79), .ZN(sum[31]));
   XNOR2_X1 i_0_131 (.A(in3[31]), .B(in1[31]), .ZN(n_0_79));
   XNOR2_X1 i_0_132 (.A(in2[32]), .B(n_0_80), .ZN(sum[32]));
   XNOR2_X1 i_0_133 (.A(in3[32]), .B(in1[32]), .ZN(n_0_80));
   XNOR2_X1 i_0_134 (.A(in2[33]), .B(n_0_81), .ZN(sum[33]));
   XNOR2_X1 i_0_135 (.A(in3[33]), .B(in1[33]), .ZN(n_0_81));
   XNOR2_X1 i_0_136 (.A(in2[34]), .B(n_0_82), .ZN(sum[34]));
   XNOR2_X1 i_0_137 (.A(in3[34]), .B(in1[34]), .ZN(n_0_82));
   XNOR2_X1 i_0_138 (.A(in2[35]), .B(n_0_83), .ZN(sum[35]));
   XNOR2_X1 i_0_139 (.A(in3[35]), .B(in1[35]), .ZN(n_0_83));
   XNOR2_X1 i_0_140 (.A(in2[36]), .B(n_0_84), .ZN(sum[36]));
   XNOR2_X1 i_0_141 (.A(in3[36]), .B(in1[36]), .ZN(n_0_84));
   XNOR2_X1 i_0_142 (.A(in2[37]), .B(n_0_85), .ZN(sum[37]));
   XNOR2_X1 i_0_143 (.A(in3[37]), .B(in1[37]), .ZN(n_0_85));
   XNOR2_X1 i_0_144 (.A(in2[38]), .B(n_0_86), .ZN(sum[38]));
   XNOR2_X1 i_0_145 (.A(in3[38]), .B(in1[38]), .ZN(n_0_86));
   XNOR2_X1 i_0_146 (.A(in2[39]), .B(n_0_87), .ZN(sum[39]));
   XNOR2_X1 i_0_147 (.A(in3[39]), .B(in1[39]), .ZN(n_0_87));
   XNOR2_X1 i_0_148 (.A(in2[40]), .B(n_0_88), .ZN(sum[40]));
   XNOR2_X1 i_0_149 (.A(in3[40]), .B(in1[40]), .ZN(n_0_88));
   XNOR2_X1 i_0_150 (.A(in2[41]), .B(n_0_89), .ZN(sum[41]));
   XNOR2_X1 i_0_151 (.A(in3[41]), .B(in1[41]), .ZN(n_0_89));
   XNOR2_X1 i_0_152 (.A(in2[42]), .B(n_0_90), .ZN(sum[42]));
   XNOR2_X1 i_0_153 (.A(in3[42]), .B(in1[42]), .ZN(n_0_90));
   XNOR2_X1 i_0_154 (.A(in2[43]), .B(n_0_91), .ZN(sum[43]));
   XNOR2_X1 i_0_155 (.A(in3[43]), .B(in1[43]), .ZN(n_0_91));
   XNOR2_X1 i_0_156 (.A(in2[44]), .B(n_0_92), .ZN(sum[44]));
   XNOR2_X1 i_0_157 (.A(in3[44]), .B(in1[44]), .ZN(n_0_92));
   XNOR2_X1 i_0_158 (.A(in2[45]), .B(n_0_93), .ZN(sum[45]));
   XNOR2_X1 i_0_159 (.A(in3[45]), .B(in1[45]), .ZN(n_0_93));
   XNOR2_X1 i_0_160 (.A(in2[46]), .B(n_0_94), .ZN(sum[46]));
   XNOR2_X1 i_0_161 (.A(in3[46]), .B(in1[63]), .ZN(n_0_94));
   XNOR2_X1 i_0_162 (.A(in2[47]), .B(n_0_95), .ZN(sum[47]));
   XNOR2_X1 i_0_163 (.A(in3[47]), .B(in1[63]), .ZN(n_0_95));
   XOR2_X1 i_0_164 (.A(in3[48]), .B(n_0_96), .Z(sum[48]));
   XOR2_X1 i_0_165 (.A(in3[63]), .B(n_0_96), .Z(sum[63]));
   XOR2_X1 i_0_166 (.A(in2[63]), .B(in1[63]), .Z(n_0_96));
endmodule

module CSA__2_5(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;

   AND2_X1 i_0_0 (.A1(in2[16]), .A2(in1[16]), .ZN(c[17]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[18]));
   OAI21_X1 i_0_2 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[19]));
   OAI21_X1 i_0_5 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[20]));
   OAI21_X1 i_0_8 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[21]));
   OAI21_X1 i_0_11 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[22]));
   OAI21_X1 i_0_14 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[23]));
   OAI21_X1 i_0_17 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[24]));
   OAI21_X1 i_0_20 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[25]));
   OAI21_X1 i_0_23 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[26]));
   OAI21_X1 i_0_26 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[27]));
   OAI21_X1 i_0_29 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[28]));
   OAI21_X1 i_0_32 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[29]));
   OAI21_X1 i_0_35 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[30]));
   OAI21_X1 i_0_38 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[31]));
   OAI21_X1 i_0_41 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[32]));
   OAI21_X1 i_0_44 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[33]));
   OAI21_X1 i_0_47 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[34]));
   OAI21_X1 i_0_50 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[35]));
   OAI21_X1 i_0_53 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[36]));
   OAI21_X1 i_0_56 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[37]));
   OAI21_X1 i_0_59 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[38]));
   OAI21_X1 i_0_62 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[39]));
   OAI21_X1 i_0_65 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[40]));
   OAI21_X1 i_0_68 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[41]));
   OAI21_X1 i_0_71 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[42]));
   OAI21_X1 i_0_74 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[43]));
   OAI21_X1 i_0_77 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[44]));
   OAI21_X1 i_0_80 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[45]));
   OAI21_X1 i_0_83 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[46]));
   OAI21_X1 i_0_86 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[47]));
   OAI21_X1 i_0_89 (.A(in2[46]), .B1(in3[46]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[46]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_62), .A2(n_0_60), .ZN(c[48]));
   OAI21_X1 i_0_92 (.A(in3[47]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(c[63]));
   OAI21_X1 i_0_94 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   XOR2_X1 i_0_96 (.A(in2[16]), .B(in1[16]), .Z(sum[16]));
   XNOR2_X1 i_0_97 (.A(in2[17]), .B(n_0_63), .ZN(sum[17]));
   XNOR2_X1 i_0_98 (.A(in3[17]), .B(in1[17]), .ZN(n_0_63));
   XNOR2_X1 i_0_99 (.A(in2[18]), .B(n_0_64), .ZN(sum[18]));
   XNOR2_X1 i_0_100 (.A(in3[18]), .B(in1[18]), .ZN(n_0_64));
   XNOR2_X1 i_0_101 (.A(in2[19]), .B(n_0_65), .ZN(sum[19]));
   XNOR2_X1 i_0_102 (.A(in3[19]), .B(in1[19]), .ZN(n_0_65));
   XNOR2_X1 i_0_103 (.A(in2[20]), .B(n_0_66), .ZN(sum[20]));
   XNOR2_X1 i_0_104 (.A(in3[20]), .B(in1[20]), .ZN(n_0_66));
   XNOR2_X1 i_0_105 (.A(in2[21]), .B(n_0_67), .ZN(sum[21]));
   XNOR2_X1 i_0_106 (.A(in3[21]), .B(in1[21]), .ZN(n_0_67));
   XNOR2_X1 i_0_107 (.A(in2[22]), .B(n_0_68), .ZN(sum[22]));
   XNOR2_X1 i_0_108 (.A(in3[22]), .B(in1[22]), .ZN(n_0_68));
   XNOR2_X1 i_0_109 (.A(in2[23]), .B(n_0_69), .ZN(sum[23]));
   XNOR2_X1 i_0_110 (.A(in3[23]), .B(in1[23]), .ZN(n_0_69));
   XNOR2_X1 i_0_111 (.A(in2[24]), .B(n_0_70), .ZN(sum[24]));
   XNOR2_X1 i_0_112 (.A(in3[24]), .B(in1[24]), .ZN(n_0_70));
   XNOR2_X1 i_0_113 (.A(in2[25]), .B(n_0_71), .ZN(sum[25]));
   XNOR2_X1 i_0_114 (.A(in3[25]), .B(in1[25]), .ZN(n_0_71));
   XNOR2_X1 i_0_115 (.A(in2[26]), .B(n_0_72), .ZN(sum[26]));
   XNOR2_X1 i_0_116 (.A(in3[26]), .B(in1[26]), .ZN(n_0_72));
   XNOR2_X1 i_0_117 (.A(in2[27]), .B(n_0_73), .ZN(sum[27]));
   XNOR2_X1 i_0_118 (.A(in3[27]), .B(in1[27]), .ZN(n_0_73));
   XNOR2_X1 i_0_119 (.A(in2[28]), .B(n_0_74), .ZN(sum[28]));
   XNOR2_X1 i_0_120 (.A(in3[28]), .B(in1[28]), .ZN(n_0_74));
   XNOR2_X1 i_0_121 (.A(in2[29]), .B(n_0_75), .ZN(sum[29]));
   XNOR2_X1 i_0_122 (.A(in3[29]), .B(in1[29]), .ZN(n_0_75));
   XNOR2_X1 i_0_123 (.A(in2[30]), .B(n_0_76), .ZN(sum[30]));
   XNOR2_X1 i_0_124 (.A(in3[30]), .B(in1[30]), .ZN(n_0_76));
   XNOR2_X1 i_0_125 (.A(in2[31]), .B(n_0_77), .ZN(sum[31]));
   XNOR2_X1 i_0_126 (.A(in3[31]), .B(in1[31]), .ZN(n_0_77));
   XNOR2_X1 i_0_127 (.A(in2[32]), .B(n_0_78), .ZN(sum[32]));
   XNOR2_X1 i_0_128 (.A(in3[32]), .B(in1[32]), .ZN(n_0_78));
   XNOR2_X1 i_0_129 (.A(in2[33]), .B(n_0_79), .ZN(sum[33]));
   XNOR2_X1 i_0_130 (.A(in3[33]), .B(in1[33]), .ZN(n_0_79));
   XNOR2_X1 i_0_131 (.A(in2[34]), .B(n_0_80), .ZN(sum[34]));
   XNOR2_X1 i_0_132 (.A(in3[34]), .B(in1[34]), .ZN(n_0_80));
   XNOR2_X1 i_0_133 (.A(in2[35]), .B(n_0_81), .ZN(sum[35]));
   XNOR2_X1 i_0_134 (.A(in3[35]), .B(in1[35]), .ZN(n_0_81));
   XNOR2_X1 i_0_135 (.A(in2[36]), .B(n_0_82), .ZN(sum[36]));
   XNOR2_X1 i_0_136 (.A(in3[36]), .B(in1[36]), .ZN(n_0_82));
   XNOR2_X1 i_0_137 (.A(in2[37]), .B(n_0_83), .ZN(sum[37]));
   XNOR2_X1 i_0_138 (.A(in3[37]), .B(in1[37]), .ZN(n_0_83));
   XNOR2_X1 i_0_139 (.A(in2[38]), .B(n_0_84), .ZN(sum[38]));
   XNOR2_X1 i_0_140 (.A(in3[38]), .B(in1[38]), .ZN(n_0_84));
   XNOR2_X1 i_0_141 (.A(in2[39]), .B(n_0_85), .ZN(sum[39]));
   XNOR2_X1 i_0_142 (.A(in3[39]), .B(in1[39]), .ZN(n_0_85));
   XNOR2_X1 i_0_143 (.A(in2[40]), .B(n_0_86), .ZN(sum[40]));
   XNOR2_X1 i_0_144 (.A(in3[40]), .B(in1[40]), .ZN(n_0_86));
   XNOR2_X1 i_0_145 (.A(in2[41]), .B(n_0_87), .ZN(sum[41]));
   XNOR2_X1 i_0_146 (.A(in3[41]), .B(in1[41]), .ZN(n_0_87));
   XNOR2_X1 i_0_147 (.A(in2[42]), .B(n_0_88), .ZN(sum[42]));
   XNOR2_X1 i_0_148 (.A(in3[42]), .B(in1[42]), .ZN(n_0_88));
   XNOR2_X1 i_0_149 (.A(in2[43]), .B(n_0_89), .ZN(sum[43]));
   XNOR2_X1 i_0_150 (.A(in3[43]), .B(in1[43]), .ZN(n_0_89));
   XNOR2_X1 i_0_151 (.A(in2[44]), .B(n_0_90), .ZN(sum[44]));
   XNOR2_X1 i_0_152 (.A(in3[44]), .B(in1[44]), .ZN(n_0_90));
   XNOR2_X1 i_0_153 (.A(in2[45]), .B(n_0_91), .ZN(sum[45]));
   XNOR2_X1 i_0_154 (.A(in3[45]), .B(in1[45]), .ZN(n_0_91));
   XNOR2_X1 i_0_155 (.A(in2[46]), .B(n_0_92), .ZN(sum[46]));
   XNOR2_X1 i_0_156 (.A(in3[46]), .B(in1[63]), .ZN(n_0_92));
   XOR2_X1 i_0_157 (.A(in3[47]), .B(n_0_93), .Z(sum[47]));
   XOR2_X1 i_0_158 (.A(in3[63]), .B(n_0_93), .Z(sum[63]));
   XOR2_X1 i_0_159 (.A(in2[63]), .B(in1[63]), .Z(n_0_93));
endmodule

module CSA__0_71(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;

   AND2_X1 i_0_0 (.A1(in2[13]), .A2(in1[13]), .ZN(c[14]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[15]));
   OAI21_X1 i_0_2 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[16]));
   OAI21_X1 i_0_5 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[17]));
   OAI21_X1 i_0_8 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[18]));
   OAI21_X1 i_0_11 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[19]));
   OAI21_X1 i_0_14 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[20]));
   OAI21_X1 i_0_17 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[21]));
   OAI21_X1 i_0_20 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[22]));
   OAI21_X1 i_0_23 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[23]));
   OAI21_X1 i_0_26 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[24]));
   OAI21_X1 i_0_29 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[25]));
   OAI21_X1 i_0_32 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[26]));
   OAI21_X1 i_0_35 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[27]));
   OAI21_X1 i_0_38 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[28]));
   OAI21_X1 i_0_41 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[29]));
   OAI21_X1 i_0_44 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[30]));
   OAI21_X1 i_0_47 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[31]));
   OAI21_X1 i_0_50 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[32]));
   OAI21_X1 i_0_53 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[33]));
   OAI21_X1 i_0_56 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[34]));
   OAI21_X1 i_0_59 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[35]));
   OAI21_X1 i_0_62 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[36]));
   OAI21_X1 i_0_65 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[37]));
   OAI21_X1 i_0_68 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[38]));
   OAI21_X1 i_0_71 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[39]));
   OAI21_X1 i_0_74 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[40]));
   OAI21_X1 i_0_77 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[41]));
   OAI21_X1 i_0_80 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[42]));
   OAI21_X1 i_0_83 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[43]));
   OAI21_X1 i_0_86 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[44]));
   OAI21_X1 i_0_89 (.A(in2[43]), .B1(in3[43]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[43]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_62), .A2(n_0_60), .ZN(c[45]));
   OAI21_X1 i_0_92 (.A(in3[44]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(c[63]));
   OAI21_X1 i_0_94 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   XOR2_X1 i_0_96 (.A(in2[13]), .B(in1[13]), .Z(sum[13]));
   XNOR2_X1 i_0_97 (.A(in2[14]), .B(n_0_63), .ZN(sum[14]));
   XNOR2_X1 i_0_98 (.A(in3[14]), .B(in1[14]), .ZN(n_0_63));
   XNOR2_X1 i_0_99 (.A(in2[15]), .B(n_0_64), .ZN(sum[15]));
   XNOR2_X1 i_0_100 (.A(in3[15]), .B(in1[15]), .ZN(n_0_64));
   XNOR2_X1 i_0_101 (.A(in2[16]), .B(n_0_65), .ZN(sum[16]));
   XNOR2_X1 i_0_102 (.A(in3[16]), .B(in1[16]), .ZN(n_0_65));
   XNOR2_X1 i_0_103 (.A(in2[17]), .B(n_0_66), .ZN(sum[17]));
   XNOR2_X1 i_0_104 (.A(in3[17]), .B(in1[17]), .ZN(n_0_66));
   XNOR2_X1 i_0_105 (.A(in2[18]), .B(n_0_67), .ZN(sum[18]));
   XNOR2_X1 i_0_106 (.A(in3[18]), .B(in1[18]), .ZN(n_0_67));
   XNOR2_X1 i_0_107 (.A(in2[19]), .B(n_0_68), .ZN(sum[19]));
   XNOR2_X1 i_0_108 (.A(in3[19]), .B(in1[19]), .ZN(n_0_68));
   XNOR2_X1 i_0_109 (.A(in2[20]), .B(n_0_69), .ZN(sum[20]));
   XNOR2_X1 i_0_110 (.A(in3[20]), .B(in1[20]), .ZN(n_0_69));
   XNOR2_X1 i_0_111 (.A(in2[21]), .B(n_0_70), .ZN(sum[21]));
   XNOR2_X1 i_0_112 (.A(in3[21]), .B(in1[21]), .ZN(n_0_70));
   XNOR2_X1 i_0_113 (.A(in2[22]), .B(n_0_71), .ZN(sum[22]));
   XNOR2_X1 i_0_114 (.A(in3[22]), .B(in1[22]), .ZN(n_0_71));
   XNOR2_X1 i_0_115 (.A(in2[23]), .B(n_0_72), .ZN(sum[23]));
   XNOR2_X1 i_0_116 (.A(in3[23]), .B(in1[23]), .ZN(n_0_72));
   XNOR2_X1 i_0_117 (.A(in2[24]), .B(n_0_73), .ZN(sum[24]));
   XNOR2_X1 i_0_118 (.A(in3[24]), .B(in1[24]), .ZN(n_0_73));
   XNOR2_X1 i_0_119 (.A(in2[25]), .B(n_0_74), .ZN(sum[25]));
   XNOR2_X1 i_0_120 (.A(in3[25]), .B(in1[25]), .ZN(n_0_74));
   XNOR2_X1 i_0_121 (.A(in2[26]), .B(n_0_75), .ZN(sum[26]));
   XNOR2_X1 i_0_122 (.A(in3[26]), .B(in1[26]), .ZN(n_0_75));
   XNOR2_X1 i_0_123 (.A(in2[27]), .B(n_0_76), .ZN(sum[27]));
   XNOR2_X1 i_0_124 (.A(in3[27]), .B(in1[27]), .ZN(n_0_76));
   XNOR2_X1 i_0_125 (.A(in2[28]), .B(n_0_77), .ZN(sum[28]));
   XNOR2_X1 i_0_126 (.A(in3[28]), .B(in1[28]), .ZN(n_0_77));
   XNOR2_X1 i_0_127 (.A(in2[29]), .B(n_0_78), .ZN(sum[29]));
   XNOR2_X1 i_0_128 (.A(in3[29]), .B(in1[29]), .ZN(n_0_78));
   XNOR2_X1 i_0_129 (.A(in2[30]), .B(n_0_79), .ZN(sum[30]));
   XNOR2_X1 i_0_130 (.A(in3[30]), .B(in1[30]), .ZN(n_0_79));
   XNOR2_X1 i_0_131 (.A(in2[31]), .B(n_0_80), .ZN(sum[31]));
   XNOR2_X1 i_0_132 (.A(in3[31]), .B(in1[31]), .ZN(n_0_80));
   XNOR2_X1 i_0_133 (.A(in2[32]), .B(n_0_81), .ZN(sum[32]));
   XNOR2_X1 i_0_134 (.A(in3[32]), .B(in1[32]), .ZN(n_0_81));
   XNOR2_X1 i_0_135 (.A(in2[33]), .B(n_0_82), .ZN(sum[33]));
   XNOR2_X1 i_0_136 (.A(in3[33]), .B(in1[33]), .ZN(n_0_82));
   XNOR2_X1 i_0_137 (.A(in2[34]), .B(n_0_83), .ZN(sum[34]));
   XNOR2_X1 i_0_138 (.A(in3[34]), .B(in1[34]), .ZN(n_0_83));
   XNOR2_X1 i_0_139 (.A(in2[35]), .B(n_0_84), .ZN(sum[35]));
   XNOR2_X1 i_0_140 (.A(in3[35]), .B(in1[35]), .ZN(n_0_84));
   XNOR2_X1 i_0_141 (.A(in2[36]), .B(n_0_85), .ZN(sum[36]));
   XNOR2_X1 i_0_142 (.A(in3[36]), .B(in1[36]), .ZN(n_0_85));
   XNOR2_X1 i_0_143 (.A(in2[37]), .B(n_0_86), .ZN(sum[37]));
   XNOR2_X1 i_0_144 (.A(in3[37]), .B(in1[37]), .ZN(n_0_86));
   XNOR2_X1 i_0_145 (.A(in2[38]), .B(n_0_87), .ZN(sum[38]));
   XNOR2_X1 i_0_146 (.A(in3[38]), .B(in1[38]), .ZN(n_0_87));
   XNOR2_X1 i_0_147 (.A(in2[39]), .B(n_0_88), .ZN(sum[39]));
   XNOR2_X1 i_0_148 (.A(in3[39]), .B(in1[39]), .ZN(n_0_88));
   XNOR2_X1 i_0_149 (.A(in2[40]), .B(n_0_89), .ZN(sum[40]));
   XNOR2_X1 i_0_150 (.A(in3[40]), .B(in1[40]), .ZN(n_0_89));
   XNOR2_X1 i_0_151 (.A(in2[41]), .B(n_0_90), .ZN(sum[41]));
   XNOR2_X1 i_0_152 (.A(in3[41]), .B(in1[41]), .ZN(n_0_90));
   XNOR2_X1 i_0_153 (.A(in2[42]), .B(n_0_91), .ZN(sum[42]));
   XNOR2_X1 i_0_154 (.A(in3[42]), .B(in1[42]), .ZN(n_0_91));
   XNOR2_X1 i_0_155 (.A(in2[43]), .B(n_0_92), .ZN(sum[43]));
   XNOR2_X1 i_0_156 (.A(in3[43]), .B(in1[63]), .ZN(n_0_92));
   XOR2_X1 i_0_157 (.A(in3[44]), .B(n_0_93), .Z(sum[44]));
   XOR2_X1 i_0_158 (.A(in3[63]), .B(n_0_93), .Z(sum[63]));
   XOR2_X1 i_0_159 (.A(in2[63]), .B(in1[63]), .Z(n_0_93));
endmodule

module CSA__3_2(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_116;
   wire n_0_115;
   wire n_0_114;
   wire n_0_113;
   wire n_0_122;
   wire n_0_112;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;

   AND2_X1 i_0_0 (.A1(in2[5]), .A2(in1[5]), .ZN(c[6]));
   AND2_X1 i_0_1 (.A1(in2[6]), .A2(in1[6]), .ZN(c[7]));
   AND2_X1 i_0_2 (.A1(in2[7]), .A2(in1[7]), .ZN(c[8]));
   AND2_X1 i_0_3 (.A1(in2[8]), .A2(in1[8]), .ZN(c[9]));
   AND2_X1 i_0_4 (.A1(in2[9]), .A2(in1[9]), .ZN(c[10]));
   NAND2_X1 i_0_5 (.A1(n_0_1), .A2(n_0_0), .ZN(c[11]));
   OAI21_X1 i_0_6 (.A(in2[10]), .B1(in3[10]), .B2(in1[10]), .ZN(n_0_0));
   NAND2_X1 i_0_7 (.A1(in3[10]), .A2(in1[10]), .ZN(n_0_1));
   NAND2_X1 i_0_8 (.A1(n_0_3), .A2(n_0_2), .ZN(c[12]));
   OAI21_X1 i_0_9 (.A(in2[11]), .B1(in3[11]), .B2(in1[11]), .ZN(n_0_2));
   NAND2_X1 i_0_10 (.A1(in3[11]), .A2(in1[11]), .ZN(n_0_3));
   NAND2_X1 i_0_11 (.A1(n_0_5), .A2(n_0_4), .ZN(c[13]));
   OAI21_X1 i_0_12 (.A(in2[12]), .B1(in3[12]), .B2(in1[12]), .ZN(n_0_4));
   NAND2_X1 i_0_13 (.A1(in3[12]), .A2(in1[12]), .ZN(n_0_5));
   NAND2_X1 i_0_14 (.A1(n_0_7), .A2(n_0_6), .ZN(c[14]));
   OAI21_X1 i_0_15 (.A(in2[13]), .B1(in3[13]), .B2(in1[13]), .ZN(n_0_6));
   NAND2_X1 i_0_16 (.A1(in3[13]), .A2(in1[13]), .ZN(n_0_7));
   NAND2_X1 i_0_17 (.A1(n_0_9), .A2(n_0_8), .ZN(c[15]));
   OAI21_X1 i_0_18 (.A(in2[14]), .B1(in3[14]), .B2(in1[14]), .ZN(n_0_8));
   NAND2_X1 i_0_19 (.A1(in3[14]), .A2(in1[14]), .ZN(n_0_9));
   NAND2_X1 i_0_20 (.A1(n_0_11), .A2(n_0_10), .ZN(c[16]));
   OAI21_X1 i_0_21 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_10));
   NAND2_X1 i_0_22 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_11));
   NAND2_X1 i_0_23 (.A1(n_0_13), .A2(n_0_12), .ZN(c[17]));
   OAI21_X1 i_0_24 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_12));
   NAND2_X1 i_0_25 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_13));
   NAND2_X1 i_0_26 (.A1(n_0_15), .A2(n_0_14), .ZN(c[18]));
   OAI21_X1 i_0_27 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_14));
   NAND2_X1 i_0_28 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_15));
   NAND2_X1 i_0_29 (.A1(n_0_17), .A2(n_0_16), .ZN(c[19]));
   OAI21_X1 i_0_30 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_16));
   NAND2_X1 i_0_31 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_17));
   NAND2_X1 i_0_32 (.A1(n_0_19), .A2(n_0_18), .ZN(c[20]));
   OAI21_X1 i_0_33 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_18));
   NAND2_X1 i_0_34 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_19));
   NAND2_X1 i_0_35 (.A1(n_0_21), .A2(n_0_20), .ZN(c[21]));
   OAI21_X1 i_0_36 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_20));
   NAND2_X1 i_0_37 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_21));
   NAND2_X1 i_0_38 (.A1(n_0_23), .A2(n_0_22), .ZN(c[22]));
   OAI21_X1 i_0_39 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_22));
   NAND2_X1 i_0_40 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_23));
   NAND2_X1 i_0_41 (.A1(n_0_25), .A2(n_0_24), .ZN(c[23]));
   OAI21_X1 i_0_42 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_24));
   NAND2_X1 i_0_43 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_25));
   NAND2_X1 i_0_44 (.A1(n_0_27), .A2(n_0_26), .ZN(c[24]));
   OAI21_X1 i_0_45 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_26));
   NAND2_X1 i_0_46 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_27));
   NAND2_X1 i_0_47 (.A1(n_0_29), .A2(n_0_28), .ZN(c[25]));
   OAI21_X1 i_0_48 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_28));
   NAND2_X1 i_0_49 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_29));
   NAND2_X1 i_0_50 (.A1(n_0_31), .A2(n_0_30), .ZN(c[26]));
   OAI21_X1 i_0_51 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_30));
   NAND2_X1 i_0_52 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_31));
   NAND2_X1 i_0_53 (.A1(n_0_33), .A2(n_0_32), .ZN(c[27]));
   OAI21_X1 i_0_54 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_32));
   NAND2_X1 i_0_55 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_33));
   NAND2_X1 i_0_56 (.A1(n_0_35), .A2(n_0_34), .ZN(c[28]));
   OAI21_X1 i_0_57 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_34));
   NAND2_X1 i_0_58 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_35));
   NAND2_X1 i_0_59 (.A1(n_0_37), .A2(n_0_36), .ZN(c[29]));
   OAI21_X1 i_0_60 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_36));
   NAND2_X1 i_0_61 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_37));
   NAND2_X1 i_0_62 (.A1(n_0_39), .A2(n_0_38), .ZN(c[30]));
   OAI21_X1 i_0_63 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_38));
   NAND2_X1 i_0_64 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_39));
   NAND2_X1 i_0_65 (.A1(n_0_41), .A2(n_0_40), .ZN(c[31]));
   OAI21_X1 i_0_66 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_40));
   NAND2_X1 i_0_67 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_41));
   NAND2_X1 i_0_68 (.A1(n_0_43), .A2(n_0_42), .ZN(c[32]));
   OAI21_X1 i_0_69 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_42));
   NAND2_X1 i_0_70 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_43));
   NAND2_X1 i_0_71 (.A1(n_0_45), .A2(n_0_44), .ZN(c[33]));
   OAI21_X1 i_0_72 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_44));
   NAND2_X1 i_0_73 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_45));
   NAND2_X1 i_0_74 (.A1(n_0_47), .A2(n_0_46), .ZN(c[34]));
   OAI21_X1 i_0_75 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_46));
   NAND2_X1 i_0_76 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_47));
   NAND2_X1 i_0_77 (.A1(n_0_49), .A2(n_0_48), .ZN(c[35]));
   OAI21_X1 i_0_78 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_48));
   NAND2_X1 i_0_79 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_49));
   NAND2_X1 i_0_80 (.A1(n_0_51), .A2(n_0_50), .ZN(c[36]));
   OAI21_X1 i_0_81 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_50));
   NAND2_X1 i_0_82 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_51));
   NAND2_X1 i_0_83 (.A1(n_0_53), .A2(n_0_52), .ZN(c[37]));
   OAI21_X1 i_0_84 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_52));
   NAND2_X1 i_0_85 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_53));
   NAND2_X1 i_0_86 (.A1(n_0_55), .A2(n_0_54), .ZN(c[38]));
   OAI21_X1 i_0_87 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_54));
   NAND2_X1 i_0_88 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_55));
   NAND2_X1 i_0_89 (.A1(n_0_57), .A2(n_0_56), .ZN(c[39]));
   OAI21_X1 i_0_90 (.A(in1[38]), .B1(in3[38]), .B2(in2[38]), .ZN(n_0_56));
   NAND2_X1 i_0_91 (.A1(in2[38]), .A2(in3[38]), .ZN(n_0_57));
   NAND2_X1 i_0_92 (.A1(n_0_59), .A2(n_0_58), .ZN(c[40]));
   OAI21_X1 i_0_93 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_58));
   NAND2_X1 i_0_94 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_59));
   NAND2_X1 i_0_95 (.A1(n_0_61), .A2(n_0_60), .ZN(c[41]));
   OAI21_X1 i_0_96 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_60));
   NAND2_X1 i_0_97 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_61));
   NAND2_X1 i_0_98 (.A1(n_0_63), .A2(n_0_62), .ZN(c[42]));
   OAI21_X1 i_0_99 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_62));
   NAND2_X1 i_0_100 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_63));
   NAND2_X1 i_0_101 (.A1(n_0_65), .A2(n_0_64), .ZN(c[43]));
   OAI21_X1 i_0_102 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_64));
   NAND2_X1 i_0_103 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_65));
   NAND2_X1 i_0_104 (.A1(n_0_67), .A2(n_0_66), .ZN(c[44]));
   OAI21_X1 i_0_105 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_66));
   NAND2_X1 i_0_106 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_67));
   NAND2_X1 i_0_107 (.A1(n_0_69), .A2(n_0_68), .ZN(c[45]));
   OAI21_X1 i_0_108 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_68));
   NAND2_X1 i_0_109 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_69));
   NAND2_X1 i_0_110 (.A1(n_0_71), .A2(n_0_70), .ZN(c[46]));
   OAI21_X1 i_0_111 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_70));
   NAND2_X1 i_0_112 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_71));
   NAND2_X1 i_0_113 (.A1(n_0_73), .A2(n_0_72), .ZN(c[47]));
   OAI21_X1 i_0_114 (.A(in2[46]), .B1(in3[46]), .B2(in1[63]), .ZN(n_0_72));
   NAND2_X1 i_0_115 (.A1(in3[46]), .A2(in1[63]), .ZN(n_0_73));
   AOI21_X1 i_0_116 (.A(n_0_75), .B1(n_0_74), .B2(n_0_114), .ZN(c[48]));
   AOI21_X1 i_0_117 (.A(n_0_75), .B1(n_0_74), .B2(n_0_115), .ZN(c[49]));
   AOI21_X1 i_0_118 (.A(n_0_75), .B1(n_0_74), .B2(n_0_116), .ZN(c[50]));
   AOI21_X1 i_0_119 (.A(n_0_75), .B1(n_0_74), .B2(n_0_117), .ZN(c[51]));
   AOI21_X1 i_0_120 (.A(n_0_75), .B1(n_0_74), .B2(n_0_118), .ZN(c[52]));
   AOI21_X1 i_0_121 (.A(n_0_75), .B1(n_0_74), .B2(n_0_119), .ZN(c[53]));
   AOI21_X1 i_0_122 (.A(n_0_75), .B1(n_0_74), .B2(n_0_120), .ZN(c[54]));
   AOI21_X1 i_0_123 (.A(n_0_75), .B1(n_0_74), .B2(n_0_121), .ZN(c[55]));
   AOI21_X1 i_0_124 (.A(n_0_75), .B1(n_0_74), .B2(n_0_122), .ZN(c[63]));
   NAND2_X1 i_0_125 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_74));
   NOR2_X1 i_0_126 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_75));
   XOR2_X1 i_0_127 (.A(in2[5]), .B(in1[5]), .Z(sum[5]));
   XOR2_X1 i_0_128 (.A(in2[6]), .B(in1[6]), .Z(sum[6]));
   XOR2_X1 i_0_129 (.A(in2[7]), .B(in1[7]), .Z(sum[7]));
   XOR2_X1 i_0_130 (.A(in2[8]), .B(in1[8]), .Z(sum[8]));
   XOR2_X1 i_0_131 (.A(in2[9]), .B(in1[9]), .Z(sum[9]));
   XNOR2_X1 i_0_132 (.A(in2[10]), .B(n_0_76), .ZN(sum[10]));
   XNOR2_X1 i_0_133 (.A(in3[10]), .B(in1[10]), .ZN(n_0_76));
   XNOR2_X1 i_0_134 (.A(in2[11]), .B(n_0_77), .ZN(sum[11]));
   XNOR2_X1 i_0_135 (.A(in3[11]), .B(in1[11]), .ZN(n_0_77));
   XNOR2_X1 i_0_136 (.A(in2[12]), .B(n_0_78), .ZN(sum[12]));
   XNOR2_X1 i_0_137 (.A(in3[12]), .B(in1[12]), .ZN(n_0_78));
   XNOR2_X1 i_0_138 (.A(in2[13]), .B(n_0_79), .ZN(sum[13]));
   XNOR2_X1 i_0_139 (.A(in3[13]), .B(in1[13]), .ZN(n_0_79));
   XNOR2_X1 i_0_140 (.A(in2[14]), .B(n_0_80), .ZN(sum[14]));
   XNOR2_X1 i_0_141 (.A(in3[14]), .B(in1[14]), .ZN(n_0_80));
   XNOR2_X1 i_0_142 (.A(in2[15]), .B(n_0_81), .ZN(sum[15]));
   XNOR2_X1 i_0_143 (.A(in3[15]), .B(in1[15]), .ZN(n_0_81));
   XNOR2_X1 i_0_144 (.A(in2[16]), .B(n_0_82), .ZN(sum[16]));
   XNOR2_X1 i_0_145 (.A(in3[16]), .B(in1[16]), .ZN(n_0_82));
   XNOR2_X1 i_0_146 (.A(in2[17]), .B(n_0_83), .ZN(sum[17]));
   XNOR2_X1 i_0_147 (.A(in3[17]), .B(in1[17]), .ZN(n_0_83));
   XNOR2_X1 i_0_148 (.A(in2[18]), .B(n_0_84), .ZN(sum[18]));
   XNOR2_X1 i_0_149 (.A(in3[18]), .B(in1[18]), .ZN(n_0_84));
   XNOR2_X1 i_0_150 (.A(in2[19]), .B(n_0_85), .ZN(sum[19]));
   XNOR2_X1 i_0_151 (.A(in3[19]), .B(in1[19]), .ZN(n_0_85));
   XNOR2_X1 i_0_152 (.A(in2[20]), .B(n_0_86), .ZN(sum[20]));
   XNOR2_X1 i_0_153 (.A(in3[20]), .B(in1[20]), .ZN(n_0_86));
   XNOR2_X1 i_0_154 (.A(in2[21]), .B(n_0_87), .ZN(sum[21]));
   XNOR2_X1 i_0_155 (.A(in3[21]), .B(in1[21]), .ZN(n_0_87));
   XNOR2_X1 i_0_156 (.A(in2[22]), .B(n_0_88), .ZN(sum[22]));
   XNOR2_X1 i_0_157 (.A(in3[22]), .B(in1[22]), .ZN(n_0_88));
   XNOR2_X1 i_0_158 (.A(in2[23]), .B(n_0_89), .ZN(sum[23]));
   XNOR2_X1 i_0_159 (.A(in3[23]), .B(in1[23]), .ZN(n_0_89));
   XNOR2_X1 i_0_160 (.A(in2[24]), .B(n_0_90), .ZN(sum[24]));
   XNOR2_X1 i_0_161 (.A(in3[24]), .B(in1[24]), .ZN(n_0_90));
   XNOR2_X1 i_0_162 (.A(in2[25]), .B(n_0_91), .ZN(sum[25]));
   XNOR2_X1 i_0_163 (.A(in3[25]), .B(in1[25]), .ZN(n_0_91));
   XNOR2_X1 i_0_164 (.A(in2[26]), .B(n_0_92), .ZN(sum[26]));
   XNOR2_X1 i_0_165 (.A(in3[26]), .B(in1[26]), .ZN(n_0_92));
   XNOR2_X1 i_0_166 (.A(in2[27]), .B(n_0_93), .ZN(sum[27]));
   XNOR2_X1 i_0_167 (.A(in3[27]), .B(in1[27]), .ZN(n_0_93));
   XNOR2_X1 i_0_168 (.A(in2[28]), .B(n_0_94), .ZN(sum[28]));
   XNOR2_X1 i_0_169 (.A(in3[28]), .B(in1[28]), .ZN(n_0_94));
   XNOR2_X1 i_0_170 (.A(in2[29]), .B(n_0_95), .ZN(sum[29]));
   XNOR2_X1 i_0_171 (.A(in3[29]), .B(in1[29]), .ZN(n_0_95));
   XNOR2_X1 i_0_172 (.A(in2[30]), .B(n_0_96), .ZN(sum[30]));
   XNOR2_X1 i_0_173 (.A(in3[30]), .B(in1[30]), .ZN(n_0_96));
   XNOR2_X1 i_0_174 (.A(in2[31]), .B(n_0_97), .ZN(sum[31]));
   XNOR2_X1 i_0_175 (.A(in3[31]), .B(in1[31]), .ZN(n_0_97));
   XNOR2_X1 i_0_176 (.A(in2[32]), .B(n_0_98), .ZN(sum[32]));
   XNOR2_X1 i_0_177 (.A(in3[32]), .B(in1[32]), .ZN(n_0_98));
   XNOR2_X1 i_0_178 (.A(in2[33]), .B(n_0_99), .ZN(sum[33]));
   XNOR2_X1 i_0_179 (.A(in3[33]), .B(in1[33]), .ZN(n_0_99));
   XNOR2_X1 i_0_180 (.A(in2[34]), .B(n_0_100), .ZN(sum[34]));
   XNOR2_X1 i_0_181 (.A(in3[34]), .B(in1[34]), .ZN(n_0_100));
   XNOR2_X1 i_0_182 (.A(in2[35]), .B(n_0_101), .ZN(sum[35]));
   XNOR2_X1 i_0_183 (.A(in3[35]), .B(in1[35]), .ZN(n_0_101));
   XNOR2_X1 i_0_184 (.A(in2[36]), .B(n_0_102), .ZN(sum[36]));
   XNOR2_X1 i_0_185 (.A(in3[36]), .B(in1[36]), .ZN(n_0_102));
   XNOR2_X1 i_0_186 (.A(in2[37]), .B(n_0_103), .ZN(sum[37]));
   XNOR2_X1 i_0_187 (.A(in3[37]), .B(in1[37]), .ZN(n_0_103));
   XNOR2_X1 i_0_188 (.A(in2[38]), .B(n_0_104), .ZN(sum[38]));
   XNOR2_X1 i_0_189 (.A(in3[38]), .B(in1[38]), .ZN(n_0_104));
   XNOR2_X1 i_0_190 (.A(in2[39]), .B(n_0_105), .ZN(sum[39]));
   XNOR2_X1 i_0_191 (.A(in3[39]), .B(in1[39]), .ZN(n_0_105));
   XNOR2_X1 i_0_192 (.A(in2[40]), .B(n_0_106), .ZN(sum[40]));
   XNOR2_X1 i_0_193 (.A(in3[40]), .B(in1[40]), .ZN(n_0_106));
   XNOR2_X1 i_0_194 (.A(in2[41]), .B(n_0_107), .ZN(sum[41]));
   XNOR2_X1 i_0_195 (.A(in3[41]), .B(in1[41]), .ZN(n_0_107));
   XNOR2_X1 i_0_196 (.A(in2[42]), .B(n_0_108), .ZN(sum[42]));
   XNOR2_X1 i_0_197 (.A(in3[42]), .B(in1[42]), .ZN(n_0_108));
   XNOR2_X1 i_0_198 (.A(in2[43]), .B(n_0_109), .ZN(sum[43]));
   XNOR2_X1 i_0_199 (.A(in3[43]), .B(in1[43]), .ZN(n_0_109));
   XNOR2_X1 i_0_200 (.A(in2[44]), .B(n_0_110), .ZN(sum[44]));
   XNOR2_X1 i_0_201 (.A(in3[44]), .B(in1[44]), .ZN(n_0_110));
   XNOR2_X1 i_0_202 (.A(in2[45]), .B(n_0_111), .ZN(sum[45]));
   XNOR2_X1 i_0_203 (.A(in3[45]), .B(in1[45]), .ZN(n_0_111));
   XNOR2_X1 i_0_209 (.A(n_0_117), .B(n_0_113), .ZN(sum[50]));
   XNOR2_X1 i_0_210 (.A(n_0_118), .B(n_0_113), .ZN(sum[51]));
   XNOR2_X1 i_0_211 (.A(n_0_119), .B(n_0_113), .ZN(sum[52]));
   XNOR2_X1 i_0_212 (.A(n_0_120), .B(n_0_113), .ZN(sum[53]));
   XNOR2_X1 i_0_213 (.A(n_0_121), .B(n_0_113), .ZN(sum[54]));
   INV_X1 i_0_219 (.A(in3[50]), .ZN(n_0_117));
   INV_X1 i_0_220 (.A(in3[51]), .ZN(n_0_118));
   INV_X1 i_0_221 (.A(in3[52]), .ZN(n_0_119));
   INV_X1 i_0_222 (.A(in3[53]), .ZN(n_0_120));
   INV_X1 i_0_223 (.A(in3[54]), .ZN(n_0_121));
   INV_X1 i_0_204 (.A(in3[49]), .ZN(n_0_116));
   INV_X1 i_0_205 (.A(in3[48]), .ZN(n_0_115));
   INV_X1 i_0_206 (.A(in3[47]), .ZN(n_0_114));
   INV_X1 i_0_207 (.A(n_0_132), .ZN(n_0_113));
   INV_X1 i_0_208 (.A(in3[63]), .ZN(n_0_122));
   NAND2_X1 i_0_214 (.A1(n_0_112), .A2(n_0_125), .ZN(sum[46]));
   NAND2_X1 i_0_215 (.A1(n_0_123), .A2(n_0_124), .ZN(n_0_112));
   NAND2_X1 i_0_216 (.A1(n_0_128), .A2(n_0_126), .ZN(n_0_123));
   INV_X1 i_0_217 (.A(in2[46]), .ZN(n_0_124));
   NAND3_X1 i_0_218 (.A1(n_0_128), .A2(in2[46]), .A3(n_0_126), .ZN(n_0_125));
   NAND2_X1 i_0_224 (.A1(in1[63]), .A2(n_0_127), .ZN(n_0_126));
   INV_X1 i_0_225 (.A(in3[46]), .ZN(n_0_127));
   NAND2_X1 i_0_226 (.A1(n_0_133), .A2(in3[46]), .ZN(n_0_128));
   NOR2_X1 i_0_227 (.A1(n_0_129), .A2(n_0_131), .ZN(sum[63]));
   INV_X1 i_0_228 (.A(n_0_130), .ZN(n_0_129));
   NAND3_X1 i_0_229 (.A1(n_0_143), .A2(in3[63]), .A3(n_0_147), .ZN(n_0_130));
   AOI21_X1 i_0_230 (.A(in3[63]), .B1(n_0_143), .B2(n_0_147), .ZN(n_0_131));
   NAND2_X1 i_0_231 (.A1(n_0_143), .A2(n_0_147), .ZN(n_0_132));
   INV_X1 i_0_232 (.A(in1[63]), .ZN(n_0_133));
   INV_X1 i_0_233 (.A(in2[63]), .ZN(n_0_134));
   NAND2_X1 i_0_234 (.A1(n_0_137), .A2(n_0_135), .ZN(sum[47]));
   NAND2_X1 i_0_235 (.A1(n_0_143), .A2(n_0_136), .ZN(n_0_135));
   AOI21_X1 i_0_236 (.A(in3[47]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_136));
   OAI21_X1 i_0_237 (.A(in3[47]), .B1(n_0_146), .B2(n_0_145), .ZN(n_0_137));
   NAND2_X1 i_0_238 (.A1(n_0_140), .A2(n_0_138), .ZN(sum[48]));
   NAND2_X1 i_0_239 (.A1(n_0_143), .A2(n_0_139), .ZN(n_0_138));
   AOI21_X1 i_0_240 (.A(in3[48]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_139));
   OAI21_X1 i_0_241 (.A(in3[48]), .B1(n_0_146), .B2(n_0_145), .ZN(n_0_140));
   NAND2_X1 i_0_242 (.A1(n_0_144), .A2(n_0_141), .ZN(sum[49]));
   NAND2_X1 i_0_243 (.A1(n_0_143), .A2(n_0_142), .ZN(n_0_141));
   AOI21_X1 i_0_244 (.A(in3[49]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_142));
   NAND2_X1 i_0_245 (.A1(n_0_133), .A2(n_0_134), .ZN(n_0_143));
   OAI21_X1 i_0_246 (.A(in3[49]), .B1(n_0_146), .B2(n_0_145), .ZN(n_0_144));
   NOR2_X1 i_0_247 (.A1(in1[63]), .A2(in2[63]), .ZN(n_0_145));
   INV_X1 i_0_248 (.A(n_0_147), .ZN(n_0_146));
   NAND2_X1 i_0_249 (.A1(in1[63]), .A2(in2[63]), .ZN(n_0_147));
endmodule

module CSA__3_5(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;

   AND2_X1 i_0_0 (.A1(in2[14]), .A2(in1[14]), .ZN(c[15]));
   AND2_X1 i_0_1 (.A1(in2[15]), .A2(in1[15]), .ZN(c[16]));
   AND2_X1 i_0_2 (.A1(in2[16]), .A2(in1[16]), .ZN(c[17]));
   NAND2_X1 i_0_3 (.A1(n_0_1), .A2(n_0_0), .ZN(c[18]));
   OAI21_X1 i_0_4 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_0));
   NAND2_X1 i_0_5 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_1));
   NAND2_X1 i_0_6 (.A1(n_0_3), .A2(n_0_2), .ZN(c[19]));
   OAI21_X1 i_0_7 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_2));
   NAND2_X1 i_0_8 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_3));
   NAND2_X1 i_0_9 (.A1(n_0_5), .A2(n_0_4), .ZN(c[20]));
   OAI21_X1 i_0_10 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_4));
   NAND2_X1 i_0_11 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_5));
   NAND2_X1 i_0_12 (.A1(n_0_7), .A2(n_0_6), .ZN(c[21]));
   OAI21_X1 i_0_13 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_6));
   NAND2_X1 i_0_14 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_7));
   NAND2_X1 i_0_15 (.A1(n_0_9), .A2(n_0_8), .ZN(c[22]));
   OAI21_X1 i_0_16 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_8));
   NAND2_X1 i_0_17 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_9));
   NAND2_X1 i_0_18 (.A1(n_0_11), .A2(n_0_10), .ZN(c[23]));
   OAI21_X1 i_0_19 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_10));
   NAND2_X1 i_0_20 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_11));
   NAND2_X1 i_0_21 (.A1(n_0_13), .A2(n_0_12), .ZN(c[24]));
   OAI21_X1 i_0_22 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_12));
   NAND2_X1 i_0_23 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_13));
   NAND2_X1 i_0_24 (.A1(n_0_15), .A2(n_0_14), .ZN(c[25]));
   OAI21_X1 i_0_25 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_14));
   NAND2_X1 i_0_26 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_15));
   NAND2_X1 i_0_27 (.A1(n_0_17), .A2(n_0_16), .ZN(c[26]));
   OAI21_X1 i_0_28 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_16));
   NAND2_X1 i_0_29 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_17));
   NAND2_X1 i_0_30 (.A1(n_0_19), .A2(n_0_18), .ZN(c[27]));
   OAI21_X1 i_0_31 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_18));
   NAND2_X1 i_0_32 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_19));
   NAND2_X1 i_0_33 (.A1(n_0_21), .A2(n_0_20), .ZN(c[28]));
   OAI21_X1 i_0_34 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_20));
   NAND2_X1 i_0_35 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_21));
   NAND2_X1 i_0_36 (.A1(n_0_23), .A2(n_0_22), .ZN(c[29]));
   OAI21_X1 i_0_37 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_22));
   NAND2_X1 i_0_38 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_23));
   NAND2_X1 i_0_39 (.A1(n_0_25), .A2(n_0_24), .ZN(c[30]));
   OAI21_X1 i_0_40 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_24));
   NAND2_X1 i_0_41 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_25));
   NAND2_X1 i_0_42 (.A1(n_0_27), .A2(n_0_26), .ZN(c[31]));
   OAI21_X1 i_0_43 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_26));
   NAND2_X1 i_0_44 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_27));
   NAND2_X1 i_0_45 (.A1(n_0_29), .A2(n_0_28), .ZN(c[32]));
   OAI21_X1 i_0_46 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_28));
   NAND2_X1 i_0_47 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_29));
   NAND2_X1 i_0_48 (.A1(n_0_31), .A2(n_0_30), .ZN(c[33]));
   OAI21_X1 i_0_49 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_30));
   NAND2_X1 i_0_50 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_31));
   NAND2_X1 i_0_51 (.A1(n_0_33), .A2(n_0_32), .ZN(c[34]));
   OAI21_X1 i_0_52 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_32));
   NAND2_X1 i_0_53 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_33));
   NAND2_X1 i_0_54 (.A1(n_0_35), .A2(n_0_34), .ZN(c[35]));
   OAI21_X1 i_0_55 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_34));
   NAND2_X1 i_0_56 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_35));
   NAND2_X1 i_0_57 (.A1(n_0_37), .A2(n_0_36), .ZN(c[36]));
   OAI21_X1 i_0_58 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_36));
   NAND2_X1 i_0_59 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_37));
   NAND2_X1 i_0_60 (.A1(n_0_39), .A2(n_0_38), .ZN(c[37]));
   OAI21_X1 i_0_61 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_38));
   NAND2_X1 i_0_62 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_39));
   NAND2_X1 i_0_63 (.A1(n_0_41), .A2(n_0_40), .ZN(c[38]));
   OAI21_X1 i_0_64 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_40));
   NAND2_X1 i_0_65 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_41));
   NAND2_X1 i_0_66 (.A1(n_0_43), .A2(n_0_42), .ZN(c[39]));
   OAI21_X1 i_0_67 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_42));
   NAND2_X1 i_0_68 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_43));
   NAND2_X1 i_0_69 (.A1(n_0_45), .A2(n_0_44), .ZN(c[40]));
   OAI21_X1 i_0_70 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_44));
   NAND2_X1 i_0_71 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_45));
   NAND2_X1 i_0_72 (.A1(n_0_47), .A2(n_0_46), .ZN(c[41]));
   OAI21_X1 i_0_73 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_46));
   NAND2_X1 i_0_74 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_47));
   NAND2_X1 i_0_75 (.A1(n_0_49), .A2(n_0_48), .ZN(c[42]));
   OAI21_X1 i_0_76 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_48));
   NAND2_X1 i_0_77 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_49));
   NAND2_X1 i_0_78 (.A1(n_0_51), .A2(n_0_50), .ZN(c[43]));
   OAI21_X1 i_0_79 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_50));
   NAND2_X1 i_0_80 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_51));
   NAND2_X1 i_0_81 (.A1(n_0_53), .A2(n_0_52), .ZN(c[44]));
   OAI21_X1 i_0_82 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_52));
   NAND2_X1 i_0_83 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_53));
   NAND2_X1 i_0_84 (.A1(n_0_55), .A2(n_0_54), .ZN(c[45]));
   OAI21_X1 i_0_85 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_54));
   NAND2_X1 i_0_86 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_55));
   NAND2_X1 i_0_87 (.A1(n_0_57), .A2(n_0_56), .ZN(c[46]));
   OAI21_X1 i_0_88 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_56));
   NAND2_X1 i_0_89 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_57));
   NAND2_X1 i_0_90 (.A1(n_0_59), .A2(n_0_58), .ZN(c[47]));
   OAI21_X1 i_0_91 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_58));
   NAND2_X1 i_0_92 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_59));
   NAND2_X1 i_0_93 (.A1(n_0_61), .A2(n_0_60), .ZN(c[48]));
   OAI21_X1 i_0_94 (.A(in2[47]), .B1(in3[47]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_95 (.A1(in3[47]), .A2(in1[63]), .ZN(n_0_61));
   NAND2_X1 i_0_96 (.A1(n_0_63), .A2(n_0_62), .ZN(c[49]));
   OAI21_X1 i_0_97 (.A(in2[48]), .B1(in3[48]), .B2(in1[63]), .ZN(n_0_62));
   NAND2_X1 i_0_98 (.A1(in3[48]), .A2(in1[63]), .ZN(n_0_63));
   NAND2_X1 i_0_99 (.A1(n_0_65), .A2(n_0_64), .ZN(c[50]));
   OAI21_X1 i_0_100 (.A(in3[49]), .B1(in1[63]), .B2(in2[49]), .ZN(n_0_64));
   NAND2_X1 i_0_101 (.A1(in2[49]), .A2(in1[63]), .ZN(n_0_65));
   NAND2_X1 i_0_102 (.A1(n_0_67), .A2(n_0_66), .ZN(c[51]));
   OAI21_X1 i_0_103 (.A(in2[50]), .B1(in3[50]), .B2(in1[63]), .ZN(n_0_66));
   NAND2_X1 i_0_104 (.A1(in3[50]), .A2(in1[63]), .ZN(n_0_67));
   NAND2_X1 i_0_105 (.A1(n_0_69), .A2(n_0_68), .ZN(c[52]));
   OAI21_X1 i_0_106 (.A(in2[51]), .B1(in3[51]), .B2(in1[63]), .ZN(n_0_68));
   NAND2_X1 i_0_107 (.A1(in3[51]), .A2(in1[63]), .ZN(n_0_69));
   NAND2_X1 i_0_108 (.A1(n_0_71), .A2(n_0_70), .ZN(c[53]));
   OAI21_X1 i_0_109 (.A(in2[52]), .B1(in3[52]), .B2(in1[63]), .ZN(n_0_70));
   NAND2_X1 i_0_110 (.A1(in3[52]), .A2(in1[63]), .ZN(n_0_71));
   NAND2_X1 i_0_111 (.A1(n_0_73), .A2(n_0_72), .ZN(c[54]));
   OAI21_X1 i_0_112 (.A(in2[53]), .B1(in3[53]), .B2(in1[63]), .ZN(n_0_72));
   NAND2_X1 i_0_113 (.A1(in3[53]), .A2(in1[63]), .ZN(n_0_73));
   NAND2_X1 i_0_114 (.A1(n_0_76), .A2(n_0_74), .ZN(c[55]));
   OAI21_X1 i_0_115 (.A(in3[54]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_74));
   NAND2_X1 i_0_116 (.A1(n_0_76), .A2(n_0_75), .ZN(c[63]));
   OAI21_X1 i_0_117 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_75));
   NAND2_X1 i_0_118 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_76));
   XOR2_X1 i_0_119 (.A(in2[14]), .B(in1[14]), .Z(sum[14]));
   XOR2_X1 i_0_120 (.A(in2[15]), .B(in1[15]), .Z(sum[15]));
   XOR2_X1 i_0_121 (.A(in2[16]), .B(in1[16]), .Z(sum[16]));
   XNOR2_X1 i_0_122 (.A(in2[17]), .B(n_0_77), .ZN(sum[17]));
   XNOR2_X1 i_0_123 (.A(in3[17]), .B(in1[17]), .ZN(n_0_77));
   XNOR2_X1 i_0_124 (.A(in2[18]), .B(n_0_78), .ZN(sum[18]));
   XNOR2_X1 i_0_125 (.A(in3[18]), .B(in1[18]), .ZN(n_0_78));
   XNOR2_X1 i_0_126 (.A(in2[19]), .B(n_0_79), .ZN(sum[19]));
   XNOR2_X1 i_0_127 (.A(in3[19]), .B(in1[19]), .ZN(n_0_79));
   XNOR2_X1 i_0_128 (.A(in2[20]), .B(n_0_80), .ZN(sum[20]));
   XNOR2_X1 i_0_129 (.A(in3[20]), .B(in1[20]), .ZN(n_0_80));
   XNOR2_X1 i_0_130 (.A(in2[21]), .B(n_0_81), .ZN(sum[21]));
   XNOR2_X1 i_0_131 (.A(in3[21]), .B(in1[21]), .ZN(n_0_81));
   XNOR2_X1 i_0_132 (.A(in2[22]), .B(n_0_82), .ZN(sum[22]));
   XNOR2_X1 i_0_133 (.A(in3[22]), .B(in1[22]), .ZN(n_0_82));
   XNOR2_X1 i_0_134 (.A(in2[23]), .B(n_0_83), .ZN(sum[23]));
   XNOR2_X1 i_0_135 (.A(in3[23]), .B(in1[23]), .ZN(n_0_83));
   XNOR2_X1 i_0_136 (.A(in2[24]), .B(n_0_84), .ZN(sum[24]));
   XNOR2_X1 i_0_137 (.A(in3[24]), .B(in1[24]), .ZN(n_0_84));
   XNOR2_X1 i_0_138 (.A(in2[25]), .B(n_0_85), .ZN(sum[25]));
   XNOR2_X1 i_0_139 (.A(in3[25]), .B(in1[25]), .ZN(n_0_85));
   XNOR2_X1 i_0_140 (.A(in2[26]), .B(n_0_86), .ZN(sum[26]));
   XNOR2_X1 i_0_141 (.A(in3[26]), .B(in1[26]), .ZN(n_0_86));
   XNOR2_X1 i_0_142 (.A(in2[27]), .B(n_0_87), .ZN(sum[27]));
   XNOR2_X1 i_0_143 (.A(in3[27]), .B(in1[27]), .ZN(n_0_87));
   XNOR2_X1 i_0_144 (.A(in2[28]), .B(n_0_88), .ZN(sum[28]));
   XNOR2_X1 i_0_145 (.A(in3[28]), .B(in1[28]), .ZN(n_0_88));
   XNOR2_X1 i_0_146 (.A(in2[29]), .B(n_0_89), .ZN(sum[29]));
   XNOR2_X1 i_0_147 (.A(in3[29]), .B(in1[29]), .ZN(n_0_89));
   XNOR2_X1 i_0_148 (.A(in2[30]), .B(n_0_90), .ZN(sum[30]));
   XNOR2_X1 i_0_149 (.A(in3[30]), .B(in1[30]), .ZN(n_0_90));
   XNOR2_X1 i_0_150 (.A(in2[31]), .B(n_0_91), .ZN(sum[31]));
   XNOR2_X1 i_0_151 (.A(in3[31]), .B(in1[31]), .ZN(n_0_91));
   XNOR2_X1 i_0_152 (.A(in2[32]), .B(n_0_92), .ZN(sum[32]));
   XNOR2_X1 i_0_153 (.A(in3[32]), .B(in1[32]), .ZN(n_0_92));
   XNOR2_X1 i_0_154 (.A(in2[33]), .B(n_0_93), .ZN(sum[33]));
   XNOR2_X1 i_0_155 (.A(in3[33]), .B(in1[33]), .ZN(n_0_93));
   XNOR2_X1 i_0_156 (.A(in2[34]), .B(n_0_94), .ZN(sum[34]));
   XNOR2_X1 i_0_157 (.A(in3[34]), .B(in1[34]), .ZN(n_0_94));
   XNOR2_X1 i_0_158 (.A(in2[35]), .B(n_0_95), .ZN(sum[35]));
   XNOR2_X1 i_0_159 (.A(in3[35]), .B(in1[35]), .ZN(n_0_95));
   XNOR2_X1 i_0_160 (.A(in2[36]), .B(n_0_96), .ZN(sum[36]));
   XNOR2_X1 i_0_161 (.A(in3[36]), .B(in1[36]), .ZN(n_0_96));
   XNOR2_X1 i_0_162 (.A(in2[37]), .B(n_0_97), .ZN(sum[37]));
   XNOR2_X1 i_0_163 (.A(in3[37]), .B(in1[37]), .ZN(n_0_97));
   XNOR2_X1 i_0_164 (.A(in2[38]), .B(n_0_98), .ZN(sum[38]));
   XNOR2_X1 i_0_165 (.A(in3[38]), .B(in1[38]), .ZN(n_0_98));
   XNOR2_X1 i_0_166 (.A(in2[39]), .B(n_0_99), .ZN(sum[39]));
   XNOR2_X1 i_0_167 (.A(in3[39]), .B(in1[39]), .ZN(n_0_99));
   XNOR2_X1 i_0_168 (.A(in2[40]), .B(n_0_100), .ZN(sum[40]));
   XNOR2_X1 i_0_169 (.A(in3[40]), .B(in1[40]), .ZN(n_0_100));
   XNOR2_X1 i_0_170 (.A(in2[41]), .B(n_0_101), .ZN(sum[41]));
   XNOR2_X1 i_0_171 (.A(in3[41]), .B(in1[41]), .ZN(n_0_101));
   XNOR2_X1 i_0_172 (.A(in2[42]), .B(n_0_102), .ZN(sum[42]));
   XNOR2_X1 i_0_173 (.A(in3[42]), .B(in1[42]), .ZN(n_0_102));
   XNOR2_X1 i_0_174 (.A(in2[43]), .B(n_0_103), .ZN(sum[43]));
   XNOR2_X1 i_0_175 (.A(in3[43]), .B(in1[43]), .ZN(n_0_103));
   XNOR2_X1 i_0_176 (.A(in2[44]), .B(n_0_104), .ZN(sum[44]));
   XNOR2_X1 i_0_177 (.A(in3[44]), .B(in1[44]), .ZN(n_0_104));
   XNOR2_X1 i_0_178 (.A(in2[45]), .B(n_0_105), .ZN(sum[45]));
   XNOR2_X1 i_0_179 (.A(in3[45]), .B(in1[45]), .ZN(n_0_105));
   XNOR2_X1 i_0_180 (.A(in2[46]), .B(n_0_106), .ZN(sum[46]));
   XNOR2_X1 i_0_181 (.A(in3[46]), .B(in1[46]), .ZN(n_0_106));
   XNOR2_X1 i_0_182 (.A(in2[47]), .B(n_0_107), .ZN(sum[47]));
   XNOR2_X1 i_0_183 (.A(in3[47]), .B(in1[63]), .ZN(n_0_107));
   XNOR2_X1 i_0_184 (.A(in2[48]), .B(n_0_108), .ZN(sum[48]));
   XNOR2_X1 i_0_185 (.A(in3[48]), .B(in1[63]), .ZN(n_0_108));
   XNOR2_X1 i_0_186 (.A(in2[49]), .B(n_0_109), .ZN(sum[49]));
   XNOR2_X1 i_0_187 (.A(in3[49]), .B(in1[63]), .ZN(n_0_109));
   XNOR2_X1 i_0_188 (.A(in2[50]), .B(n_0_110), .ZN(sum[50]));
   XNOR2_X1 i_0_189 (.A(in3[50]), .B(in1[63]), .ZN(n_0_110));
   XNOR2_X1 i_0_190 (.A(in2[51]), .B(n_0_111), .ZN(sum[51]));
   XNOR2_X1 i_0_191 (.A(in3[51]), .B(in1[63]), .ZN(n_0_111));
   XNOR2_X1 i_0_192 (.A(in2[52]), .B(n_0_112), .ZN(sum[52]));
   XNOR2_X1 i_0_193 (.A(in3[52]), .B(in1[63]), .ZN(n_0_112));
   XNOR2_X1 i_0_194 (.A(in2[53]), .B(n_0_113), .ZN(sum[53]));
   XNOR2_X1 i_0_195 (.A(in3[53]), .B(in1[63]), .ZN(n_0_113));
   XOR2_X1 i_0_196 (.A(in3[54]), .B(n_0_114), .Z(sum[54]));
   XOR2_X1 i_0_197 (.A(in3[63]), .B(n_0_114), .Z(sum[63]));
   XOR2_X1 i_0_198 (.A(in2[63]), .B(in1[63]), .Z(n_0_114));
endmodule

module CSA__3_8(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;

   AND2_X1 i_0_0 (.A1(in2[16]), .A2(in1[16]), .ZN(c[17]));
   AND2_X1 i_0_1 (.A1(in2[17]), .A2(in1[17]), .ZN(c[18]));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_0), .ZN(c[19]));
   OAI21_X1 i_0_3 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_0));
   NAND2_X1 i_0_4 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .ZN(c[20]));
   OAI21_X1 i_0_6 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_2));
   NAND2_X1 i_0_7 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_4), .ZN(c[21]));
   OAI21_X1 i_0_9 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_4));
   NAND2_X1 i_0_10 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(n_0_7), .A2(n_0_6), .ZN(c[22]));
   OAI21_X1 i_0_12 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_6));
   NAND2_X1 i_0_13 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_7));
   NAND2_X1 i_0_14 (.A1(n_0_9), .A2(n_0_8), .ZN(c[23]));
   OAI21_X1 i_0_15 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_8));
   NAND2_X1 i_0_16 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_9));
   NAND2_X1 i_0_17 (.A1(n_0_11), .A2(n_0_10), .ZN(c[24]));
   OAI21_X1 i_0_18 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_10));
   NAND2_X1 i_0_19 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_11));
   NAND2_X1 i_0_20 (.A1(n_0_13), .A2(n_0_12), .ZN(c[25]));
   OAI21_X1 i_0_21 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_12));
   NAND2_X1 i_0_22 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_13));
   NAND2_X1 i_0_23 (.A1(n_0_15), .A2(n_0_14), .ZN(c[26]));
   OAI21_X1 i_0_24 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_14));
   NAND2_X1 i_0_25 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_15));
   NAND2_X1 i_0_26 (.A1(n_0_17), .A2(n_0_16), .ZN(c[27]));
   OAI21_X1 i_0_27 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_16));
   NAND2_X1 i_0_28 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_17));
   NAND2_X1 i_0_29 (.A1(n_0_19), .A2(n_0_18), .ZN(c[28]));
   OAI21_X1 i_0_30 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_18));
   NAND2_X1 i_0_31 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_19));
   NAND2_X1 i_0_32 (.A1(n_0_21), .A2(n_0_20), .ZN(c[29]));
   OAI21_X1 i_0_33 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_20));
   NAND2_X1 i_0_34 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_21));
   NAND2_X1 i_0_35 (.A1(n_0_23), .A2(n_0_22), .ZN(c[30]));
   OAI21_X1 i_0_36 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_22));
   NAND2_X1 i_0_37 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_23));
   NAND2_X1 i_0_38 (.A1(n_0_25), .A2(n_0_24), .ZN(c[31]));
   OAI21_X1 i_0_39 (.A(in1[30]), .B1(in3[30]), .B2(in2[30]), .ZN(n_0_24));
   NAND2_X1 i_0_40 (.A1(in2[30]), .A2(in3[30]), .ZN(n_0_25));
   NAND2_X1 i_0_41 (.A1(n_0_27), .A2(n_0_26), .ZN(c[32]));
   OAI21_X1 i_0_42 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_26));
   NAND2_X1 i_0_43 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_27));
   NAND2_X1 i_0_44 (.A1(n_0_29), .A2(n_0_28), .ZN(c[33]));
   OAI21_X1 i_0_45 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_28));
   NAND2_X1 i_0_46 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_29));
   NAND2_X1 i_0_47 (.A1(n_0_31), .A2(n_0_30), .ZN(c[34]));
   OAI21_X1 i_0_48 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_30));
   NAND2_X1 i_0_49 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_31));
   NAND2_X1 i_0_50 (.A1(n_0_33), .A2(n_0_32), .ZN(c[35]));
   OAI21_X1 i_0_51 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_32));
   NAND2_X1 i_0_52 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_33));
   NAND2_X1 i_0_53 (.A1(n_0_35), .A2(n_0_34), .ZN(c[36]));
   OAI21_X1 i_0_54 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_34));
   NAND2_X1 i_0_55 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_35));
   NAND2_X1 i_0_56 (.A1(n_0_37), .A2(n_0_36), .ZN(c[37]));
   OAI21_X1 i_0_57 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_36));
   NAND2_X1 i_0_58 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_37));
   NAND2_X1 i_0_59 (.A1(n_0_39), .A2(n_0_38), .ZN(c[38]));
   OAI21_X1 i_0_60 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_38));
   NAND2_X1 i_0_61 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_39));
   NAND2_X1 i_0_62 (.A1(n_0_41), .A2(n_0_40), .ZN(c[39]));
   OAI21_X1 i_0_63 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_40));
   NAND2_X1 i_0_64 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_41));
   NAND2_X1 i_0_65 (.A1(n_0_43), .A2(n_0_42), .ZN(c[40]));
   OAI21_X1 i_0_66 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_42));
   NAND2_X1 i_0_67 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_43));
   NAND2_X1 i_0_68 (.A1(n_0_45), .A2(n_0_44), .ZN(c[41]));
   OAI21_X1 i_0_69 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_44));
   NAND2_X1 i_0_70 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_45));
   NAND2_X1 i_0_71 (.A1(n_0_47), .A2(n_0_46), .ZN(c[42]));
   OAI21_X1 i_0_72 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_46));
   NAND2_X1 i_0_73 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_47));
   NAND2_X1 i_0_74 (.A1(n_0_49), .A2(n_0_48), .ZN(c[43]));
   OAI21_X1 i_0_75 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_48));
   NAND2_X1 i_0_76 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_49));
   NAND2_X1 i_0_77 (.A1(n_0_51), .A2(n_0_50), .ZN(c[44]));
   OAI21_X1 i_0_78 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_50));
   NAND2_X1 i_0_79 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_51));
   NAND2_X1 i_0_80 (.A1(n_0_53), .A2(n_0_52), .ZN(c[45]));
   OAI21_X1 i_0_81 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_52));
   NAND2_X1 i_0_82 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_53));
   NAND2_X1 i_0_83 (.A1(n_0_55), .A2(n_0_54), .ZN(c[46]));
   OAI21_X1 i_0_84 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_54));
   NAND2_X1 i_0_85 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_55));
   NAND2_X1 i_0_86 (.A1(n_0_57), .A2(n_0_56), .ZN(c[47]));
   OAI21_X1 i_0_87 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_56));
   NAND2_X1 i_0_88 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_57));
   NAND2_X1 i_0_89 (.A1(n_0_59), .A2(n_0_58), .ZN(c[48]));
   OAI21_X1 i_0_90 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_58));
   NAND2_X1 i_0_91 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_59));
   NAND2_X1 i_0_92 (.A1(n_0_61), .A2(n_0_60), .ZN(c[49]));
   OAI21_X1 i_0_93 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_60));
   NAND2_X1 i_0_94 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(n_0_63), .A2(n_0_62), .ZN(c[50]));
   OAI21_X1 i_0_96 (.A(in2[49]), .B1(in3[49]), .B2(in1[63]), .ZN(n_0_62));
   NAND2_X1 i_0_97 (.A1(in3[49]), .A2(in1[63]), .ZN(n_0_63));
   AOI21_X1 i_0_98 (.A(n_0_65), .B1(n_0_64), .B2(n_0_99), .ZN(c[51]));
   AOI21_X1 i_0_99 (.A(n_0_65), .B1(n_0_64), .B2(n_0_100), .ZN(c[52]));
   AOI21_X1 i_0_100 (.A(n_0_65), .B1(n_0_64), .B2(n_0_101), .ZN(c[53]));
   AOI21_X1 i_0_101 (.A(n_0_65), .B1(n_0_64), .B2(n_0_102), .ZN(c[54]));
   AOI21_X1 i_0_102 (.A(n_0_65), .B1(n_0_64), .B2(n_0_103), .ZN(c[63]));
   NAND2_X1 i_0_103 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_64));
   NOR2_X1 i_0_104 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_65));
   XOR2_X1 i_0_105 (.A(in2[16]), .B(in1[16]), .Z(sum[16]));
   XOR2_X1 i_0_106 (.A(in2[17]), .B(in1[17]), .Z(sum[17]));
   XNOR2_X1 i_0_107 (.A(in2[18]), .B(n_0_66), .ZN(sum[18]));
   XNOR2_X1 i_0_108 (.A(in3[18]), .B(in1[18]), .ZN(n_0_66));
   XNOR2_X1 i_0_109 (.A(in2[19]), .B(n_0_67), .ZN(sum[19]));
   XNOR2_X1 i_0_110 (.A(in3[19]), .B(in1[19]), .ZN(n_0_67));
   XNOR2_X1 i_0_111 (.A(in2[20]), .B(n_0_68), .ZN(sum[20]));
   XNOR2_X1 i_0_112 (.A(in3[20]), .B(in1[20]), .ZN(n_0_68));
   XNOR2_X1 i_0_113 (.A(in2[21]), .B(n_0_69), .ZN(sum[21]));
   XNOR2_X1 i_0_114 (.A(in3[21]), .B(in1[21]), .ZN(n_0_69));
   XNOR2_X1 i_0_115 (.A(in2[22]), .B(n_0_70), .ZN(sum[22]));
   XNOR2_X1 i_0_116 (.A(in3[22]), .B(in1[22]), .ZN(n_0_70));
   XNOR2_X1 i_0_117 (.A(in2[23]), .B(n_0_71), .ZN(sum[23]));
   XNOR2_X1 i_0_118 (.A(in3[23]), .B(in1[23]), .ZN(n_0_71));
   XNOR2_X1 i_0_119 (.A(in2[24]), .B(n_0_72), .ZN(sum[24]));
   XNOR2_X1 i_0_120 (.A(in3[24]), .B(in1[24]), .ZN(n_0_72));
   XNOR2_X1 i_0_121 (.A(in2[25]), .B(n_0_73), .ZN(sum[25]));
   XNOR2_X1 i_0_122 (.A(in3[25]), .B(in1[25]), .ZN(n_0_73));
   XNOR2_X1 i_0_123 (.A(in2[26]), .B(n_0_74), .ZN(sum[26]));
   XNOR2_X1 i_0_124 (.A(in3[26]), .B(in1[26]), .ZN(n_0_74));
   XNOR2_X1 i_0_125 (.A(in2[27]), .B(n_0_75), .ZN(sum[27]));
   XNOR2_X1 i_0_126 (.A(in3[27]), .B(in1[27]), .ZN(n_0_75));
   XNOR2_X1 i_0_127 (.A(in2[28]), .B(n_0_76), .ZN(sum[28]));
   XNOR2_X1 i_0_128 (.A(in3[28]), .B(in1[28]), .ZN(n_0_76));
   XNOR2_X1 i_0_129 (.A(in2[29]), .B(n_0_77), .ZN(sum[29]));
   XNOR2_X1 i_0_130 (.A(in3[29]), .B(in1[29]), .ZN(n_0_77));
   XNOR2_X1 i_0_131 (.A(in2[30]), .B(n_0_78), .ZN(sum[30]));
   XNOR2_X1 i_0_132 (.A(in3[30]), .B(in1[30]), .ZN(n_0_78));
   XNOR2_X1 i_0_133 (.A(in2[31]), .B(n_0_79), .ZN(sum[31]));
   XNOR2_X1 i_0_134 (.A(in3[31]), .B(in1[31]), .ZN(n_0_79));
   XNOR2_X1 i_0_135 (.A(in2[32]), .B(n_0_80), .ZN(sum[32]));
   XNOR2_X1 i_0_136 (.A(in3[32]), .B(in1[32]), .ZN(n_0_80));
   XNOR2_X1 i_0_137 (.A(in2[33]), .B(n_0_81), .ZN(sum[33]));
   XNOR2_X1 i_0_138 (.A(in3[33]), .B(in1[33]), .ZN(n_0_81));
   XNOR2_X1 i_0_139 (.A(in2[34]), .B(n_0_82), .ZN(sum[34]));
   XNOR2_X1 i_0_140 (.A(in3[34]), .B(in1[34]), .ZN(n_0_82));
   XNOR2_X1 i_0_141 (.A(in2[35]), .B(n_0_83), .ZN(sum[35]));
   XNOR2_X1 i_0_142 (.A(in3[35]), .B(in1[35]), .ZN(n_0_83));
   XNOR2_X1 i_0_143 (.A(in2[36]), .B(n_0_84), .ZN(sum[36]));
   XNOR2_X1 i_0_144 (.A(in3[36]), .B(in1[36]), .ZN(n_0_84));
   XNOR2_X1 i_0_145 (.A(in2[37]), .B(n_0_85), .ZN(sum[37]));
   XNOR2_X1 i_0_146 (.A(in3[37]), .B(in1[37]), .ZN(n_0_85));
   XNOR2_X1 i_0_147 (.A(in2[38]), .B(n_0_86), .ZN(sum[38]));
   XNOR2_X1 i_0_148 (.A(in3[38]), .B(in1[38]), .ZN(n_0_86));
   XNOR2_X1 i_0_149 (.A(in2[39]), .B(n_0_87), .ZN(sum[39]));
   XNOR2_X1 i_0_150 (.A(in3[39]), .B(in1[39]), .ZN(n_0_87));
   XNOR2_X1 i_0_151 (.A(in2[40]), .B(n_0_88), .ZN(sum[40]));
   XNOR2_X1 i_0_152 (.A(in3[40]), .B(in1[40]), .ZN(n_0_88));
   XNOR2_X1 i_0_153 (.A(in2[41]), .B(n_0_89), .ZN(sum[41]));
   XNOR2_X1 i_0_154 (.A(in3[41]), .B(in1[41]), .ZN(n_0_89));
   XNOR2_X1 i_0_155 (.A(in2[42]), .B(n_0_90), .ZN(sum[42]));
   XNOR2_X1 i_0_156 (.A(in3[42]), .B(in1[42]), .ZN(n_0_90));
   XNOR2_X1 i_0_157 (.A(in2[43]), .B(n_0_91), .ZN(sum[43]));
   XNOR2_X1 i_0_158 (.A(in3[43]), .B(in1[43]), .ZN(n_0_91));
   XNOR2_X1 i_0_159 (.A(in2[44]), .B(n_0_92), .ZN(sum[44]));
   XNOR2_X1 i_0_160 (.A(in3[44]), .B(in1[44]), .ZN(n_0_92));
   XNOR2_X1 i_0_161 (.A(in2[45]), .B(n_0_93), .ZN(sum[45]));
   XNOR2_X1 i_0_162 (.A(in3[45]), .B(in1[45]), .ZN(n_0_93));
   XNOR2_X1 i_0_163 (.A(in2[46]), .B(n_0_94), .ZN(sum[46]));
   XNOR2_X1 i_0_164 (.A(in3[46]), .B(in1[46]), .ZN(n_0_94));
   XNOR2_X1 i_0_165 (.A(in2[47]), .B(n_0_95), .ZN(sum[47]));
   XNOR2_X1 i_0_166 (.A(in3[47]), .B(in1[47]), .ZN(n_0_95));
   XNOR2_X1 i_0_167 (.A(in2[48]), .B(n_0_96), .ZN(sum[48]));
   XNOR2_X1 i_0_168 (.A(in3[48]), .B(in1[48]), .ZN(n_0_96));
   XNOR2_X1 i_0_169 (.A(in2[49]), .B(n_0_97), .ZN(sum[49]));
   XNOR2_X1 i_0_170 (.A(in3[49]), .B(in1[63]), .ZN(n_0_97));
   XNOR2_X1 i_0_171 (.A(n_0_99), .B(n_0_98), .ZN(sum[50]));
   XNOR2_X1 i_0_172 (.A(n_0_100), .B(n_0_98), .ZN(sum[51]));
   XNOR2_X1 i_0_173 (.A(n_0_101), .B(n_0_98), .ZN(sum[52]));
   XNOR2_X1 i_0_174 (.A(n_0_102), .B(n_0_98), .ZN(sum[53]));
   XNOR2_X1 i_0_175 (.A(n_0_103), .B(n_0_98), .ZN(sum[63]));
   XOR2_X1 i_0_176 (.A(in2[63]), .B(in1[63]), .Z(n_0_98));
   INV_X1 i_0_177 (.A(in3[50]), .ZN(n_0_99));
   INV_X1 i_0_178 (.A(in3[51]), .ZN(n_0_100));
   INV_X1 i_0_179 (.A(in3[52]), .ZN(n_0_101));
   INV_X1 i_0_180 (.A(in3[53]), .ZN(n_0_102));
   INV_X1 i_0_181 (.A(in3[63]), .ZN(n_0_103));
endmodule

module CSA__3_11(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;

   AND2_X1 i_0_0 (.A1(in2[20]), .A2(in1[20]), .ZN(c[21]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[22]));
   OAI21_X1 i_0_2 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[23]));
   OAI21_X1 i_0_5 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[24]));
   OAI21_X1 i_0_8 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[25]));
   OAI21_X1 i_0_11 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[26]));
   OAI21_X1 i_0_14 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[27]));
   OAI21_X1 i_0_17 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[28]));
   OAI21_X1 i_0_20 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[29]));
   OAI21_X1 i_0_23 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[30]));
   OAI21_X1 i_0_26 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[31]));
   OAI21_X1 i_0_29 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[32]));
   OAI21_X1 i_0_32 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[33]));
   OAI21_X1 i_0_35 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[34]));
   OAI21_X1 i_0_38 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[35]));
   OAI21_X1 i_0_41 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[36]));
   OAI21_X1 i_0_44 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[37]));
   OAI21_X1 i_0_47 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[38]));
   OAI21_X1 i_0_50 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[39]));
   OAI21_X1 i_0_53 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[40]));
   OAI21_X1 i_0_56 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[41]));
   OAI21_X1 i_0_59 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[42]));
   OAI21_X1 i_0_62 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[43]));
   OAI21_X1 i_0_65 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[44]));
   OAI21_X1 i_0_68 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[45]));
   OAI21_X1 i_0_71 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[46]));
   OAI21_X1 i_0_74 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[47]));
   OAI21_X1 i_0_77 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[48]));
   OAI21_X1 i_0_80 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[49]));
   OAI21_X1 i_0_83 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[50]));
   OAI21_X1 i_0_86 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[51]));
   OAI21_X1 i_0_89 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_61), .A2(n_0_60), .ZN(c[52]));
   OAI21_X1 i_0_92 (.A(in2[51]), .B1(in3[51]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(in3[51]), .A2(in1[63]), .ZN(n_0_61));
   AOI21_X1 i_0_94 (.A(n_0_63), .B1(n_0_62), .B2(n_0_96), .ZN(c[53]));
   AOI21_X1 i_0_95 (.A(n_0_63), .B1(n_0_62), .B2(n_0_97), .ZN(c[54]));
   AOI21_X1 i_0_96 (.A(n_0_63), .B1(n_0_62), .B2(n_0_98), .ZN(c[63]));
   NAND2_X1 i_0_97 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   NOR2_X1 i_0_98 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_63));
   XOR2_X1 i_0_99 (.A(in2[20]), .B(in1[20]), .Z(sum[20]));
   XNOR2_X1 i_0_100 (.A(in2[21]), .B(n_0_64), .ZN(sum[21]));
   XNOR2_X1 i_0_101 (.A(in3[21]), .B(in1[21]), .ZN(n_0_64));
   XNOR2_X1 i_0_102 (.A(in2[22]), .B(n_0_65), .ZN(sum[22]));
   XNOR2_X1 i_0_103 (.A(in3[22]), .B(in1[22]), .ZN(n_0_65));
   XNOR2_X1 i_0_104 (.A(in2[23]), .B(n_0_66), .ZN(sum[23]));
   XNOR2_X1 i_0_105 (.A(in3[23]), .B(in1[23]), .ZN(n_0_66));
   XNOR2_X1 i_0_106 (.A(in2[24]), .B(n_0_67), .ZN(sum[24]));
   XNOR2_X1 i_0_107 (.A(in3[24]), .B(in1[24]), .ZN(n_0_67));
   XNOR2_X1 i_0_108 (.A(in2[25]), .B(n_0_68), .ZN(sum[25]));
   XNOR2_X1 i_0_109 (.A(in3[25]), .B(in1[25]), .ZN(n_0_68));
   XNOR2_X1 i_0_110 (.A(in2[26]), .B(n_0_69), .ZN(sum[26]));
   XNOR2_X1 i_0_111 (.A(in3[26]), .B(in1[26]), .ZN(n_0_69));
   XNOR2_X1 i_0_112 (.A(in2[27]), .B(n_0_70), .ZN(sum[27]));
   XNOR2_X1 i_0_113 (.A(in3[27]), .B(in1[27]), .ZN(n_0_70));
   XNOR2_X1 i_0_114 (.A(in2[28]), .B(n_0_71), .ZN(sum[28]));
   XNOR2_X1 i_0_115 (.A(in3[28]), .B(in1[28]), .ZN(n_0_71));
   XNOR2_X1 i_0_116 (.A(in2[29]), .B(n_0_72), .ZN(sum[29]));
   XNOR2_X1 i_0_117 (.A(in3[29]), .B(in1[29]), .ZN(n_0_72));
   XNOR2_X1 i_0_118 (.A(in2[30]), .B(n_0_73), .ZN(sum[30]));
   XNOR2_X1 i_0_119 (.A(in3[30]), .B(in1[30]), .ZN(n_0_73));
   XNOR2_X1 i_0_120 (.A(in2[31]), .B(n_0_74), .ZN(sum[31]));
   XNOR2_X1 i_0_121 (.A(in3[31]), .B(in1[31]), .ZN(n_0_74));
   XNOR2_X1 i_0_122 (.A(in2[32]), .B(n_0_75), .ZN(sum[32]));
   XNOR2_X1 i_0_123 (.A(in3[32]), .B(in1[32]), .ZN(n_0_75));
   XNOR2_X1 i_0_124 (.A(in2[33]), .B(n_0_76), .ZN(sum[33]));
   XNOR2_X1 i_0_125 (.A(in3[33]), .B(in1[33]), .ZN(n_0_76));
   XNOR2_X1 i_0_126 (.A(in2[34]), .B(n_0_77), .ZN(sum[34]));
   XNOR2_X1 i_0_127 (.A(in3[34]), .B(in1[34]), .ZN(n_0_77));
   XNOR2_X1 i_0_128 (.A(in2[35]), .B(n_0_78), .ZN(sum[35]));
   XNOR2_X1 i_0_129 (.A(in3[35]), .B(in1[35]), .ZN(n_0_78));
   XNOR2_X1 i_0_130 (.A(in2[36]), .B(n_0_79), .ZN(sum[36]));
   XNOR2_X1 i_0_131 (.A(in3[36]), .B(in1[36]), .ZN(n_0_79));
   XNOR2_X1 i_0_132 (.A(in2[37]), .B(n_0_80), .ZN(sum[37]));
   XNOR2_X1 i_0_133 (.A(in3[37]), .B(in1[37]), .ZN(n_0_80));
   XNOR2_X1 i_0_134 (.A(in2[38]), .B(n_0_81), .ZN(sum[38]));
   XNOR2_X1 i_0_135 (.A(in3[38]), .B(in1[38]), .ZN(n_0_81));
   XNOR2_X1 i_0_136 (.A(in2[39]), .B(n_0_82), .ZN(sum[39]));
   XNOR2_X1 i_0_137 (.A(in3[39]), .B(in1[39]), .ZN(n_0_82));
   XNOR2_X1 i_0_138 (.A(in2[40]), .B(n_0_83), .ZN(sum[40]));
   XNOR2_X1 i_0_139 (.A(in3[40]), .B(in1[40]), .ZN(n_0_83));
   XNOR2_X1 i_0_140 (.A(in2[41]), .B(n_0_84), .ZN(sum[41]));
   XNOR2_X1 i_0_141 (.A(in3[41]), .B(in1[41]), .ZN(n_0_84));
   XNOR2_X1 i_0_142 (.A(in2[42]), .B(n_0_85), .ZN(sum[42]));
   XNOR2_X1 i_0_143 (.A(in3[42]), .B(in1[42]), .ZN(n_0_85));
   XNOR2_X1 i_0_144 (.A(in2[43]), .B(n_0_86), .ZN(sum[43]));
   XNOR2_X1 i_0_145 (.A(in3[43]), .B(in1[43]), .ZN(n_0_86));
   XNOR2_X1 i_0_146 (.A(in2[44]), .B(n_0_87), .ZN(sum[44]));
   XNOR2_X1 i_0_147 (.A(in3[44]), .B(in1[44]), .ZN(n_0_87));
   XNOR2_X1 i_0_148 (.A(in2[45]), .B(n_0_88), .ZN(sum[45]));
   XNOR2_X1 i_0_149 (.A(in3[45]), .B(in1[45]), .ZN(n_0_88));
   XNOR2_X1 i_0_150 (.A(in2[46]), .B(n_0_89), .ZN(sum[46]));
   XNOR2_X1 i_0_151 (.A(in3[46]), .B(in1[46]), .ZN(n_0_89));
   XNOR2_X1 i_0_152 (.A(in2[47]), .B(n_0_90), .ZN(sum[47]));
   XNOR2_X1 i_0_153 (.A(in3[47]), .B(in1[47]), .ZN(n_0_90));
   XNOR2_X1 i_0_154 (.A(in2[48]), .B(n_0_91), .ZN(sum[48]));
   XNOR2_X1 i_0_155 (.A(in3[48]), .B(in1[48]), .ZN(n_0_91));
   XNOR2_X1 i_0_156 (.A(in2[49]), .B(n_0_92), .ZN(sum[49]));
   XNOR2_X1 i_0_157 (.A(in3[49]), .B(in1[49]), .ZN(n_0_92));
   XNOR2_X1 i_0_158 (.A(in2[50]), .B(n_0_93), .ZN(sum[50]));
   XNOR2_X1 i_0_159 (.A(in3[50]), .B(in1[50]), .ZN(n_0_93));
   XNOR2_X1 i_0_160 (.A(in2[51]), .B(n_0_94), .ZN(sum[51]));
   XNOR2_X1 i_0_161 (.A(in3[51]), .B(in1[63]), .ZN(n_0_94));
   XNOR2_X1 i_0_162 (.A(n_0_96), .B(n_0_95), .ZN(sum[52]));
   XNOR2_X1 i_0_163 (.A(n_0_97), .B(n_0_95), .ZN(sum[53]));
   XNOR2_X1 i_0_164 (.A(n_0_98), .B(n_0_95), .ZN(sum[63]));
   XOR2_X1 i_0_165 (.A(in2[63]), .B(in1[63]), .Z(n_0_95));
   INV_X1 i_0_166 (.A(in3[52]), .ZN(n_0_96));
   INV_X1 i_0_167 (.A(in3[53]), .ZN(n_0_97));
   INV_X1 i_0_168 (.A(in3[63]), .ZN(n_0_98));
endmodule

module CSA__0_74(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;

   AND2_X1 i_0_0 (.A1(in2[19]), .A2(in1[19]), .ZN(c[20]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[21]));
   OAI21_X1 i_0_2 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[22]));
   OAI21_X1 i_0_5 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[23]));
   OAI21_X1 i_0_8 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[24]));
   OAI21_X1 i_0_11 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[25]));
   OAI21_X1 i_0_14 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[26]));
   OAI21_X1 i_0_17 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[27]));
   OAI21_X1 i_0_20 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[28]));
   OAI21_X1 i_0_23 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[29]));
   OAI21_X1 i_0_26 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[30]));
   OAI21_X1 i_0_29 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[31]));
   OAI21_X1 i_0_32 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[32]));
   OAI21_X1 i_0_35 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[33]));
   OAI21_X1 i_0_38 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[34]));
   OAI21_X1 i_0_41 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[35]));
   OAI21_X1 i_0_44 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[36]));
   OAI21_X1 i_0_47 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[37]));
   OAI21_X1 i_0_50 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[38]));
   OAI21_X1 i_0_53 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[39]));
   OAI21_X1 i_0_56 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[40]));
   OAI21_X1 i_0_59 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[41]));
   OAI21_X1 i_0_62 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[42]));
   OAI21_X1 i_0_65 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[43]));
   OAI21_X1 i_0_68 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[44]));
   OAI21_X1 i_0_71 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[45]));
   OAI21_X1 i_0_74 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[46]));
   OAI21_X1 i_0_77 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[47]));
   OAI21_X1 i_0_80 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[48]));
   OAI21_X1 i_0_83 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[49]));
   OAI21_X1 i_0_86 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[50]));
   OAI21_X1 i_0_89 (.A(in2[49]), .B1(in3[49]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[49]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_62), .A2(n_0_60), .ZN(c[51]));
   OAI21_X1 i_0_92 (.A(in3[50]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(c[63]));
   OAI21_X1 i_0_94 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   XOR2_X1 i_0_96 (.A(in2[19]), .B(in1[19]), .Z(sum[19]));
   XNOR2_X1 i_0_97 (.A(in2[20]), .B(n_0_63), .ZN(sum[20]));
   XNOR2_X1 i_0_98 (.A(in3[20]), .B(in1[20]), .ZN(n_0_63));
   XNOR2_X1 i_0_99 (.A(in2[21]), .B(n_0_64), .ZN(sum[21]));
   XNOR2_X1 i_0_100 (.A(in3[21]), .B(in1[21]), .ZN(n_0_64));
   XNOR2_X1 i_0_101 (.A(in2[22]), .B(n_0_65), .ZN(sum[22]));
   XNOR2_X1 i_0_102 (.A(in3[22]), .B(in1[22]), .ZN(n_0_65));
   XNOR2_X1 i_0_103 (.A(in2[23]), .B(n_0_66), .ZN(sum[23]));
   XNOR2_X1 i_0_104 (.A(in3[23]), .B(in1[23]), .ZN(n_0_66));
   XNOR2_X1 i_0_105 (.A(in2[24]), .B(n_0_67), .ZN(sum[24]));
   XNOR2_X1 i_0_106 (.A(in3[24]), .B(in1[24]), .ZN(n_0_67));
   XNOR2_X1 i_0_107 (.A(in2[25]), .B(n_0_68), .ZN(sum[25]));
   XNOR2_X1 i_0_108 (.A(in3[25]), .B(in1[25]), .ZN(n_0_68));
   XNOR2_X1 i_0_109 (.A(in2[26]), .B(n_0_69), .ZN(sum[26]));
   XNOR2_X1 i_0_110 (.A(in3[26]), .B(in1[26]), .ZN(n_0_69));
   XNOR2_X1 i_0_111 (.A(in2[27]), .B(n_0_70), .ZN(sum[27]));
   XNOR2_X1 i_0_112 (.A(in3[27]), .B(in1[27]), .ZN(n_0_70));
   XNOR2_X1 i_0_113 (.A(in2[28]), .B(n_0_71), .ZN(sum[28]));
   XNOR2_X1 i_0_114 (.A(in3[28]), .B(in1[28]), .ZN(n_0_71));
   XNOR2_X1 i_0_115 (.A(in2[29]), .B(n_0_72), .ZN(sum[29]));
   XNOR2_X1 i_0_116 (.A(in3[29]), .B(in1[29]), .ZN(n_0_72));
   XNOR2_X1 i_0_117 (.A(in2[30]), .B(n_0_73), .ZN(sum[30]));
   XNOR2_X1 i_0_118 (.A(in3[30]), .B(in1[30]), .ZN(n_0_73));
   XNOR2_X1 i_0_119 (.A(in2[31]), .B(n_0_74), .ZN(sum[31]));
   XNOR2_X1 i_0_120 (.A(in3[31]), .B(in1[31]), .ZN(n_0_74));
   XNOR2_X1 i_0_121 (.A(in2[32]), .B(n_0_75), .ZN(sum[32]));
   XNOR2_X1 i_0_122 (.A(in3[32]), .B(in1[32]), .ZN(n_0_75));
   XNOR2_X1 i_0_123 (.A(in2[33]), .B(n_0_76), .ZN(sum[33]));
   XNOR2_X1 i_0_124 (.A(in3[33]), .B(in1[33]), .ZN(n_0_76));
   XNOR2_X1 i_0_125 (.A(in2[34]), .B(n_0_77), .ZN(sum[34]));
   XNOR2_X1 i_0_126 (.A(in3[34]), .B(in1[34]), .ZN(n_0_77));
   XNOR2_X1 i_0_127 (.A(in2[35]), .B(n_0_78), .ZN(sum[35]));
   XNOR2_X1 i_0_128 (.A(in3[35]), .B(in1[35]), .ZN(n_0_78));
   XNOR2_X1 i_0_129 (.A(in2[36]), .B(n_0_79), .ZN(sum[36]));
   XNOR2_X1 i_0_130 (.A(in3[36]), .B(in1[36]), .ZN(n_0_79));
   XNOR2_X1 i_0_131 (.A(in2[37]), .B(n_0_80), .ZN(sum[37]));
   XNOR2_X1 i_0_132 (.A(in3[37]), .B(in1[37]), .ZN(n_0_80));
   XNOR2_X1 i_0_133 (.A(in2[38]), .B(n_0_81), .ZN(sum[38]));
   XNOR2_X1 i_0_134 (.A(in3[38]), .B(in1[38]), .ZN(n_0_81));
   XNOR2_X1 i_0_135 (.A(in2[39]), .B(n_0_82), .ZN(sum[39]));
   XNOR2_X1 i_0_136 (.A(in3[39]), .B(in1[39]), .ZN(n_0_82));
   XNOR2_X1 i_0_137 (.A(in2[40]), .B(n_0_83), .ZN(sum[40]));
   XNOR2_X1 i_0_138 (.A(in3[40]), .B(in1[40]), .ZN(n_0_83));
   XNOR2_X1 i_0_139 (.A(in2[41]), .B(n_0_84), .ZN(sum[41]));
   XNOR2_X1 i_0_140 (.A(in3[41]), .B(in1[41]), .ZN(n_0_84));
   XNOR2_X1 i_0_141 (.A(in2[42]), .B(n_0_85), .ZN(sum[42]));
   XNOR2_X1 i_0_142 (.A(in3[42]), .B(in1[42]), .ZN(n_0_85));
   XNOR2_X1 i_0_143 (.A(in2[43]), .B(n_0_86), .ZN(sum[43]));
   XNOR2_X1 i_0_144 (.A(in3[43]), .B(in1[43]), .ZN(n_0_86));
   XNOR2_X1 i_0_145 (.A(in2[44]), .B(n_0_87), .ZN(sum[44]));
   XNOR2_X1 i_0_146 (.A(in3[44]), .B(in1[44]), .ZN(n_0_87));
   XNOR2_X1 i_0_147 (.A(in2[45]), .B(n_0_88), .ZN(sum[45]));
   XNOR2_X1 i_0_148 (.A(in3[45]), .B(in1[45]), .ZN(n_0_88));
   XNOR2_X1 i_0_149 (.A(in2[46]), .B(n_0_89), .ZN(sum[46]));
   XNOR2_X1 i_0_150 (.A(in3[46]), .B(in1[46]), .ZN(n_0_89));
   XNOR2_X1 i_0_151 (.A(in2[47]), .B(n_0_90), .ZN(sum[47]));
   XNOR2_X1 i_0_152 (.A(in3[47]), .B(in1[47]), .ZN(n_0_90));
   XNOR2_X1 i_0_153 (.A(in2[48]), .B(n_0_91), .ZN(sum[48]));
   XNOR2_X1 i_0_154 (.A(in3[48]), .B(in1[48]), .ZN(n_0_91));
   XNOR2_X1 i_0_155 (.A(in2[49]), .B(n_0_92), .ZN(sum[49]));
   XNOR2_X1 i_0_156 (.A(in3[49]), .B(in1[63]), .ZN(n_0_92));
   XOR2_X1 i_0_157 (.A(in3[50]), .B(n_0_93), .Z(sum[50]));
   XOR2_X1 i_0_158 (.A(in3[63]), .B(n_0_93), .Z(sum[63]));
   XOR2_X1 i_0_159 (.A(in2[63]), .B(in1[63]), .Z(n_0_93));
endmodule

module CSA__4_2(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;

   AND2_X1 i_0_0 (.A1(in2[29]), .A2(in1[29]), .ZN(c[30]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[31]));
   OAI21_X1 i_0_2 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[32]));
   OAI21_X1 i_0_5 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[33]));
   OAI21_X1 i_0_8 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[34]));
   OAI21_X1 i_0_11 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[35]));
   OAI21_X1 i_0_14 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[36]));
   OAI21_X1 i_0_17 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[37]));
   OAI21_X1 i_0_20 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[38]));
   OAI21_X1 i_0_23 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[39]));
   OAI21_X1 i_0_26 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[40]));
   OAI21_X1 i_0_29 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[41]));
   OAI21_X1 i_0_32 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[42]));
   OAI21_X1 i_0_35 (.A(in1[41]), .B1(in3[41]), .B2(in2[41]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in2[41]), .A2(in3[41]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[43]));
   OAI21_X1 i_0_38 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[44]));
   OAI21_X1 i_0_41 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[45]));
   OAI21_X1 i_0_44 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[46]));
   OAI21_X1 i_0_47 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[47]));
   OAI21_X1 i_0_50 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[48]));
   OAI21_X1 i_0_53 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[49]));
   OAI21_X1 i_0_56 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[50]));
   OAI21_X1 i_0_59 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[51]));
   OAI21_X1 i_0_62 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[52]));
   OAI21_X1 i_0_65 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[53]));
   OAI21_X1 i_0_68 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[54]));
   OAI21_X1 i_0_71 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[55]));
   OAI21_X1 i_0_74 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[56]));
   OAI21_X1 i_0_77 (.A(in2[55]), .B1(in3[55]), .B2(in1[55]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[55]), .A2(in1[55]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[57]));
   OAI21_X1 i_0_80 (.A(in2[56]), .B1(in3[56]), .B2(in1[56]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[56]), .A2(in1[56]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[58]));
   OAI21_X1 i_0_83 (.A(in2[57]), .B1(in3[57]), .B2(in1[57]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[57]), .A2(in1[57]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[59]));
   OAI21_X1 i_0_86 (.A(in2[58]), .B1(in3[58]), .B2(in1[58]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[58]), .A2(in1[58]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[60]));
   OAI21_X1 i_0_89 (.A(in2[59]), .B1(in3[59]), .B2(in1[59]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[59]), .A2(in1[59]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_61), .A2(n_0_60), .ZN(c[61]));
   OAI21_X1 i_0_92 (.A(in2[60]), .B1(in3[60]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(in3[60]), .A2(in1[63]), .ZN(n_0_61));
   NAND2_X1 i_0_94 (.A1(n_0_63), .A2(n_0_62), .ZN(c[63]));
   OAI21_X1 i_0_95 (.A(in2[63]), .B1(in3[63]), .B2(in1[63]), .ZN(n_0_62));
   NAND2_X1 i_0_96 (.A1(in3[63]), .A2(in1[63]), .ZN(n_0_63));
   XOR2_X1 i_0_97 (.A(in2[29]), .B(in1[29]), .Z(sum[29]));
   XNOR2_X1 i_0_98 (.A(in2[30]), .B(n_0_64), .ZN(sum[30]));
   XNOR2_X1 i_0_99 (.A(in3[30]), .B(in1[30]), .ZN(n_0_64));
   XNOR2_X1 i_0_100 (.A(in2[31]), .B(n_0_65), .ZN(sum[31]));
   XNOR2_X1 i_0_101 (.A(in3[31]), .B(in1[31]), .ZN(n_0_65));
   XNOR2_X1 i_0_102 (.A(in2[32]), .B(n_0_66), .ZN(sum[32]));
   XNOR2_X1 i_0_103 (.A(in3[32]), .B(in1[32]), .ZN(n_0_66));
   XNOR2_X1 i_0_104 (.A(in2[33]), .B(n_0_67), .ZN(sum[33]));
   XNOR2_X1 i_0_105 (.A(in3[33]), .B(in1[33]), .ZN(n_0_67));
   XNOR2_X1 i_0_106 (.A(in2[34]), .B(n_0_68), .ZN(sum[34]));
   XNOR2_X1 i_0_107 (.A(in3[34]), .B(in1[34]), .ZN(n_0_68));
   XNOR2_X1 i_0_108 (.A(in2[35]), .B(n_0_69), .ZN(sum[35]));
   XNOR2_X1 i_0_109 (.A(in3[35]), .B(in1[35]), .ZN(n_0_69));
   XNOR2_X1 i_0_110 (.A(in2[36]), .B(n_0_70), .ZN(sum[36]));
   XNOR2_X1 i_0_111 (.A(in3[36]), .B(in1[36]), .ZN(n_0_70));
   XNOR2_X1 i_0_112 (.A(in2[37]), .B(n_0_71), .ZN(sum[37]));
   XNOR2_X1 i_0_113 (.A(in3[37]), .B(in1[37]), .ZN(n_0_71));
   XNOR2_X1 i_0_114 (.A(in2[38]), .B(n_0_72), .ZN(sum[38]));
   XNOR2_X1 i_0_115 (.A(in3[38]), .B(in1[38]), .ZN(n_0_72));
   XNOR2_X1 i_0_116 (.A(in2[39]), .B(n_0_73), .ZN(sum[39]));
   XNOR2_X1 i_0_117 (.A(in3[39]), .B(in1[39]), .ZN(n_0_73));
   XNOR2_X1 i_0_118 (.A(in2[40]), .B(n_0_74), .ZN(sum[40]));
   XNOR2_X1 i_0_119 (.A(in3[40]), .B(in1[40]), .ZN(n_0_74));
   XNOR2_X1 i_0_120 (.A(in2[41]), .B(n_0_75), .ZN(sum[41]));
   XNOR2_X1 i_0_121 (.A(in3[41]), .B(in1[41]), .ZN(n_0_75));
   XNOR2_X1 i_0_122 (.A(in2[42]), .B(n_0_76), .ZN(sum[42]));
   XNOR2_X1 i_0_123 (.A(in3[42]), .B(in1[42]), .ZN(n_0_76));
   XNOR2_X1 i_0_124 (.A(in2[43]), .B(n_0_77), .ZN(sum[43]));
   XNOR2_X1 i_0_125 (.A(in3[43]), .B(in1[43]), .ZN(n_0_77));
   XNOR2_X1 i_0_126 (.A(in2[44]), .B(n_0_78), .ZN(sum[44]));
   XNOR2_X1 i_0_127 (.A(in3[44]), .B(in1[44]), .ZN(n_0_78));
   XNOR2_X1 i_0_128 (.A(in2[45]), .B(n_0_79), .ZN(sum[45]));
   XNOR2_X1 i_0_129 (.A(in3[45]), .B(in1[45]), .ZN(n_0_79));
   XNOR2_X1 i_0_130 (.A(in2[46]), .B(n_0_80), .ZN(sum[46]));
   XNOR2_X1 i_0_131 (.A(in3[46]), .B(in1[46]), .ZN(n_0_80));
   XNOR2_X1 i_0_132 (.A(in2[47]), .B(n_0_81), .ZN(sum[47]));
   XNOR2_X1 i_0_133 (.A(in3[47]), .B(in1[47]), .ZN(n_0_81));
   XNOR2_X1 i_0_134 (.A(in2[48]), .B(n_0_82), .ZN(sum[48]));
   XNOR2_X1 i_0_135 (.A(in3[48]), .B(in1[48]), .ZN(n_0_82));
   XNOR2_X1 i_0_136 (.A(in2[49]), .B(n_0_83), .ZN(sum[49]));
   XNOR2_X1 i_0_137 (.A(in3[49]), .B(in1[49]), .ZN(n_0_83));
   XNOR2_X1 i_0_138 (.A(in2[50]), .B(n_0_84), .ZN(sum[50]));
   XNOR2_X1 i_0_139 (.A(in3[50]), .B(in1[50]), .ZN(n_0_84));
   XNOR2_X1 i_0_140 (.A(in2[51]), .B(n_0_85), .ZN(sum[51]));
   XNOR2_X1 i_0_141 (.A(in3[51]), .B(in1[51]), .ZN(n_0_85));
   XNOR2_X1 i_0_142 (.A(in2[52]), .B(n_0_86), .ZN(sum[52]));
   XNOR2_X1 i_0_143 (.A(in3[52]), .B(in1[52]), .ZN(n_0_86));
   XNOR2_X1 i_0_144 (.A(in2[53]), .B(n_0_87), .ZN(sum[53]));
   XNOR2_X1 i_0_145 (.A(in3[53]), .B(in1[53]), .ZN(n_0_87));
   XNOR2_X1 i_0_146 (.A(in2[54]), .B(n_0_88), .ZN(sum[54]));
   XNOR2_X1 i_0_147 (.A(in3[54]), .B(in1[54]), .ZN(n_0_88));
   XNOR2_X1 i_0_148 (.A(in2[55]), .B(n_0_89), .ZN(sum[55]));
   XNOR2_X1 i_0_149 (.A(in3[55]), .B(in1[55]), .ZN(n_0_89));
   XNOR2_X1 i_0_150 (.A(in2[56]), .B(n_0_90), .ZN(sum[56]));
   XNOR2_X1 i_0_151 (.A(in3[56]), .B(in1[56]), .ZN(n_0_90));
   XNOR2_X1 i_0_152 (.A(in2[57]), .B(n_0_91), .ZN(sum[57]));
   XNOR2_X1 i_0_153 (.A(in3[57]), .B(in1[57]), .ZN(n_0_91));
   XNOR2_X1 i_0_154 (.A(in2[58]), .B(n_0_92), .ZN(sum[58]));
   XNOR2_X1 i_0_155 (.A(in3[58]), .B(in1[58]), .ZN(n_0_92));
   XNOR2_X1 i_0_156 (.A(in2[59]), .B(n_0_93), .ZN(sum[59]));
   XNOR2_X1 i_0_157 (.A(in3[59]), .B(in1[59]), .ZN(n_0_93));
   XNOR2_X1 i_0_158 (.A(in2[60]), .B(n_0_94), .ZN(sum[60]));
   XNOR2_X1 i_0_159 (.A(in3[60]), .B(in1[63]), .ZN(n_0_94));
   XNOR2_X1 i_0_160 (.A(in2[63]), .B(n_0_95), .ZN(sum[63]));
   XNOR2_X1 i_0_161 (.A(in3[63]), .B(in1[63]), .ZN(n_0_95));
endmodule

module CSA__4_5(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;

   AND2_X1 i_0_0 (.A1(in2[30]), .A2(in1[30]), .ZN(c[31]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[32]));
   OAI21_X1 i_0_2 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[33]));
   OAI21_X1 i_0_5 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[34]));
   OAI21_X1 i_0_8 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[35]));
   OAI21_X1 i_0_11 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[36]));
   OAI21_X1 i_0_14 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[37]));
   OAI21_X1 i_0_17 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[38]));
   OAI21_X1 i_0_20 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[39]));
   OAI21_X1 i_0_23 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[40]));
   OAI21_X1 i_0_26 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[41]));
   OAI21_X1 i_0_29 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[42]));
   OAI21_X1 i_0_32 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[43]));
   OAI21_X1 i_0_35 (.A(in1[42]), .B1(in3[42]), .B2(in2[42]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in2[42]), .A2(in3[42]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[44]));
   OAI21_X1 i_0_38 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[45]));
   OAI21_X1 i_0_41 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[46]));
   OAI21_X1 i_0_44 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[47]));
   OAI21_X1 i_0_47 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[48]));
   OAI21_X1 i_0_50 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[49]));
   OAI21_X1 i_0_53 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[50]));
   OAI21_X1 i_0_56 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[51]));
   OAI21_X1 i_0_59 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[52]));
   OAI21_X1 i_0_62 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[53]));
   OAI21_X1 i_0_65 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[54]));
   OAI21_X1 i_0_68 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[55]));
   OAI21_X1 i_0_71 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[56]));
   OAI21_X1 i_0_74 (.A(in2[55]), .B1(in3[55]), .B2(in1[55]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[55]), .A2(in1[55]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[57]));
   OAI21_X1 i_0_77 (.A(in2[56]), .B1(in3[56]), .B2(in1[56]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[56]), .A2(in1[56]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[58]));
   OAI21_X1 i_0_80 (.A(in2[57]), .B1(in3[57]), .B2(in1[57]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[57]), .A2(in1[57]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[59]));
   OAI21_X1 i_0_83 (.A(in2[58]), .B1(in3[58]), .B2(in1[58]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[58]), .A2(in1[58]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[60]));
   OAI21_X1 i_0_86 (.A(in2[59]), .B1(in3[59]), .B2(in1[59]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[59]), .A2(in1[59]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[61]));
   OAI21_X1 i_0_89 (.A(in2[60]), .B1(in3[60]), .B2(in1[60]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[60]), .A2(in1[60]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_61), .A2(n_0_60), .ZN(c[62]));
   OAI21_X1 i_0_92 (.A(in2[61]), .B1(in3[61]), .B2(in1[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(in3[61]), .A2(in1[63]), .ZN(n_0_61));
   NAND2_X1 i_0_94 (.A1(n_0_63), .A2(n_0_62), .ZN(c[63]));
   OAI21_X1 i_0_95 (.A(in2[63]), .B1(in3[63]), .B2(in1[63]), .ZN(n_0_62));
   NAND2_X1 i_0_96 (.A1(in3[63]), .A2(in1[63]), .ZN(n_0_63));
   XOR2_X1 i_0_97 (.A(in2[30]), .B(in1[30]), .Z(sum[30]));
   XNOR2_X1 i_0_98 (.A(in2[31]), .B(n_0_64), .ZN(sum[31]));
   XNOR2_X1 i_0_99 (.A(in3[31]), .B(in1[31]), .ZN(n_0_64));
   XNOR2_X1 i_0_100 (.A(in2[32]), .B(n_0_65), .ZN(sum[32]));
   XNOR2_X1 i_0_101 (.A(in3[32]), .B(in1[32]), .ZN(n_0_65));
   XNOR2_X1 i_0_102 (.A(in2[33]), .B(n_0_66), .ZN(sum[33]));
   XNOR2_X1 i_0_103 (.A(in3[33]), .B(in1[33]), .ZN(n_0_66));
   XNOR2_X1 i_0_104 (.A(in2[34]), .B(n_0_67), .ZN(sum[34]));
   XNOR2_X1 i_0_105 (.A(in3[34]), .B(in1[34]), .ZN(n_0_67));
   XNOR2_X1 i_0_106 (.A(in2[35]), .B(n_0_68), .ZN(sum[35]));
   XNOR2_X1 i_0_107 (.A(in3[35]), .B(in1[35]), .ZN(n_0_68));
   XNOR2_X1 i_0_108 (.A(in2[36]), .B(n_0_69), .ZN(sum[36]));
   XNOR2_X1 i_0_109 (.A(in3[36]), .B(in1[36]), .ZN(n_0_69));
   XNOR2_X1 i_0_110 (.A(in2[37]), .B(n_0_70), .ZN(sum[37]));
   XNOR2_X1 i_0_111 (.A(in3[37]), .B(in1[37]), .ZN(n_0_70));
   XNOR2_X1 i_0_112 (.A(in2[38]), .B(n_0_71), .ZN(sum[38]));
   XNOR2_X1 i_0_113 (.A(in3[38]), .B(in1[38]), .ZN(n_0_71));
   XNOR2_X1 i_0_114 (.A(in2[39]), .B(n_0_72), .ZN(sum[39]));
   XNOR2_X1 i_0_115 (.A(in3[39]), .B(in1[39]), .ZN(n_0_72));
   XNOR2_X1 i_0_116 (.A(in2[40]), .B(n_0_73), .ZN(sum[40]));
   XNOR2_X1 i_0_117 (.A(in3[40]), .B(in1[40]), .ZN(n_0_73));
   XNOR2_X1 i_0_118 (.A(in2[41]), .B(n_0_74), .ZN(sum[41]));
   XNOR2_X1 i_0_119 (.A(in3[41]), .B(in1[41]), .ZN(n_0_74));
   XNOR2_X1 i_0_120 (.A(in2[42]), .B(n_0_75), .ZN(sum[42]));
   XNOR2_X1 i_0_121 (.A(in3[42]), .B(in1[42]), .ZN(n_0_75));
   XNOR2_X1 i_0_122 (.A(in2[43]), .B(n_0_76), .ZN(sum[43]));
   XNOR2_X1 i_0_123 (.A(in3[43]), .B(in1[43]), .ZN(n_0_76));
   XNOR2_X1 i_0_124 (.A(in2[44]), .B(n_0_77), .ZN(sum[44]));
   XNOR2_X1 i_0_125 (.A(in3[44]), .B(in1[44]), .ZN(n_0_77));
   XNOR2_X1 i_0_126 (.A(in2[45]), .B(n_0_78), .ZN(sum[45]));
   XNOR2_X1 i_0_127 (.A(in3[45]), .B(in1[45]), .ZN(n_0_78));
   XNOR2_X1 i_0_128 (.A(in2[46]), .B(n_0_79), .ZN(sum[46]));
   XNOR2_X1 i_0_129 (.A(in3[46]), .B(in1[46]), .ZN(n_0_79));
   XNOR2_X1 i_0_130 (.A(in2[47]), .B(n_0_80), .ZN(sum[47]));
   XNOR2_X1 i_0_131 (.A(in3[47]), .B(in1[47]), .ZN(n_0_80));
   XNOR2_X1 i_0_132 (.A(in2[48]), .B(n_0_81), .ZN(sum[48]));
   XNOR2_X1 i_0_133 (.A(in3[48]), .B(in1[48]), .ZN(n_0_81));
   XNOR2_X1 i_0_134 (.A(in2[49]), .B(n_0_82), .ZN(sum[49]));
   XNOR2_X1 i_0_135 (.A(in3[49]), .B(in1[49]), .ZN(n_0_82));
   XNOR2_X1 i_0_136 (.A(in2[50]), .B(n_0_83), .ZN(sum[50]));
   XNOR2_X1 i_0_137 (.A(in3[50]), .B(in1[50]), .ZN(n_0_83));
   XNOR2_X1 i_0_138 (.A(in2[51]), .B(n_0_84), .ZN(sum[51]));
   XNOR2_X1 i_0_139 (.A(in3[51]), .B(in1[51]), .ZN(n_0_84));
   XNOR2_X1 i_0_140 (.A(in2[52]), .B(n_0_85), .ZN(sum[52]));
   XNOR2_X1 i_0_141 (.A(in3[52]), .B(in1[52]), .ZN(n_0_85));
   XNOR2_X1 i_0_142 (.A(in2[53]), .B(n_0_86), .ZN(sum[53]));
   XNOR2_X1 i_0_143 (.A(in3[53]), .B(in1[53]), .ZN(n_0_86));
   XNOR2_X1 i_0_144 (.A(in2[54]), .B(n_0_87), .ZN(sum[54]));
   XNOR2_X1 i_0_145 (.A(in3[54]), .B(in1[54]), .ZN(n_0_87));
   XNOR2_X1 i_0_146 (.A(in2[55]), .B(n_0_88), .ZN(sum[55]));
   XNOR2_X1 i_0_147 (.A(in3[55]), .B(in1[55]), .ZN(n_0_88));
   XNOR2_X1 i_0_148 (.A(in2[56]), .B(n_0_89), .ZN(sum[56]));
   XNOR2_X1 i_0_149 (.A(in3[56]), .B(in1[56]), .ZN(n_0_89));
   XNOR2_X1 i_0_150 (.A(in2[57]), .B(n_0_90), .ZN(sum[57]));
   XNOR2_X1 i_0_151 (.A(in3[57]), .B(in1[57]), .ZN(n_0_90));
   XNOR2_X1 i_0_152 (.A(in2[58]), .B(n_0_91), .ZN(sum[58]));
   XNOR2_X1 i_0_153 (.A(in3[58]), .B(in1[58]), .ZN(n_0_91));
   XNOR2_X1 i_0_154 (.A(in2[59]), .B(n_0_92), .ZN(sum[59]));
   XNOR2_X1 i_0_155 (.A(in3[59]), .B(in1[59]), .ZN(n_0_92));
   XNOR2_X1 i_0_156 (.A(in2[60]), .B(n_0_93), .ZN(sum[60]));
   XNOR2_X1 i_0_157 (.A(in3[60]), .B(in1[60]), .ZN(n_0_93));
   XNOR2_X1 i_0_158 (.A(in2[61]), .B(n_0_94), .ZN(sum[61]));
   XNOR2_X1 i_0_159 (.A(in3[61]), .B(in1[63]), .ZN(n_0_94));
   XNOR2_X1 i_0_160 (.A(in2[63]), .B(n_0_95), .ZN(sum[63]));
   XNOR2_X1 i_0_161 (.A(in3[63]), .B(in1[63]), .ZN(n_0_95));
endmodule

module CSA__4_8(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;

   AND2_X1 i_0_0 (.A1(in2[24]), .A2(in1[24]), .ZN(c[25]));
   AND2_X1 i_0_1 (.A1(in2[25]), .A2(in1[25]), .ZN(c[26]));
   AND2_X1 i_0_2 (.A1(in2[26]), .A2(in1[26]), .ZN(c[27]));
   NAND2_X1 i_0_3 (.A1(n_0_1), .A2(n_0_0), .ZN(c[28]));
   OAI21_X1 i_0_4 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_0));
   NAND2_X1 i_0_5 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_1));
   NAND2_X1 i_0_6 (.A1(n_0_3), .A2(n_0_2), .ZN(c[29]));
   OAI21_X1 i_0_7 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_2));
   NAND2_X1 i_0_8 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_3));
   NAND2_X1 i_0_9 (.A1(n_0_5), .A2(n_0_4), .ZN(c[30]));
   OAI21_X1 i_0_10 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_4));
   NAND2_X1 i_0_11 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_5));
   NAND2_X1 i_0_12 (.A1(n_0_7), .A2(n_0_6), .ZN(c[31]));
   OAI21_X1 i_0_13 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_6));
   NAND2_X1 i_0_14 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_7));
   NAND2_X1 i_0_15 (.A1(n_0_9), .A2(n_0_8), .ZN(c[32]));
   OAI21_X1 i_0_16 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_8));
   NAND2_X1 i_0_17 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_9));
   NAND2_X1 i_0_18 (.A1(n_0_11), .A2(n_0_10), .ZN(c[33]));
   OAI21_X1 i_0_19 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_10));
   NAND2_X1 i_0_20 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_11));
   NAND2_X1 i_0_21 (.A1(n_0_13), .A2(n_0_12), .ZN(c[34]));
   OAI21_X1 i_0_22 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_12));
   NAND2_X1 i_0_23 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_13));
   NAND2_X1 i_0_24 (.A1(n_0_15), .A2(n_0_14), .ZN(c[35]));
   OAI21_X1 i_0_25 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_14));
   NAND2_X1 i_0_26 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_15));
   NAND2_X1 i_0_27 (.A1(n_0_17), .A2(n_0_16), .ZN(c[36]));
   OAI21_X1 i_0_28 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_16));
   NAND2_X1 i_0_29 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_17));
   NAND2_X1 i_0_30 (.A1(n_0_19), .A2(n_0_18), .ZN(c[37]));
   OAI21_X1 i_0_31 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_18));
   NAND2_X1 i_0_32 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_19));
   NAND2_X1 i_0_33 (.A1(n_0_21), .A2(n_0_20), .ZN(c[38]));
   OAI21_X1 i_0_34 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_20));
   NAND2_X1 i_0_35 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_21));
   NAND2_X1 i_0_36 (.A1(n_0_23), .A2(n_0_22), .ZN(c[39]));
   OAI21_X1 i_0_37 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_22));
   NAND2_X1 i_0_38 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_23));
   NAND2_X1 i_0_39 (.A1(n_0_25), .A2(n_0_24), .ZN(c[40]));
   OAI21_X1 i_0_40 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_24));
   NAND2_X1 i_0_41 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_25));
   NAND2_X1 i_0_42 (.A1(n_0_27), .A2(n_0_26), .ZN(c[41]));
   OAI21_X1 i_0_43 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_26));
   NAND2_X1 i_0_44 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_27));
   NAND2_X1 i_0_45 (.A1(n_0_29), .A2(n_0_28), .ZN(c[42]));
   OAI21_X1 i_0_46 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_28));
   NAND2_X1 i_0_47 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_29));
   NAND2_X1 i_0_48 (.A1(n_0_31), .A2(n_0_30), .ZN(c[43]));
   OAI21_X1 i_0_49 (.A(in3[42]), .B1(in1[42]), .B2(in2[42]), .ZN(n_0_30));
   NAND2_X1 i_0_50 (.A1(in2[42]), .A2(in1[42]), .ZN(n_0_31));
   NAND2_X1 i_0_51 (.A1(n_0_33), .A2(n_0_32), .ZN(c[44]));
   OAI21_X1 i_0_52 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_32));
   NAND2_X1 i_0_53 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_33));
   NAND2_X1 i_0_54 (.A1(n_0_35), .A2(n_0_34), .ZN(c[45]));
   OAI21_X1 i_0_55 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_34));
   NAND2_X1 i_0_56 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_35));
   NAND2_X1 i_0_57 (.A1(n_0_37), .A2(n_0_36), .ZN(c[46]));
   OAI21_X1 i_0_58 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_36));
   NAND2_X1 i_0_59 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_37));
   NAND2_X1 i_0_60 (.A1(n_0_39), .A2(n_0_38), .ZN(c[47]));
   OAI21_X1 i_0_61 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_38));
   NAND2_X1 i_0_62 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_39));
   NAND2_X1 i_0_63 (.A1(n_0_41), .A2(n_0_40), .ZN(c[48]));
   OAI21_X1 i_0_64 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_40));
   NAND2_X1 i_0_65 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_41));
   NAND2_X1 i_0_66 (.A1(n_0_43), .A2(n_0_42), .ZN(c[49]));
   OAI21_X1 i_0_67 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_42));
   NAND2_X1 i_0_68 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_43));
   NAND2_X1 i_0_69 (.A1(n_0_45), .A2(n_0_44), .ZN(c[50]));
   OAI21_X1 i_0_70 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_44));
   NAND2_X1 i_0_71 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_45));
   NAND2_X1 i_0_72 (.A1(n_0_47), .A2(n_0_46), .ZN(c[51]));
   OAI21_X1 i_0_73 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_46));
   NAND2_X1 i_0_74 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_47));
   NAND2_X1 i_0_75 (.A1(n_0_49), .A2(n_0_48), .ZN(c[52]));
   OAI21_X1 i_0_76 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_48));
   NAND2_X1 i_0_77 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_49));
   NAND2_X1 i_0_78 (.A1(n_0_51), .A2(n_0_50), .ZN(c[53]));
   OAI21_X1 i_0_79 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_50));
   NAND2_X1 i_0_80 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_51));
   NAND2_X1 i_0_81 (.A1(n_0_53), .A2(n_0_52), .ZN(c[54]));
   OAI21_X1 i_0_82 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_52));
   NAND2_X1 i_0_83 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_53));
   NAND2_X1 i_0_84 (.A1(n_0_55), .A2(n_0_54), .ZN(c[55]));
   OAI21_X1 i_0_85 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_54));
   NAND2_X1 i_0_86 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_55));
   NAND2_X1 i_0_87 (.A1(n_0_57), .A2(n_0_56), .ZN(c[56]));
   OAI21_X1 i_0_88 (.A(in2[55]), .B1(in3[55]), .B2(in1[55]), .ZN(n_0_56));
   NAND2_X1 i_0_89 (.A1(in3[55]), .A2(in1[55]), .ZN(n_0_57));
   NAND2_X1 i_0_90 (.A1(n_0_59), .A2(n_0_58), .ZN(c[57]));
   OAI21_X1 i_0_91 (.A(in2[56]), .B1(in3[56]), .B2(in1[56]), .ZN(n_0_58));
   NAND2_X1 i_0_92 (.A1(in3[56]), .A2(in1[56]), .ZN(n_0_59));
   NAND2_X1 i_0_93 (.A1(n_0_61), .A2(n_0_60), .ZN(c[58]));
   OAI21_X1 i_0_94 (.A(in2[57]), .B1(in3[57]), .B2(in1[57]), .ZN(n_0_60));
   NAND2_X1 i_0_95 (.A1(in3[57]), .A2(in1[57]), .ZN(n_0_61));
   NAND2_X1 i_0_96 (.A1(n_0_63), .A2(n_0_62), .ZN(c[59]));
   OAI21_X1 i_0_97 (.A(in2[58]), .B1(in3[58]), .B2(in1[58]), .ZN(n_0_62));
   NAND2_X1 i_0_98 (.A1(in3[58]), .A2(in1[58]), .ZN(n_0_63));
   NAND2_X1 i_0_99 (.A1(n_0_65), .A2(n_0_64), .ZN(c[60]));
   OAI21_X1 i_0_100 (.A(in2[59]), .B1(in3[59]), .B2(in1[63]), .ZN(n_0_64));
   NAND2_X1 i_0_101 (.A1(in3[59]), .A2(in1[63]), .ZN(n_0_65));
   AOI21_X1 i_0_102 (.A(n_0_67), .B1(n_0_66), .B2(n_0_102), .ZN(c[61]));
   AOI21_X1 i_0_103 (.A(n_0_67), .B1(n_0_66), .B2(n_0_103), .ZN(c[62]));
   AOI21_X1 i_0_104 (.A(n_0_67), .B1(n_0_66), .B2(n_0_104), .ZN(c[63]));
   NAND2_X1 i_0_105 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_66));
   NOR2_X1 i_0_106 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_67));
   XOR2_X1 i_0_107 (.A(in2[24]), .B(in1[24]), .Z(sum[24]));
   XOR2_X1 i_0_108 (.A(in2[25]), .B(in1[25]), .Z(sum[25]));
   XOR2_X1 i_0_109 (.A(in2[26]), .B(in1[26]), .Z(sum[26]));
   XNOR2_X1 i_0_110 (.A(in2[27]), .B(n_0_68), .ZN(sum[27]));
   XNOR2_X1 i_0_111 (.A(in3[27]), .B(in1[27]), .ZN(n_0_68));
   XNOR2_X1 i_0_112 (.A(in2[28]), .B(n_0_69), .ZN(sum[28]));
   XNOR2_X1 i_0_113 (.A(in3[28]), .B(in1[28]), .ZN(n_0_69));
   XNOR2_X1 i_0_114 (.A(in2[29]), .B(n_0_70), .ZN(sum[29]));
   XNOR2_X1 i_0_115 (.A(in3[29]), .B(in1[29]), .ZN(n_0_70));
   XNOR2_X1 i_0_116 (.A(in2[30]), .B(n_0_71), .ZN(sum[30]));
   XNOR2_X1 i_0_117 (.A(in3[30]), .B(in1[30]), .ZN(n_0_71));
   XNOR2_X1 i_0_118 (.A(in2[31]), .B(n_0_72), .ZN(sum[31]));
   XNOR2_X1 i_0_119 (.A(in3[31]), .B(in1[31]), .ZN(n_0_72));
   XNOR2_X1 i_0_120 (.A(in2[32]), .B(n_0_73), .ZN(sum[32]));
   XNOR2_X1 i_0_121 (.A(in3[32]), .B(in1[32]), .ZN(n_0_73));
   XNOR2_X1 i_0_122 (.A(in2[33]), .B(n_0_74), .ZN(sum[33]));
   XNOR2_X1 i_0_123 (.A(in3[33]), .B(in1[33]), .ZN(n_0_74));
   XNOR2_X1 i_0_124 (.A(in2[34]), .B(n_0_75), .ZN(sum[34]));
   XNOR2_X1 i_0_125 (.A(in3[34]), .B(in1[34]), .ZN(n_0_75));
   XNOR2_X1 i_0_126 (.A(in2[35]), .B(n_0_76), .ZN(sum[35]));
   XNOR2_X1 i_0_127 (.A(in3[35]), .B(in1[35]), .ZN(n_0_76));
   XNOR2_X1 i_0_128 (.A(in2[36]), .B(n_0_77), .ZN(sum[36]));
   XNOR2_X1 i_0_129 (.A(in3[36]), .B(in1[36]), .ZN(n_0_77));
   XNOR2_X1 i_0_130 (.A(in2[37]), .B(n_0_78), .ZN(sum[37]));
   XNOR2_X1 i_0_131 (.A(in3[37]), .B(in1[37]), .ZN(n_0_78));
   XNOR2_X1 i_0_132 (.A(in2[38]), .B(n_0_79), .ZN(sum[38]));
   XNOR2_X1 i_0_133 (.A(in3[38]), .B(in1[38]), .ZN(n_0_79));
   XNOR2_X1 i_0_134 (.A(in2[39]), .B(n_0_80), .ZN(sum[39]));
   XNOR2_X1 i_0_135 (.A(in3[39]), .B(in1[39]), .ZN(n_0_80));
   XNOR2_X1 i_0_136 (.A(in2[40]), .B(n_0_81), .ZN(sum[40]));
   XNOR2_X1 i_0_137 (.A(in3[40]), .B(in1[40]), .ZN(n_0_81));
   XNOR2_X1 i_0_138 (.A(in2[41]), .B(n_0_82), .ZN(sum[41]));
   XNOR2_X1 i_0_139 (.A(in3[41]), .B(in1[41]), .ZN(n_0_82));
   XNOR2_X1 i_0_140 (.A(in2[42]), .B(n_0_83), .ZN(sum[42]));
   XNOR2_X1 i_0_141 (.A(in3[42]), .B(in1[42]), .ZN(n_0_83));
   XNOR2_X1 i_0_142 (.A(in2[43]), .B(n_0_84), .ZN(sum[43]));
   XNOR2_X1 i_0_143 (.A(in3[43]), .B(in1[43]), .ZN(n_0_84));
   XNOR2_X1 i_0_144 (.A(in2[44]), .B(n_0_85), .ZN(sum[44]));
   XNOR2_X1 i_0_145 (.A(in3[44]), .B(in1[44]), .ZN(n_0_85));
   XNOR2_X1 i_0_146 (.A(in2[45]), .B(n_0_86), .ZN(sum[45]));
   XNOR2_X1 i_0_147 (.A(in3[45]), .B(in1[45]), .ZN(n_0_86));
   XNOR2_X1 i_0_148 (.A(in2[46]), .B(n_0_87), .ZN(sum[46]));
   XNOR2_X1 i_0_149 (.A(in3[46]), .B(in1[46]), .ZN(n_0_87));
   XNOR2_X1 i_0_150 (.A(in2[47]), .B(n_0_88), .ZN(sum[47]));
   XNOR2_X1 i_0_151 (.A(in3[47]), .B(in1[47]), .ZN(n_0_88));
   XNOR2_X1 i_0_152 (.A(in2[48]), .B(n_0_89), .ZN(sum[48]));
   XNOR2_X1 i_0_153 (.A(in3[48]), .B(in1[48]), .ZN(n_0_89));
   XNOR2_X1 i_0_154 (.A(in2[49]), .B(n_0_90), .ZN(sum[49]));
   XNOR2_X1 i_0_155 (.A(in3[49]), .B(in1[49]), .ZN(n_0_90));
   XNOR2_X1 i_0_156 (.A(in2[50]), .B(n_0_91), .ZN(sum[50]));
   XNOR2_X1 i_0_157 (.A(in3[50]), .B(in1[50]), .ZN(n_0_91));
   XNOR2_X1 i_0_158 (.A(in2[51]), .B(n_0_92), .ZN(sum[51]));
   XNOR2_X1 i_0_159 (.A(in3[51]), .B(in1[51]), .ZN(n_0_92));
   XNOR2_X1 i_0_160 (.A(in2[52]), .B(n_0_93), .ZN(sum[52]));
   XNOR2_X1 i_0_161 (.A(in3[52]), .B(in1[52]), .ZN(n_0_93));
   XNOR2_X1 i_0_162 (.A(in2[53]), .B(n_0_94), .ZN(sum[53]));
   XNOR2_X1 i_0_163 (.A(in3[53]), .B(in1[53]), .ZN(n_0_94));
   XNOR2_X1 i_0_164 (.A(in2[54]), .B(n_0_95), .ZN(sum[54]));
   XNOR2_X1 i_0_165 (.A(in3[54]), .B(in1[54]), .ZN(n_0_95));
   XNOR2_X1 i_0_166 (.A(in2[55]), .B(n_0_96), .ZN(sum[55]));
   XNOR2_X1 i_0_167 (.A(in3[55]), .B(in1[55]), .ZN(n_0_96));
   XNOR2_X1 i_0_168 (.A(in2[56]), .B(n_0_97), .ZN(sum[56]));
   XNOR2_X1 i_0_169 (.A(in3[56]), .B(in1[56]), .ZN(n_0_97));
   XNOR2_X1 i_0_170 (.A(in2[57]), .B(n_0_98), .ZN(sum[57]));
   XNOR2_X1 i_0_171 (.A(in3[57]), .B(in1[57]), .ZN(n_0_98));
   XNOR2_X1 i_0_172 (.A(in2[58]), .B(n_0_99), .ZN(sum[58]));
   XNOR2_X1 i_0_173 (.A(in3[58]), .B(in1[58]), .ZN(n_0_99));
   XNOR2_X1 i_0_174 (.A(in2[59]), .B(n_0_100), .ZN(sum[59]));
   XNOR2_X1 i_0_175 (.A(in3[59]), .B(in1[63]), .ZN(n_0_100));
   XNOR2_X1 i_0_176 (.A(n_0_102), .B(n_0_101), .ZN(sum[60]));
   XNOR2_X1 i_0_177 (.A(n_0_103), .B(n_0_101), .ZN(sum[61]));
   XNOR2_X1 i_0_178 (.A(n_0_104), .B(n_0_101), .ZN(sum[63]));
   XOR2_X1 i_0_179 (.A(in2[63]), .B(in1[63]), .Z(n_0_101));
   INV_X1 i_0_180 (.A(in3[60]), .ZN(n_0_102));
   INV_X1 i_0_181 (.A(in3[61]), .ZN(n_0_103));
   INV_X1 i_0_182 (.A(in3[63]), .ZN(n_0_104));
endmodule

module CSA__4_11(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;

   AND2_X1 i_0_0 (.A1(in2[21]), .A2(in1[21]), .ZN(c[22]));
   AND2_X1 i_0_1 (.A1(in2[22]), .A2(in1[22]), .ZN(c[23]));
   AND2_X1 i_0_2 (.A1(in2[23]), .A2(in1[23]), .ZN(c[24]));
   AND2_X1 i_0_3 (.A1(in2[24]), .A2(in1[24]), .ZN(c[25]));
   NAND2_X1 i_0_4 (.A1(n_0_1), .A2(n_0_0), .ZN(c[26]));
   OAI21_X1 i_0_5 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_1));
   NAND2_X1 i_0_7 (.A1(n_0_3), .A2(n_0_2), .ZN(c[27]));
   OAI21_X1 i_0_8 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_2));
   NAND2_X1 i_0_9 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_3));
   NAND2_X1 i_0_10 (.A1(n_0_5), .A2(n_0_4), .ZN(c[28]));
   OAI21_X1 i_0_11 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_4));
   NAND2_X1 i_0_12 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_5));
   NAND2_X1 i_0_13 (.A1(n_0_7), .A2(n_0_6), .ZN(c[29]));
   OAI21_X1 i_0_14 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_6));
   NAND2_X1 i_0_15 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_7));
   NAND2_X1 i_0_16 (.A1(n_0_9), .A2(n_0_8), .ZN(c[30]));
   OAI21_X1 i_0_17 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_8));
   NAND2_X1 i_0_18 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_9));
   NAND2_X1 i_0_19 (.A1(n_0_11), .A2(n_0_10), .ZN(c[31]));
   OAI21_X1 i_0_20 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_10));
   NAND2_X1 i_0_21 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_11));
   NAND2_X1 i_0_22 (.A1(n_0_13), .A2(n_0_12), .ZN(c[32]));
   OAI21_X1 i_0_23 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_12));
   NAND2_X1 i_0_24 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_13));
   NAND2_X1 i_0_25 (.A1(n_0_15), .A2(n_0_14), .ZN(c[33]));
   OAI21_X1 i_0_26 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_14));
   NAND2_X1 i_0_27 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_15));
   NAND2_X1 i_0_28 (.A1(n_0_17), .A2(n_0_16), .ZN(c[34]));
   OAI21_X1 i_0_29 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_16));
   NAND2_X1 i_0_30 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_17));
   NAND2_X1 i_0_31 (.A1(n_0_19), .A2(n_0_18), .ZN(c[35]));
   OAI21_X1 i_0_32 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_18));
   NAND2_X1 i_0_33 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_19));
   NAND2_X1 i_0_34 (.A1(n_0_21), .A2(n_0_20), .ZN(c[36]));
   OAI21_X1 i_0_35 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_20));
   NAND2_X1 i_0_36 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_21));
   NAND2_X1 i_0_37 (.A1(n_0_23), .A2(n_0_22), .ZN(c[37]));
   OAI21_X1 i_0_38 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_22));
   NAND2_X1 i_0_39 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_23));
   NAND2_X1 i_0_40 (.A1(n_0_25), .A2(n_0_24), .ZN(c[38]));
   OAI21_X1 i_0_41 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_24));
   NAND2_X1 i_0_42 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_25));
   NAND2_X1 i_0_43 (.A1(n_0_27), .A2(n_0_26), .ZN(c[39]));
   OAI21_X1 i_0_44 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_26));
   NAND2_X1 i_0_45 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_27));
   NAND2_X1 i_0_46 (.A1(n_0_29), .A2(n_0_28), .ZN(c[40]));
   OAI21_X1 i_0_47 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_28));
   NAND2_X1 i_0_48 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_29));
   NAND2_X1 i_0_49 (.A1(n_0_31), .A2(n_0_30), .ZN(c[41]));
   OAI21_X1 i_0_50 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_30));
   NAND2_X1 i_0_51 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_31));
   NAND2_X1 i_0_52 (.A1(n_0_33), .A2(n_0_32), .ZN(c[42]));
   OAI21_X1 i_0_53 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_32));
   NAND2_X1 i_0_54 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_33));
   NAND2_X1 i_0_55 (.A1(n_0_35), .A2(n_0_34), .ZN(c[43]));
   OAI21_X1 i_0_56 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_34));
   NAND2_X1 i_0_57 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_35));
   NAND2_X1 i_0_58 (.A1(n_0_37), .A2(n_0_36), .ZN(c[44]));
   OAI21_X1 i_0_59 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_36));
   NAND2_X1 i_0_60 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_37));
   NAND2_X1 i_0_61 (.A1(n_0_39), .A2(n_0_38), .ZN(c[45]));
   OAI21_X1 i_0_62 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_38));
   NAND2_X1 i_0_63 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_39));
   NAND2_X1 i_0_64 (.A1(n_0_41), .A2(n_0_40), .ZN(c[46]));
   OAI21_X1 i_0_65 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_40));
   NAND2_X1 i_0_66 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_41));
   NAND2_X1 i_0_67 (.A1(n_0_43), .A2(n_0_42), .ZN(c[47]));
   OAI21_X1 i_0_68 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_42));
   NAND2_X1 i_0_69 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_43));
   NAND2_X1 i_0_70 (.A1(n_0_45), .A2(n_0_44), .ZN(c[48]));
   OAI21_X1 i_0_71 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_44));
   NAND2_X1 i_0_72 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_45));
   NAND2_X1 i_0_73 (.A1(n_0_47), .A2(n_0_46), .ZN(c[49]));
   OAI21_X1 i_0_74 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_46));
   NAND2_X1 i_0_75 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_47));
   NAND2_X1 i_0_76 (.A1(n_0_49), .A2(n_0_48), .ZN(c[50]));
   OAI21_X1 i_0_77 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_48));
   NAND2_X1 i_0_78 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_49));
   NAND2_X1 i_0_79 (.A1(n_0_51), .A2(n_0_50), .ZN(c[51]));
   OAI21_X1 i_0_80 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_50));
   NAND2_X1 i_0_81 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_51));
   NAND2_X1 i_0_82 (.A1(n_0_53), .A2(n_0_52), .ZN(c[52]));
   OAI21_X1 i_0_83 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_52));
   NAND2_X1 i_0_84 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_53));
   NAND2_X1 i_0_85 (.A1(n_0_55), .A2(n_0_54), .ZN(c[53]));
   OAI21_X1 i_0_86 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_54));
   NAND2_X1 i_0_87 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_55));
   NAND2_X1 i_0_88 (.A1(n_0_57), .A2(n_0_56), .ZN(c[54]));
   OAI21_X1 i_0_89 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_56));
   NAND2_X1 i_0_90 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_57));
   NAND2_X1 i_0_91 (.A1(n_0_59), .A2(n_0_58), .ZN(c[55]));
   OAI21_X1 i_0_92 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_58));
   NAND2_X1 i_0_93 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_59));
   NAND2_X1 i_0_94 (.A1(n_0_61), .A2(n_0_60), .ZN(c[56]));
   OAI21_X1 i_0_95 (.A(in2[55]), .B1(in3[55]), .B2(in1[55]), .ZN(n_0_60));
   NAND2_X1 i_0_96 (.A1(in3[55]), .A2(in1[55]), .ZN(n_0_61));
   NAND2_X1 i_0_97 (.A1(n_0_63), .A2(n_0_62), .ZN(c[57]));
   OAI21_X1 i_0_98 (.A(in3[56]), .B1(in1[63]), .B2(in2[56]), .ZN(n_0_62));
   NAND2_X1 i_0_99 (.A1(in2[56]), .A2(in1[63]), .ZN(n_0_63));
   NAND2_X1 i_0_100 (.A1(n_0_65), .A2(n_0_64), .ZN(c[58]));
   OAI21_X1 i_0_101 (.A(in2[57]), .B1(in3[57]), .B2(in1[63]), .ZN(n_0_64));
   NAND2_X1 i_0_102 (.A1(in3[57]), .A2(in1[63]), .ZN(n_0_65));
   NAND2_X1 i_0_103 (.A1(n_0_67), .A2(n_0_66), .ZN(c[59]));
   OAI21_X1 i_0_104 (.A(in2[58]), .B1(in3[58]), .B2(in1[63]), .ZN(n_0_66));
   NAND2_X1 i_0_105 (.A1(in3[58]), .A2(in1[63]), .ZN(n_0_67));
   NAND2_X1 i_0_106 (.A1(n_0_69), .A2(n_0_68), .ZN(c[60]));
   OAI21_X1 i_0_107 (.A(in2[59]), .B1(in3[59]), .B2(in1[63]), .ZN(n_0_68));
   NAND2_X1 i_0_108 (.A1(in3[59]), .A2(in1[63]), .ZN(n_0_69));
   NAND2_X1 i_0_109 (.A1(n_0_71), .A2(n_0_70), .ZN(c[61]));
   OAI21_X1 i_0_110 (.A(in2[60]), .B1(in3[60]), .B2(in1[63]), .ZN(n_0_70));
   NAND2_X1 i_0_111 (.A1(in3[60]), .A2(in1[63]), .ZN(n_0_71));
   NAND2_X1 i_0_112 (.A1(n_0_73), .A2(n_0_72), .ZN(c[62]));
   OAI21_X1 i_0_113 (.A(in2[61]), .B1(in3[61]), .B2(in1[63]), .ZN(n_0_72));
   NAND2_X1 i_0_114 (.A1(in3[61]), .A2(in1[63]), .ZN(n_0_73));
   NAND2_X1 i_0_115 (.A1(n_0_75), .A2(n_0_74), .ZN(c[63]));
   OAI21_X1 i_0_116 (.A(in3[62]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_74));
   NAND2_X1 i_0_117 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_75));
   XOR2_X1 i_0_118 (.A(in2[21]), .B(in1[21]), .Z(sum[21]));
   XOR2_X1 i_0_119 (.A(in2[22]), .B(in1[22]), .Z(sum[22]));
   XOR2_X1 i_0_120 (.A(in2[23]), .B(in1[23]), .Z(sum[23]));
   XOR2_X1 i_0_121 (.A(in2[24]), .B(in1[24]), .Z(sum[24]));
   XNOR2_X1 i_0_122 (.A(in2[25]), .B(n_0_76), .ZN(sum[25]));
   XNOR2_X1 i_0_123 (.A(in3[25]), .B(in1[25]), .ZN(n_0_76));
   XNOR2_X1 i_0_124 (.A(in2[26]), .B(n_0_77), .ZN(sum[26]));
   XNOR2_X1 i_0_125 (.A(in3[26]), .B(in1[26]), .ZN(n_0_77));
   XNOR2_X1 i_0_126 (.A(in2[27]), .B(n_0_78), .ZN(sum[27]));
   XNOR2_X1 i_0_127 (.A(in3[27]), .B(in1[27]), .ZN(n_0_78));
   XNOR2_X1 i_0_128 (.A(in2[28]), .B(n_0_79), .ZN(sum[28]));
   XNOR2_X1 i_0_129 (.A(in3[28]), .B(in1[28]), .ZN(n_0_79));
   XNOR2_X1 i_0_130 (.A(in2[29]), .B(n_0_80), .ZN(sum[29]));
   XNOR2_X1 i_0_131 (.A(in3[29]), .B(in1[29]), .ZN(n_0_80));
   XNOR2_X1 i_0_132 (.A(in2[30]), .B(n_0_81), .ZN(sum[30]));
   XNOR2_X1 i_0_133 (.A(in3[30]), .B(in1[30]), .ZN(n_0_81));
   XNOR2_X1 i_0_134 (.A(in2[31]), .B(n_0_82), .ZN(sum[31]));
   XNOR2_X1 i_0_135 (.A(in3[31]), .B(in1[31]), .ZN(n_0_82));
   XNOR2_X1 i_0_136 (.A(in2[32]), .B(n_0_83), .ZN(sum[32]));
   XNOR2_X1 i_0_137 (.A(in3[32]), .B(in1[32]), .ZN(n_0_83));
   XNOR2_X1 i_0_138 (.A(in2[33]), .B(n_0_84), .ZN(sum[33]));
   XNOR2_X1 i_0_139 (.A(in3[33]), .B(in1[33]), .ZN(n_0_84));
   XNOR2_X1 i_0_140 (.A(in2[34]), .B(n_0_85), .ZN(sum[34]));
   XNOR2_X1 i_0_141 (.A(in3[34]), .B(in1[34]), .ZN(n_0_85));
   XNOR2_X1 i_0_142 (.A(in2[35]), .B(n_0_86), .ZN(sum[35]));
   XNOR2_X1 i_0_143 (.A(in3[35]), .B(in1[35]), .ZN(n_0_86));
   XNOR2_X1 i_0_144 (.A(in2[36]), .B(n_0_87), .ZN(sum[36]));
   XNOR2_X1 i_0_145 (.A(in3[36]), .B(in1[36]), .ZN(n_0_87));
   XNOR2_X1 i_0_146 (.A(in2[37]), .B(n_0_88), .ZN(sum[37]));
   XNOR2_X1 i_0_147 (.A(in3[37]), .B(in1[37]), .ZN(n_0_88));
   XNOR2_X1 i_0_148 (.A(in2[38]), .B(n_0_89), .ZN(sum[38]));
   XNOR2_X1 i_0_149 (.A(in3[38]), .B(in1[38]), .ZN(n_0_89));
   XNOR2_X1 i_0_150 (.A(in2[39]), .B(n_0_90), .ZN(sum[39]));
   XNOR2_X1 i_0_151 (.A(in3[39]), .B(in1[39]), .ZN(n_0_90));
   XNOR2_X1 i_0_152 (.A(in2[40]), .B(n_0_91), .ZN(sum[40]));
   XNOR2_X1 i_0_153 (.A(in3[40]), .B(in1[40]), .ZN(n_0_91));
   XNOR2_X1 i_0_154 (.A(in2[41]), .B(n_0_92), .ZN(sum[41]));
   XNOR2_X1 i_0_155 (.A(in3[41]), .B(in1[41]), .ZN(n_0_92));
   XNOR2_X1 i_0_156 (.A(in2[42]), .B(n_0_93), .ZN(sum[42]));
   XNOR2_X1 i_0_157 (.A(in3[42]), .B(in1[42]), .ZN(n_0_93));
   XNOR2_X1 i_0_158 (.A(in2[43]), .B(n_0_94), .ZN(sum[43]));
   XNOR2_X1 i_0_159 (.A(in3[43]), .B(in1[43]), .ZN(n_0_94));
   XNOR2_X1 i_0_160 (.A(in2[44]), .B(n_0_95), .ZN(sum[44]));
   XNOR2_X1 i_0_161 (.A(in3[44]), .B(in1[44]), .ZN(n_0_95));
   XNOR2_X1 i_0_162 (.A(in2[45]), .B(n_0_96), .ZN(sum[45]));
   XNOR2_X1 i_0_163 (.A(in3[45]), .B(in1[45]), .ZN(n_0_96));
   XNOR2_X1 i_0_164 (.A(in2[46]), .B(n_0_97), .ZN(sum[46]));
   XNOR2_X1 i_0_165 (.A(in3[46]), .B(in1[46]), .ZN(n_0_97));
   XNOR2_X1 i_0_166 (.A(in2[47]), .B(n_0_98), .ZN(sum[47]));
   XNOR2_X1 i_0_167 (.A(in3[47]), .B(in1[47]), .ZN(n_0_98));
   XNOR2_X1 i_0_168 (.A(in2[48]), .B(n_0_99), .ZN(sum[48]));
   XNOR2_X1 i_0_169 (.A(in3[48]), .B(in1[48]), .ZN(n_0_99));
   XNOR2_X1 i_0_170 (.A(in2[49]), .B(n_0_100), .ZN(sum[49]));
   XNOR2_X1 i_0_171 (.A(in3[49]), .B(in1[49]), .ZN(n_0_100));
   XNOR2_X1 i_0_172 (.A(in2[50]), .B(n_0_101), .ZN(sum[50]));
   XNOR2_X1 i_0_173 (.A(in3[50]), .B(in1[50]), .ZN(n_0_101));
   XNOR2_X1 i_0_174 (.A(in2[51]), .B(n_0_102), .ZN(sum[51]));
   XNOR2_X1 i_0_175 (.A(in3[51]), .B(in1[51]), .ZN(n_0_102));
   XNOR2_X1 i_0_176 (.A(in2[52]), .B(n_0_103), .ZN(sum[52]));
   XNOR2_X1 i_0_177 (.A(in3[52]), .B(in1[52]), .ZN(n_0_103));
   XNOR2_X1 i_0_178 (.A(in2[53]), .B(n_0_104), .ZN(sum[53]));
   XNOR2_X1 i_0_179 (.A(in3[53]), .B(in1[53]), .ZN(n_0_104));
   XNOR2_X1 i_0_180 (.A(in2[54]), .B(n_0_105), .ZN(sum[54]));
   XNOR2_X1 i_0_181 (.A(in3[54]), .B(in1[54]), .ZN(n_0_105));
   XNOR2_X1 i_0_182 (.A(in2[55]), .B(n_0_106), .ZN(sum[55]));
   XNOR2_X1 i_0_183 (.A(in3[55]), .B(in1[55]), .ZN(n_0_106));
   XNOR2_X1 i_0_184 (.A(in2[56]), .B(n_0_107), .ZN(sum[56]));
   XNOR2_X1 i_0_185 (.A(in3[56]), .B(in1[63]), .ZN(n_0_107));
   XNOR2_X1 i_0_186 (.A(in2[57]), .B(n_0_108), .ZN(sum[57]));
   XNOR2_X1 i_0_187 (.A(in3[57]), .B(in1[63]), .ZN(n_0_108));
   XNOR2_X1 i_0_188 (.A(in2[58]), .B(n_0_109), .ZN(sum[58]));
   XNOR2_X1 i_0_189 (.A(in3[58]), .B(in1[63]), .ZN(n_0_109));
   XNOR2_X1 i_0_190 (.A(in2[59]), .B(n_0_110), .ZN(sum[59]));
   XNOR2_X1 i_0_191 (.A(in3[59]), .B(in1[63]), .ZN(n_0_110));
   XNOR2_X1 i_0_192 (.A(in2[60]), .B(n_0_111), .ZN(sum[60]));
   XNOR2_X1 i_0_193 (.A(in3[60]), .B(in1[63]), .ZN(n_0_111));
   XNOR2_X1 i_0_194 (.A(in2[61]), .B(n_0_112), .ZN(sum[61]));
   XNOR2_X1 i_0_195 (.A(in3[61]), .B(in1[63]), .ZN(n_0_112));
   XOR2_X1 i_0_196 (.A(in3[62]), .B(n_0_113), .Z(sum[62]));
   XOR2_X1 i_0_197 (.A(in3[63]), .B(n_0_113), .Z(sum[63]));
   XOR2_X1 i_0_198 (.A(in2[63]), .B(in1[63]), .Z(n_0_113));
endmodule

module CSA__4_14(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;

   AND2_X1 i_0_0 (.A1(in2[6]), .A2(in1[6]), .ZN(c[7]));
   AND2_X1 i_0_1 (.A1(in2[7]), .A2(in1[7]), .ZN(c[8]));
   AND2_X1 i_0_2 (.A1(in2[8]), .A2(in1[8]), .ZN(c[9]));
   AND2_X1 i_0_3 (.A1(in2[9]), .A2(in1[9]), .ZN(c[10]));
   AND2_X1 i_0_4 (.A1(in2[10]), .A2(in1[10]), .ZN(c[11]));
   AND2_X1 i_0_5 (.A1(in2[11]), .A2(in1[11]), .ZN(c[12]));
   AND2_X1 i_0_6 (.A1(in2[12]), .A2(in1[12]), .ZN(c[13]));
   AND2_X1 i_0_7 (.A1(in2[13]), .A2(in1[13]), .ZN(c[14]));
   AND2_X1 i_0_8 (.A1(in2[14]), .A2(in1[14]), .ZN(c[15]));
   NAND2_X1 i_0_9 (.A1(n_0_1), .A2(n_0_0), .ZN(c[16]));
   OAI21_X1 i_0_10 (.A(in2[15]), .B1(in3[15]), .B2(in1[15]), .ZN(n_0_0));
   NAND2_X1 i_0_11 (.A1(in3[15]), .A2(in1[15]), .ZN(n_0_1));
   NAND2_X1 i_0_12 (.A1(n_0_3), .A2(n_0_2), .ZN(c[17]));
   OAI21_X1 i_0_13 (.A(in2[16]), .B1(in3[16]), .B2(in1[16]), .ZN(n_0_2));
   NAND2_X1 i_0_14 (.A1(in3[16]), .A2(in1[16]), .ZN(n_0_3));
   NAND2_X1 i_0_15 (.A1(n_0_5), .A2(n_0_4), .ZN(c[18]));
   OAI21_X1 i_0_16 (.A(in2[17]), .B1(in3[17]), .B2(in1[17]), .ZN(n_0_4));
   NAND2_X1 i_0_17 (.A1(in3[17]), .A2(in1[17]), .ZN(n_0_5));
   NAND2_X1 i_0_18 (.A1(n_0_7), .A2(n_0_6), .ZN(c[19]));
   OAI21_X1 i_0_19 (.A(in2[18]), .B1(in3[18]), .B2(in1[18]), .ZN(n_0_6));
   NAND2_X1 i_0_20 (.A1(in3[18]), .A2(in1[18]), .ZN(n_0_7));
   NAND2_X1 i_0_21 (.A1(n_0_9), .A2(n_0_8), .ZN(c[20]));
   OAI21_X1 i_0_22 (.A(in2[19]), .B1(in3[19]), .B2(in1[19]), .ZN(n_0_8));
   NAND2_X1 i_0_23 (.A1(in3[19]), .A2(in1[19]), .ZN(n_0_9));
   NAND2_X1 i_0_24 (.A1(n_0_11), .A2(n_0_10), .ZN(c[21]));
   OAI21_X1 i_0_25 (.A(in2[20]), .B1(in3[20]), .B2(in1[20]), .ZN(n_0_10));
   NAND2_X1 i_0_26 (.A1(in3[20]), .A2(in1[20]), .ZN(n_0_11));
   NAND2_X1 i_0_27 (.A1(n_0_13), .A2(n_0_12), .ZN(c[22]));
   OAI21_X1 i_0_28 (.A(in2[21]), .B1(in3[21]), .B2(in1[21]), .ZN(n_0_12));
   NAND2_X1 i_0_29 (.A1(in3[21]), .A2(in1[21]), .ZN(n_0_13));
   NAND2_X1 i_0_30 (.A1(n_0_15), .A2(n_0_14), .ZN(c[23]));
   OAI21_X1 i_0_31 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_14));
   NAND2_X1 i_0_32 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_15));
   NAND2_X1 i_0_33 (.A1(n_0_17), .A2(n_0_16), .ZN(c[24]));
   OAI21_X1 i_0_34 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_16));
   NAND2_X1 i_0_35 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_17));
   NAND2_X1 i_0_36 (.A1(n_0_19), .A2(n_0_18), .ZN(c[25]));
   OAI21_X1 i_0_37 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_18));
   NAND2_X1 i_0_38 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_19));
   NAND2_X1 i_0_39 (.A1(n_0_21), .A2(n_0_20), .ZN(c[26]));
   OAI21_X1 i_0_40 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_20));
   NAND2_X1 i_0_41 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_21));
   NAND2_X1 i_0_42 (.A1(n_0_23), .A2(n_0_22), .ZN(c[27]));
   OAI21_X1 i_0_43 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_22));
   NAND2_X1 i_0_44 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_23));
   NAND2_X1 i_0_45 (.A1(n_0_25), .A2(n_0_24), .ZN(c[28]));
   OAI21_X1 i_0_46 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_24));
   NAND2_X1 i_0_47 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_25));
   NAND2_X1 i_0_48 (.A1(n_0_27), .A2(n_0_26), .ZN(c[29]));
   OAI21_X1 i_0_49 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_26));
   NAND2_X1 i_0_50 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_27));
   NAND2_X1 i_0_51 (.A1(n_0_29), .A2(n_0_28), .ZN(c[30]));
   OAI21_X1 i_0_52 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_28));
   NAND2_X1 i_0_53 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_29));
   NAND2_X1 i_0_54 (.A1(n_0_31), .A2(n_0_30), .ZN(c[31]));
   OAI21_X1 i_0_55 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_30));
   NAND2_X1 i_0_56 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_31));
   NAND2_X1 i_0_57 (.A1(n_0_33), .A2(n_0_32), .ZN(c[32]));
   OAI21_X1 i_0_58 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_32));
   NAND2_X1 i_0_59 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_33));
   NAND2_X1 i_0_60 (.A1(n_0_35), .A2(n_0_34), .ZN(c[33]));
   OAI21_X1 i_0_61 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_34));
   NAND2_X1 i_0_62 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_35));
   NAND2_X1 i_0_63 (.A1(n_0_37), .A2(n_0_36), .ZN(c[34]));
   OAI21_X1 i_0_64 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_36));
   NAND2_X1 i_0_65 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_37));
   NAND2_X1 i_0_66 (.A1(n_0_39), .A2(n_0_38), .ZN(c[35]));
   OAI21_X1 i_0_67 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_38));
   NAND2_X1 i_0_68 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_39));
   NAND2_X1 i_0_69 (.A1(n_0_41), .A2(n_0_40), .ZN(c[36]));
   OAI21_X1 i_0_70 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_40));
   NAND2_X1 i_0_71 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_41));
   NAND2_X1 i_0_72 (.A1(n_0_43), .A2(n_0_42), .ZN(c[37]));
   OAI21_X1 i_0_73 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_42));
   NAND2_X1 i_0_74 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_43));
   NAND2_X1 i_0_75 (.A1(n_0_45), .A2(n_0_44), .ZN(c[38]));
   OAI21_X1 i_0_76 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_44));
   NAND2_X1 i_0_77 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_45));
   NAND2_X1 i_0_78 (.A1(n_0_47), .A2(n_0_46), .ZN(c[39]));
   OAI21_X1 i_0_79 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_46));
   NAND2_X1 i_0_80 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_47));
   NAND2_X1 i_0_81 (.A1(n_0_49), .A2(n_0_48), .ZN(c[40]));
   OAI21_X1 i_0_82 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_48));
   NAND2_X1 i_0_83 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_49));
   NAND2_X1 i_0_84 (.A1(n_0_51), .A2(n_0_50), .ZN(c[41]));
   OAI21_X1 i_0_85 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_50));
   NAND2_X1 i_0_86 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_51));
   NAND2_X1 i_0_87 (.A1(n_0_53), .A2(n_0_52), .ZN(c[42]));
   OAI21_X1 i_0_88 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_52));
   NAND2_X1 i_0_89 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_53));
   NAND2_X1 i_0_90 (.A1(n_0_55), .A2(n_0_54), .ZN(c[43]));
   OAI21_X1 i_0_91 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_54));
   NAND2_X1 i_0_92 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_55));
   NAND2_X1 i_0_93 (.A1(n_0_57), .A2(n_0_56), .ZN(c[44]));
   OAI21_X1 i_0_94 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_56));
   NAND2_X1 i_0_95 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_57));
   NAND2_X1 i_0_96 (.A1(n_0_59), .A2(n_0_58), .ZN(c[45]));
   OAI21_X1 i_0_97 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_58));
   NAND2_X1 i_0_98 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_59));
   NAND2_X1 i_0_99 (.A1(n_0_61), .A2(n_0_60), .ZN(c[46]));
   OAI21_X1 i_0_100 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_60));
   NAND2_X1 i_0_101 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_61));
   NAND2_X1 i_0_102 (.A1(n_0_63), .A2(n_0_62), .ZN(c[47]));
   OAI21_X1 i_0_103 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_62));
   NAND2_X1 i_0_104 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_63));
   NAND2_X1 i_0_105 (.A1(n_0_65), .A2(n_0_64), .ZN(c[48]));
   OAI21_X1 i_0_106 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_64));
   NAND2_X1 i_0_107 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_65));
   NAND2_X1 i_0_108 (.A1(n_0_67), .A2(n_0_66), .ZN(c[49]));
   OAI21_X1 i_0_109 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_66));
   NAND2_X1 i_0_110 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_67));
   NAND2_X1 i_0_111 (.A1(n_0_69), .A2(n_0_68), .ZN(c[50]));
   OAI21_X1 i_0_112 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_68));
   NAND2_X1 i_0_113 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_69));
   NAND2_X1 i_0_114 (.A1(n_0_71), .A2(n_0_70), .ZN(c[51]));
   OAI21_X1 i_0_115 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_70));
   NAND2_X1 i_0_116 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_71));
   NAND2_X1 i_0_117 (.A1(n_0_73), .A2(n_0_72), .ZN(c[52]));
   OAI21_X1 i_0_118 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_72));
   NAND2_X1 i_0_119 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_73));
   NAND2_X1 i_0_120 (.A1(n_0_75), .A2(n_0_74), .ZN(c[53]));
   OAI21_X1 i_0_121 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_74));
   NAND2_X1 i_0_122 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_75));
   NAND2_X1 i_0_123 (.A1(n_0_77), .A2(n_0_76), .ZN(c[54]));
   OAI21_X1 i_0_124 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_76));
   NAND2_X1 i_0_125 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_77));
   NAND2_X1 i_0_126 (.A1(n_0_79), .A2(n_0_78), .ZN(c[55]));
   OAI21_X1 i_0_127 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_78));
   NAND2_X1 i_0_128 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_79));
   NAND2_X1 i_0_129 (.A1(n_0_81), .A2(n_0_80), .ZN(c[56]));
   OAI21_X1 i_0_130 (.A(in2[55]), .B1(in3[55]), .B2(in1[63]), .ZN(n_0_80));
   NAND2_X1 i_0_131 (.A1(in3[55]), .A2(in1[63]), .ZN(n_0_81));
   AOI21_X1 i_0_132 (.A(n_0_83), .B1(n_0_82), .B2(n_0_126), .ZN(c[57]));
   AOI21_X1 i_0_133 (.A(n_0_83), .B1(n_0_82), .B2(n_0_127), .ZN(c[58]));
   AOI21_X1 i_0_134 (.A(n_0_83), .B1(n_0_82), .B2(n_0_128), .ZN(c[59]));
   AOI21_X1 i_0_135 (.A(n_0_83), .B1(n_0_82), .B2(n_0_129), .ZN(c[60]));
   AOI21_X1 i_0_136 (.A(n_0_83), .B1(n_0_82), .B2(n_0_130), .ZN(c[61]));
   AOI21_X1 i_0_137 (.A(n_0_83), .B1(n_0_82), .B2(n_0_131), .ZN(c[62]));
   AOI21_X1 i_0_138 (.A(n_0_83), .B1(n_0_82), .B2(n_0_132), .ZN(c[63]));
   NAND2_X1 i_0_139 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_82));
   NOR2_X1 i_0_140 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_83));
   XOR2_X1 i_0_141 (.A(in2[6]), .B(in1[6]), .Z(sum[6]));
   XOR2_X1 i_0_142 (.A(in2[7]), .B(in1[7]), .Z(sum[7]));
   XOR2_X1 i_0_143 (.A(in2[8]), .B(in1[8]), .Z(sum[8]));
   XOR2_X1 i_0_144 (.A(in2[9]), .B(in1[9]), .Z(sum[9]));
   XOR2_X1 i_0_145 (.A(in2[10]), .B(in1[10]), .Z(sum[10]));
   XOR2_X1 i_0_146 (.A(in2[11]), .B(in1[11]), .Z(sum[11]));
   XOR2_X1 i_0_147 (.A(in2[12]), .B(in1[12]), .Z(sum[12]));
   XOR2_X1 i_0_148 (.A(in2[13]), .B(in1[13]), .Z(sum[13]));
   XOR2_X1 i_0_149 (.A(in2[14]), .B(in1[14]), .Z(sum[14]));
   XNOR2_X1 i_0_150 (.A(in2[15]), .B(n_0_84), .ZN(sum[15]));
   XNOR2_X1 i_0_151 (.A(in3[15]), .B(in1[15]), .ZN(n_0_84));
   XNOR2_X1 i_0_152 (.A(in2[16]), .B(n_0_85), .ZN(sum[16]));
   XNOR2_X1 i_0_153 (.A(in3[16]), .B(in1[16]), .ZN(n_0_85));
   XNOR2_X1 i_0_154 (.A(in2[17]), .B(n_0_86), .ZN(sum[17]));
   XNOR2_X1 i_0_155 (.A(in3[17]), .B(in1[17]), .ZN(n_0_86));
   XNOR2_X1 i_0_156 (.A(in2[18]), .B(n_0_87), .ZN(sum[18]));
   XNOR2_X1 i_0_157 (.A(in3[18]), .B(in1[18]), .ZN(n_0_87));
   XNOR2_X1 i_0_158 (.A(in2[19]), .B(n_0_88), .ZN(sum[19]));
   XNOR2_X1 i_0_159 (.A(in3[19]), .B(in1[19]), .ZN(n_0_88));
   XNOR2_X1 i_0_160 (.A(in2[20]), .B(n_0_89), .ZN(sum[20]));
   XNOR2_X1 i_0_161 (.A(in3[20]), .B(in1[20]), .ZN(n_0_89));
   XNOR2_X1 i_0_162 (.A(in2[21]), .B(n_0_90), .ZN(sum[21]));
   XNOR2_X1 i_0_163 (.A(in3[21]), .B(in1[21]), .ZN(n_0_90));
   XNOR2_X1 i_0_164 (.A(in2[22]), .B(n_0_91), .ZN(sum[22]));
   XNOR2_X1 i_0_165 (.A(in3[22]), .B(in1[22]), .ZN(n_0_91));
   XNOR2_X1 i_0_166 (.A(in2[23]), .B(n_0_92), .ZN(sum[23]));
   XNOR2_X1 i_0_167 (.A(in3[23]), .B(in1[23]), .ZN(n_0_92));
   XNOR2_X1 i_0_168 (.A(in2[24]), .B(n_0_93), .ZN(sum[24]));
   XNOR2_X1 i_0_169 (.A(in3[24]), .B(in1[24]), .ZN(n_0_93));
   XNOR2_X1 i_0_170 (.A(in2[25]), .B(n_0_94), .ZN(sum[25]));
   XNOR2_X1 i_0_171 (.A(in3[25]), .B(in1[25]), .ZN(n_0_94));
   XNOR2_X1 i_0_172 (.A(in2[26]), .B(n_0_95), .ZN(sum[26]));
   XNOR2_X1 i_0_173 (.A(in3[26]), .B(in1[26]), .ZN(n_0_95));
   XNOR2_X1 i_0_174 (.A(in2[27]), .B(n_0_96), .ZN(sum[27]));
   XNOR2_X1 i_0_175 (.A(in3[27]), .B(in1[27]), .ZN(n_0_96));
   XNOR2_X1 i_0_176 (.A(in2[28]), .B(n_0_97), .ZN(sum[28]));
   XNOR2_X1 i_0_177 (.A(in3[28]), .B(in1[28]), .ZN(n_0_97));
   XNOR2_X1 i_0_178 (.A(in2[29]), .B(n_0_98), .ZN(sum[29]));
   XNOR2_X1 i_0_179 (.A(in3[29]), .B(in1[29]), .ZN(n_0_98));
   XNOR2_X1 i_0_180 (.A(in2[30]), .B(n_0_99), .ZN(sum[30]));
   XNOR2_X1 i_0_181 (.A(in3[30]), .B(in1[30]), .ZN(n_0_99));
   XNOR2_X1 i_0_182 (.A(in2[31]), .B(n_0_100), .ZN(sum[31]));
   XNOR2_X1 i_0_183 (.A(in3[31]), .B(in1[31]), .ZN(n_0_100));
   XNOR2_X1 i_0_184 (.A(in2[32]), .B(n_0_101), .ZN(sum[32]));
   XNOR2_X1 i_0_185 (.A(in3[32]), .B(in1[32]), .ZN(n_0_101));
   XNOR2_X1 i_0_186 (.A(in2[33]), .B(n_0_102), .ZN(sum[33]));
   XNOR2_X1 i_0_187 (.A(in3[33]), .B(in1[33]), .ZN(n_0_102));
   XNOR2_X1 i_0_188 (.A(in2[34]), .B(n_0_103), .ZN(sum[34]));
   XNOR2_X1 i_0_189 (.A(in3[34]), .B(in1[34]), .ZN(n_0_103));
   XNOR2_X1 i_0_190 (.A(in2[35]), .B(n_0_104), .ZN(sum[35]));
   XNOR2_X1 i_0_191 (.A(in3[35]), .B(in1[35]), .ZN(n_0_104));
   XNOR2_X1 i_0_192 (.A(in2[36]), .B(n_0_105), .ZN(sum[36]));
   XNOR2_X1 i_0_193 (.A(in3[36]), .B(in1[36]), .ZN(n_0_105));
   XNOR2_X1 i_0_194 (.A(in2[37]), .B(n_0_106), .ZN(sum[37]));
   XNOR2_X1 i_0_195 (.A(in3[37]), .B(in1[37]), .ZN(n_0_106));
   XNOR2_X1 i_0_196 (.A(in2[38]), .B(n_0_107), .ZN(sum[38]));
   XNOR2_X1 i_0_197 (.A(in3[38]), .B(in1[38]), .ZN(n_0_107));
   XNOR2_X1 i_0_198 (.A(in2[39]), .B(n_0_108), .ZN(sum[39]));
   XNOR2_X1 i_0_199 (.A(in3[39]), .B(in1[39]), .ZN(n_0_108));
   XNOR2_X1 i_0_200 (.A(in2[40]), .B(n_0_109), .ZN(sum[40]));
   XNOR2_X1 i_0_201 (.A(in3[40]), .B(in1[40]), .ZN(n_0_109));
   XNOR2_X1 i_0_202 (.A(in2[41]), .B(n_0_110), .ZN(sum[41]));
   XNOR2_X1 i_0_203 (.A(in3[41]), .B(in1[41]), .ZN(n_0_110));
   XNOR2_X1 i_0_204 (.A(in2[42]), .B(n_0_111), .ZN(sum[42]));
   XNOR2_X1 i_0_205 (.A(in3[42]), .B(in1[42]), .ZN(n_0_111));
   XNOR2_X1 i_0_206 (.A(in2[43]), .B(n_0_112), .ZN(sum[43]));
   XNOR2_X1 i_0_207 (.A(in3[43]), .B(in1[43]), .ZN(n_0_112));
   XNOR2_X1 i_0_208 (.A(in2[44]), .B(n_0_113), .ZN(sum[44]));
   XNOR2_X1 i_0_209 (.A(in3[44]), .B(in1[44]), .ZN(n_0_113));
   XNOR2_X1 i_0_210 (.A(in2[45]), .B(n_0_114), .ZN(sum[45]));
   XNOR2_X1 i_0_211 (.A(in3[45]), .B(in1[45]), .ZN(n_0_114));
   XNOR2_X1 i_0_212 (.A(in2[46]), .B(n_0_115), .ZN(sum[46]));
   XNOR2_X1 i_0_213 (.A(in3[46]), .B(in1[46]), .ZN(n_0_115));
   XNOR2_X1 i_0_220 (.A(in2[50]), .B(n_0_119), .ZN(sum[50]));
   XNOR2_X1 i_0_221 (.A(in3[50]), .B(in1[50]), .ZN(n_0_119));
   XNOR2_X1 i_0_222 (.A(in2[51]), .B(n_0_120), .ZN(sum[51]));
   XNOR2_X1 i_0_223 (.A(in3[51]), .B(in1[51]), .ZN(n_0_120));
   XNOR2_X1 i_0_224 (.A(in2[52]), .B(n_0_121), .ZN(sum[52]));
   XNOR2_X1 i_0_225 (.A(in3[52]), .B(in1[52]), .ZN(n_0_121));
   XNOR2_X1 i_0_226 (.A(in2[53]), .B(n_0_122), .ZN(sum[53]));
   XNOR2_X1 i_0_227 (.A(in3[53]), .B(in1[53]), .ZN(n_0_122));
   XNOR2_X1 i_0_228 (.A(in2[54]), .B(n_0_123), .ZN(sum[54]));
   XNOR2_X1 i_0_229 (.A(in3[54]), .B(in1[54]), .ZN(n_0_123));
   XNOR2_X1 i_0_230 (.A(in2[55]), .B(n_0_124), .ZN(sum[55]));
   XNOR2_X1 i_0_231 (.A(in3[55]), .B(in1[63]), .ZN(n_0_124));
   XNOR2_X1 i_0_232 (.A(n_0_126), .B(n_0_125), .ZN(sum[56]));
   XNOR2_X1 i_0_233 (.A(n_0_127), .B(n_0_125), .ZN(sum[57]));
   XNOR2_X1 i_0_234 (.A(n_0_128), .B(n_0_125), .ZN(sum[58]));
   XNOR2_X1 i_0_235 (.A(n_0_129), .B(n_0_125), .ZN(sum[59]));
   XNOR2_X1 i_0_236 (.A(n_0_130), .B(n_0_125), .ZN(sum[60]));
   XNOR2_X1 i_0_237 (.A(n_0_131), .B(n_0_125), .ZN(sum[61]));
   XNOR2_X1 i_0_238 (.A(n_0_132), .B(n_0_125), .ZN(sum[62]));
   XOR2_X1 i_0_239 (.A(in3[63]), .B(n_0_125), .Z(sum[63]));
   XOR2_X1 i_0_240 (.A(in2[63]), .B(in1[63]), .Z(n_0_125));
   INV_X1 i_0_241 (.A(in3[56]), .ZN(n_0_126));
   INV_X1 i_0_242 (.A(in3[57]), .ZN(n_0_127));
   INV_X1 i_0_243 (.A(in3[58]), .ZN(n_0_128));
   INV_X1 i_0_244 (.A(in3[59]), .ZN(n_0_129));
   INV_X1 i_0_245 (.A(in3[60]), .ZN(n_0_130));
   INV_X1 i_0_246 (.A(in3[61]), .ZN(n_0_131));
   INV_X1 i_0_247 (.A(in3[62]), .ZN(n_0_132));
   XOR2_X1 i_0_214 (.A(in2[47]), .B(n_0_116), .Z(sum[47]));
   XOR2_X1 i_0_215 (.A(in3[47]), .B(in1[47]), .Z(n_0_116));
   XOR2_X1 i_0_216 (.A(in2[48]), .B(n_0_117), .Z(sum[48]));
   XOR2_X1 i_0_217 (.A(in3[48]), .B(in1[48]), .Z(n_0_117));
   XOR2_X1 i_0_218 (.A(in2[49]), .B(n_0_118), .Z(sum[49]));
   XOR2_X1 i_0_219 (.A(in3[49]), .B(in1[49]), .Z(n_0_118));
endmodule

module CSA__4_17(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;

   AND2_X1 i_0_0 (.A1(in2[7]), .A2(in1[7]), .ZN(c[8]));
   AND2_X1 i_0_1 (.A1(in2[8]), .A2(in1[8]), .ZN(c[9]));
   AND2_X1 i_0_2 (.A1(in2[9]), .A2(in1[9]), .ZN(c[10]));
   AND2_X1 i_0_3 (.A1(in2[10]), .A2(in1[10]), .ZN(c[11]));
   AND2_X1 i_0_4 (.A1(in2[11]), .A2(in1[11]), .ZN(c[12]));
   AND2_X1 i_0_5 (.A1(in2[12]), .A2(in1[12]), .ZN(c[13]));
   AND2_X1 i_0_6 (.A1(in2[13]), .A2(in1[13]), .ZN(c[14]));
   AND2_X1 i_0_7 (.A1(in2[14]), .A2(in1[14]), .ZN(c[15]));
   AND2_X1 i_0_8 (.A1(in2[15]), .A2(in1[15]), .ZN(c[16]));
   AND2_X1 i_0_9 (.A1(in2[16]), .A2(in1[16]), .ZN(c[17]));
   AND2_X1 i_0_10 (.A1(in2[17]), .A2(in1[17]), .ZN(c[18]));
   AND2_X1 i_0_11 (.A1(in2[18]), .A2(in1[18]), .ZN(c[19]));
   AND2_X1 i_0_12 (.A1(in2[19]), .A2(in1[19]), .ZN(c[20]));
   AND2_X1 i_0_13 (.A1(in2[20]), .A2(in1[20]), .ZN(c[21]));
   AND2_X1 i_0_14 (.A1(in2[21]), .A2(in1[21]), .ZN(c[22]));
   NAND2_X1 i_0_15 (.A1(n_0_1), .A2(n_0_0), .ZN(c[23]));
   OAI21_X1 i_0_16 (.A(in2[22]), .B1(in3[22]), .B2(in1[22]), .ZN(n_0_0));
   NAND2_X1 i_0_17 (.A1(in3[22]), .A2(in1[22]), .ZN(n_0_1));
   NAND2_X1 i_0_18 (.A1(n_0_3), .A2(n_0_2), .ZN(c[24]));
   OAI21_X1 i_0_19 (.A(in2[23]), .B1(in3[23]), .B2(in1[23]), .ZN(n_0_2));
   NAND2_X1 i_0_20 (.A1(in3[23]), .A2(in1[23]), .ZN(n_0_3));
   NAND2_X1 i_0_21 (.A1(n_0_5), .A2(n_0_4), .ZN(c[25]));
   OAI21_X1 i_0_22 (.A(in2[24]), .B1(in3[24]), .B2(in1[24]), .ZN(n_0_4));
   NAND2_X1 i_0_23 (.A1(in3[24]), .A2(in1[24]), .ZN(n_0_5));
   NAND2_X1 i_0_24 (.A1(n_0_7), .A2(n_0_6), .ZN(c[26]));
   OAI21_X1 i_0_25 (.A(in2[25]), .B1(in3[25]), .B2(in1[25]), .ZN(n_0_6));
   NAND2_X1 i_0_26 (.A1(in3[25]), .A2(in1[25]), .ZN(n_0_7));
   NAND2_X1 i_0_27 (.A1(n_0_9), .A2(n_0_8), .ZN(c[27]));
   OAI21_X1 i_0_28 (.A(in2[26]), .B1(in3[26]), .B2(in1[26]), .ZN(n_0_8));
   NAND2_X1 i_0_29 (.A1(in3[26]), .A2(in1[26]), .ZN(n_0_9));
   NAND2_X1 i_0_30 (.A1(n_0_11), .A2(n_0_10), .ZN(c[28]));
   OAI21_X1 i_0_31 (.A(in2[27]), .B1(in3[27]), .B2(in1[27]), .ZN(n_0_10));
   NAND2_X1 i_0_32 (.A1(in3[27]), .A2(in1[27]), .ZN(n_0_11));
   NAND2_X1 i_0_33 (.A1(n_0_13), .A2(n_0_12), .ZN(c[29]));
   OAI21_X1 i_0_34 (.A(in2[28]), .B1(in3[28]), .B2(in1[28]), .ZN(n_0_12));
   NAND2_X1 i_0_35 (.A1(in3[28]), .A2(in1[28]), .ZN(n_0_13));
   NAND2_X1 i_0_36 (.A1(n_0_15), .A2(n_0_14), .ZN(c[30]));
   OAI21_X1 i_0_37 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_14));
   NAND2_X1 i_0_38 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_15));
   NAND2_X1 i_0_39 (.A1(n_0_17), .A2(n_0_16), .ZN(c[31]));
   OAI21_X1 i_0_40 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_16));
   NAND2_X1 i_0_41 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_17));
   NAND2_X1 i_0_42 (.A1(n_0_19), .A2(n_0_18), .ZN(c[32]));
   OAI21_X1 i_0_43 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_18));
   NAND2_X1 i_0_44 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_19));
   NAND2_X1 i_0_45 (.A1(n_0_21), .A2(n_0_20), .ZN(c[33]));
   OAI21_X1 i_0_46 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_20));
   NAND2_X1 i_0_47 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_21));
   NAND2_X1 i_0_48 (.A1(n_0_23), .A2(n_0_22), .ZN(c[34]));
   OAI21_X1 i_0_49 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_22));
   NAND2_X1 i_0_50 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_23));
   NAND2_X1 i_0_51 (.A1(n_0_25), .A2(n_0_24), .ZN(c[35]));
   OAI21_X1 i_0_52 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_24));
   NAND2_X1 i_0_53 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_25));
   NAND2_X1 i_0_54 (.A1(n_0_27), .A2(n_0_26), .ZN(c[36]));
   OAI21_X1 i_0_55 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_26));
   NAND2_X1 i_0_56 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_27));
   NAND2_X1 i_0_57 (.A1(n_0_29), .A2(n_0_28), .ZN(c[37]));
   OAI21_X1 i_0_58 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_28));
   NAND2_X1 i_0_59 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_29));
   NAND2_X1 i_0_60 (.A1(n_0_31), .A2(n_0_30), .ZN(c[38]));
   OAI21_X1 i_0_61 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_30));
   NAND2_X1 i_0_62 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_31));
   NAND2_X1 i_0_63 (.A1(n_0_33), .A2(n_0_32), .ZN(c[39]));
   OAI21_X1 i_0_64 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_32));
   NAND2_X1 i_0_65 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_33));
   NAND2_X1 i_0_66 (.A1(n_0_35), .A2(n_0_34), .ZN(c[40]));
   OAI21_X1 i_0_67 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_34));
   NAND2_X1 i_0_68 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_35));
   NAND2_X1 i_0_69 (.A1(n_0_37), .A2(n_0_36), .ZN(c[41]));
   OAI21_X1 i_0_70 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_36));
   NAND2_X1 i_0_71 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_37));
   NAND2_X1 i_0_72 (.A1(n_0_39), .A2(n_0_38), .ZN(c[42]));
   OAI21_X1 i_0_73 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_38));
   NAND2_X1 i_0_74 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_39));
   NAND2_X1 i_0_75 (.A1(n_0_41), .A2(n_0_40), .ZN(c[43]));
   OAI21_X1 i_0_76 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_40));
   NAND2_X1 i_0_77 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_41));
   NAND2_X1 i_0_78 (.A1(n_0_43), .A2(n_0_42), .ZN(c[44]));
   OAI21_X1 i_0_79 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_42));
   NAND2_X1 i_0_80 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_43));
   NAND2_X1 i_0_81 (.A1(n_0_45), .A2(n_0_44), .ZN(c[45]));
   OAI21_X1 i_0_82 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_44));
   NAND2_X1 i_0_83 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_45));
   NAND2_X1 i_0_84 (.A1(n_0_47), .A2(n_0_46), .ZN(c[46]));
   OAI21_X1 i_0_85 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_46));
   NAND2_X1 i_0_86 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_47));
   NAND2_X1 i_0_87 (.A1(n_0_49), .A2(n_0_48), .ZN(c[47]));
   OAI21_X1 i_0_88 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_48));
   NAND2_X1 i_0_89 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_49));
   NAND2_X1 i_0_90 (.A1(n_0_51), .A2(n_0_50), .ZN(c[48]));
   OAI21_X1 i_0_91 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_50));
   NAND2_X1 i_0_92 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_51));
   NAND2_X1 i_0_93 (.A1(n_0_53), .A2(n_0_52), .ZN(c[49]));
   OAI21_X1 i_0_94 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_52));
   NAND2_X1 i_0_95 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_53));
   NAND2_X1 i_0_96 (.A1(n_0_55), .A2(n_0_54), .ZN(c[50]));
   OAI21_X1 i_0_97 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_54));
   NAND2_X1 i_0_98 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_55));
   NAND2_X1 i_0_99 (.A1(n_0_57), .A2(n_0_56), .ZN(c[51]));
   OAI21_X1 i_0_100 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_56));
   NAND2_X1 i_0_101 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_57));
   NAND2_X1 i_0_102 (.A1(n_0_59), .A2(n_0_58), .ZN(c[52]));
   OAI21_X1 i_0_103 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_58));
   NAND2_X1 i_0_104 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_59));
   NAND2_X1 i_0_105 (.A1(n_0_61), .A2(n_0_60), .ZN(c[53]));
   OAI21_X1 i_0_106 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_60));
   NAND2_X1 i_0_107 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_61));
   NAND2_X1 i_0_108 (.A1(n_0_63), .A2(n_0_62), .ZN(c[54]));
   OAI21_X1 i_0_109 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_62));
   NAND2_X1 i_0_110 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_63));
   NAND2_X1 i_0_111 (.A1(n_0_65), .A2(n_0_64), .ZN(c[55]));
   OAI21_X1 i_0_112 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_64));
   NAND2_X1 i_0_113 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_65));
   NAND2_X1 i_0_114 (.A1(n_0_67), .A2(n_0_66), .ZN(c[56]));
   OAI21_X1 i_0_115 (.A(in2[55]), .B1(in3[55]), .B2(in1[55]), .ZN(n_0_66));
   NAND2_X1 i_0_116 (.A1(in3[55]), .A2(in1[55]), .ZN(n_0_67));
   NAND2_X1 i_0_117 (.A1(n_0_69), .A2(n_0_68), .ZN(c[57]));
   OAI21_X1 i_0_118 (.A(in2[56]), .B1(in3[56]), .B2(in1[56]), .ZN(n_0_68));
   NAND2_X1 i_0_119 (.A1(in3[56]), .A2(in1[56]), .ZN(n_0_69));
   NAND2_X1 i_0_120 (.A1(n_0_71), .A2(n_0_70), .ZN(c[58]));
   OAI21_X1 i_0_121 (.A(in2[57]), .B1(in3[57]), .B2(in1[57]), .ZN(n_0_70));
   NAND2_X1 i_0_122 (.A1(in3[57]), .A2(in1[57]), .ZN(n_0_71));
   NAND2_X1 i_0_123 (.A1(n_0_73), .A2(n_0_72), .ZN(c[59]));
   OAI21_X1 i_0_124 (.A(in2[58]), .B1(in3[58]), .B2(in1[58]), .ZN(n_0_72));
   NAND2_X1 i_0_125 (.A1(in3[58]), .A2(in1[58]), .ZN(n_0_73));
   NAND2_X1 i_0_126 (.A1(n_0_75), .A2(n_0_74), .ZN(c[60]));
   OAI21_X1 i_0_127 (.A(in2[59]), .B1(in3[59]), .B2(in1[59]), .ZN(n_0_74));
   NAND2_X1 i_0_128 (.A1(in3[59]), .A2(in1[59]), .ZN(n_0_75));
   NAND2_X1 i_0_129 (.A1(n_0_77), .A2(n_0_76), .ZN(c[61]));
   OAI21_X1 i_0_130 (.A(in2[60]), .B1(in3[60]), .B2(in1[60]), .ZN(n_0_76));
   NAND2_X1 i_0_131 (.A1(in3[60]), .A2(in1[60]), .ZN(n_0_77));
   NAND2_X1 i_0_132 (.A1(n_0_79), .A2(n_0_78), .ZN(c[62]));
   OAI21_X1 i_0_133 (.A(in2[61]), .B1(in3[61]), .B2(in1[61]), .ZN(n_0_78));
   NAND2_X1 i_0_134 (.A1(in3[61]), .A2(in1[61]), .ZN(n_0_79));
   NAND2_X1 i_0_135 (.A1(n_0_81), .A2(n_0_80), .ZN(c[63]));
   OAI21_X1 i_0_136 (.A(in2[62]), .B1(in3[62]), .B2(in1[62]), .ZN(n_0_80));
   NAND2_X1 i_0_137 (.A1(in3[62]), .A2(in1[62]), .ZN(n_0_81));
   XOR2_X1 i_0_138 (.A(in2[7]), .B(in1[7]), .Z(sum[7]));
   XOR2_X1 i_0_139 (.A(in2[8]), .B(in1[8]), .Z(sum[8]));
   XOR2_X1 i_0_140 (.A(in2[9]), .B(in1[9]), .Z(sum[9]));
   XOR2_X1 i_0_141 (.A(in2[10]), .B(in1[10]), .Z(sum[10]));
   XOR2_X1 i_0_142 (.A(in2[11]), .B(in1[11]), .Z(sum[11]));
   XOR2_X1 i_0_143 (.A(in2[12]), .B(in1[12]), .Z(sum[12]));
   XOR2_X1 i_0_144 (.A(in2[13]), .B(in1[13]), .Z(sum[13]));
   XOR2_X1 i_0_145 (.A(in2[14]), .B(in1[14]), .Z(sum[14]));
   XOR2_X1 i_0_146 (.A(in2[15]), .B(in1[15]), .Z(sum[15]));
   XOR2_X1 i_0_147 (.A(in2[16]), .B(in1[16]), .Z(sum[16]));
   XOR2_X1 i_0_148 (.A(in2[17]), .B(in1[17]), .Z(sum[17]));
   XOR2_X1 i_0_149 (.A(in2[18]), .B(in1[18]), .Z(sum[18]));
   XOR2_X1 i_0_150 (.A(in2[19]), .B(in1[19]), .Z(sum[19]));
   XOR2_X1 i_0_151 (.A(in2[20]), .B(in1[20]), .Z(sum[20]));
   XOR2_X1 i_0_152 (.A(in2[21]), .B(in1[21]), .Z(sum[21]));
   XNOR2_X1 i_0_153 (.A(in2[22]), .B(n_0_82), .ZN(sum[22]));
   XNOR2_X1 i_0_154 (.A(in3[22]), .B(in1[22]), .ZN(n_0_82));
   XNOR2_X1 i_0_155 (.A(in2[23]), .B(n_0_83), .ZN(sum[23]));
   XNOR2_X1 i_0_156 (.A(in3[23]), .B(in1[23]), .ZN(n_0_83));
   XNOR2_X1 i_0_157 (.A(in2[24]), .B(n_0_84), .ZN(sum[24]));
   XNOR2_X1 i_0_158 (.A(in3[24]), .B(in1[24]), .ZN(n_0_84));
   XNOR2_X1 i_0_159 (.A(in2[25]), .B(n_0_85), .ZN(sum[25]));
   XNOR2_X1 i_0_160 (.A(in3[25]), .B(in1[25]), .ZN(n_0_85));
   XNOR2_X1 i_0_161 (.A(in2[26]), .B(n_0_86), .ZN(sum[26]));
   XNOR2_X1 i_0_162 (.A(in3[26]), .B(in1[26]), .ZN(n_0_86));
   XNOR2_X1 i_0_163 (.A(in2[27]), .B(n_0_87), .ZN(sum[27]));
   XNOR2_X1 i_0_164 (.A(in3[27]), .B(in1[27]), .ZN(n_0_87));
   XNOR2_X1 i_0_165 (.A(in2[28]), .B(n_0_88), .ZN(sum[28]));
   XNOR2_X1 i_0_166 (.A(in3[28]), .B(in1[28]), .ZN(n_0_88));
   XNOR2_X1 i_0_167 (.A(in2[29]), .B(n_0_89), .ZN(sum[29]));
   XNOR2_X1 i_0_168 (.A(in3[29]), .B(in1[29]), .ZN(n_0_89));
   XNOR2_X1 i_0_169 (.A(in2[30]), .B(n_0_90), .ZN(sum[30]));
   XNOR2_X1 i_0_170 (.A(in3[30]), .B(in1[30]), .ZN(n_0_90));
   XNOR2_X1 i_0_171 (.A(in2[31]), .B(n_0_91), .ZN(sum[31]));
   XNOR2_X1 i_0_172 (.A(in3[31]), .B(in1[31]), .ZN(n_0_91));
   XNOR2_X1 i_0_173 (.A(in2[32]), .B(n_0_92), .ZN(sum[32]));
   XNOR2_X1 i_0_174 (.A(in3[32]), .B(in1[32]), .ZN(n_0_92));
   XNOR2_X1 i_0_175 (.A(in2[33]), .B(n_0_93), .ZN(sum[33]));
   XNOR2_X1 i_0_176 (.A(in3[33]), .B(in1[33]), .ZN(n_0_93));
   XNOR2_X1 i_0_177 (.A(in2[34]), .B(n_0_94), .ZN(sum[34]));
   XNOR2_X1 i_0_178 (.A(in3[34]), .B(in1[34]), .ZN(n_0_94));
   XNOR2_X1 i_0_179 (.A(in2[35]), .B(n_0_95), .ZN(sum[35]));
   XNOR2_X1 i_0_180 (.A(in3[35]), .B(in1[35]), .ZN(n_0_95));
   XNOR2_X1 i_0_181 (.A(in2[36]), .B(n_0_96), .ZN(sum[36]));
   XNOR2_X1 i_0_182 (.A(in3[36]), .B(in1[36]), .ZN(n_0_96));
   XNOR2_X1 i_0_183 (.A(in2[37]), .B(n_0_97), .ZN(sum[37]));
   XNOR2_X1 i_0_184 (.A(in3[37]), .B(in1[37]), .ZN(n_0_97));
   XNOR2_X1 i_0_185 (.A(in2[38]), .B(n_0_98), .ZN(sum[38]));
   XNOR2_X1 i_0_186 (.A(in3[38]), .B(in1[38]), .ZN(n_0_98));
   XNOR2_X1 i_0_187 (.A(in2[39]), .B(n_0_99), .ZN(sum[39]));
   XNOR2_X1 i_0_188 (.A(in3[39]), .B(in1[39]), .ZN(n_0_99));
   XNOR2_X1 i_0_189 (.A(in2[40]), .B(n_0_100), .ZN(sum[40]));
   XNOR2_X1 i_0_190 (.A(in3[40]), .B(in1[40]), .ZN(n_0_100));
   XNOR2_X1 i_0_191 (.A(in2[41]), .B(n_0_101), .ZN(sum[41]));
   XNOR2_X1 i_0_192 (.A(in3[41]), .B(in1[41]), .ZN(n_0_101));
   XNOR2_X1 i_0_193 (.A(in2[42]), .B(n_0_102), .ZN(sum[42]));
   XNOR2_X1 i_0_194 (.A(in3[42]), .B(in1[42]), .ZN(n_0_102));
   XNOR2_X1 i_0_195 (.A(in2[43]), .B(n_0_103), .ZN(sum[43]));
   XNOR2_X1 i_0_196 (.A(in3[43]), .B(in1[43]), .ZN(n_0_103));
   XNOR2_X1 i_0_197 (.A(in2[44]), .B(n_0_104), .ZN(sum[44]));
   XNOR2_X1 i_0_198 (.A(in3[44]), .B(in1[44]), .ZN(n_0_104));
   XNOR2_X1 i_0_199 (.A(in2[45]), .B(n_0_105), .ZN(sum[45]));
   XNOR2_X1 i_0_200 (.A(in3[45]), .B(in1[45]), .ZN(n_0_105));
   XNOR2_X1 i_0_201 (.A(in2[46]), .B(n_0_106), .ZN(sum[46]));
   XNOR2_X1 i_0_202 (.A(in3[46]), .B(in1[46]), .ZN(n_0_106));
   XNOR2_X1 i_0_209 (.A(in2[50]), .B(n_0_110), .ZN(sum[50]));
   XNOR2_X1 i_0_210 (.A(in3[50]), .B(in1[50]), .ZN(n_0_110));
   XNOR2_X1 i_0_211 (.A(in2[51]), .B(n_0_111), .ZN(sum[51]));
   XNOR2_X1 i_0_212 (.A(in3[51]), .B(in1[51]), .ZN(n_0_111));
   XNOR2_X1 i_0_213 (.A(in2[52]), .B(n_0_112), .ZN(sum[52]));
   XNOR2_X1 i_0_214 (.A(in3[52]), .B(in1[52]), .ZN(n_0_112));
   XNOR2_X1 i_0_215 (.A(in2[53]), .B(n_0_113), .ZN(sum[53]));
   XNOR2_X1 i_0_216 (.A(in3[53]), .B(in1[53]), .ZN(n_0_113));
   XNOR2_X1 i_0_217 (.A(in2[54]), .B(n_0_114), .ZN(sum[54]));
   XNOR2_X1 i_0_218 (.A(in3[54]), .B(in1[54]), .ZN(n_0_114));
   XNOR2_X1 i_0_219 (.A(in2[55]), .B(n_0_115), .ZN(sum[55]));
   XNOR2_X1 i_0_220 (.A(in3[55]), .B(in1[55]), .ZN(n_0_115));
   XNOR2_X1 i_0_221 (.A(in2[56]), .B(n_0_116), .ZN(sum[56]));
   XNOR2_X1 i_0_222 (.A(in3[56]), .B(in1[56]), .ZN(n_0_116));
   XNOR2_X1 i_0_223 (.A(in2[57]), .B(n_0_117), .ZN(sum[57]));
   XNOR2_X1 i_0_224 (.A(in3[57]), .B(in1[57]), .ZN(n_0_117));
   XNOR2_X1 i_0_225 (.A(in2[58]), .B(n_0_118), .ZN(sum[58]));
   XNOR2_X1 i_0_226 (.A(in3[58]), .B(in1[58]), .ZN(n_0_118));
   XNOR2_X1 i_0_227 (.A(in2[59]), .B(n_0_119), .ZN(sum[59]));
   XNOR2_X1 i_0_228 (.A(in3[59]), .B(in1[59]), .ZN(n_0_119));
   XNOR2_X1 i_0_229 (.A(in2[60]), .B(n_0_120), .ZN(sum[60]));
   XNOR2_X1 i_0_230 (.A(in3[60]), .B(in1[60]), .ZN(n_0_120));
   XNOR2_X1 i_0_231 (.A(in2[61]), .B(n_0_121), .ZN(sum[61]));
   XNOR2_X1 i_0_232 (.A(in3[61]), .B(in1[61]), .ZN(n_0_121));
   XNOR2_X1 i_0_233 (.A(in2[62]), .B(n_0_122), .ZN(sum[62]));
   XNOR2_X1 i_0_234 (.A(in3[62]), .B(in1[62]), .ZN(n_0_122));
   XNOR2_X1 i_0_235 (.A(in2[63]), .B(n_0_123), .ZN(sum[63]));
   XNOR2_X1 i_0_236 (.A(in3[63]), .B(in1[63]), .ZN(n_0_123));
   INV_X1 i_0_203 (.A(in1[47]), .ZN(n_0_107));
   XNOR2_X1 i_0_204 (.A(in2[47]), .B(in3[47]), .ZN(n_0_108));
   INV_X1 i_0_205 (.A(n_0_108), .ZN(n_0_109));
   AOI22_X1 i_0_206 (.A1(n_0_107), .A2(n_0_108), .B1(in1[47]), .B2(n_0_109), 
      .ZN(sum[47]));
   OR2_X1 i_0_207 (.A1(in2[48]), .A2(in3[48]), .ZN(n_0_124));
   NAND2_X1 i_0_208 (.A1(in2[48]), .A2(in3[48]), .ZN(n_0_125));
   AND3_X1 i_0_237 (.A1(in1[48]), .A2(n_0_124), .A3(n_0_125), .ZN(n_0_126));
   AOI21_X1 i_0_238 (.A(in1[48]), .B1(n_0_124), .B2(n_0_125), .ZN(n_0_127));
   NOR2_X1 i_0_239 (.A1(n_0_126), .A2(n_0_127), .ZN(sum[48]));
   OR2_X1 i_0_240 (.A1(in2[49]), .A2(in3[49]), .ZN(n_0_128));
   NAND2_X1 i_0_241 (.A1(in2[49]), .A2(in3[49]), .ZN(n_0_129));
   AND3_X1 i_0_242 (.A1(in1[49]), .A2(n_0_128), .A3(n_0_129), .ZN(n_0_130));
   AOI21_X1 i_0_243 (.A(in1[49]), .B1(n_0_128), .B2(n_0_129), .ZN(n_0_131));
   NOR2_X1 i_0_244 (.A1(n_0_130), .A2(n_0_131), .ZN(sum[49]));
endmodule

module CSA__4_20(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;

   AND2_X1 i_0_0 (.A1(in2[8]), .A2(in1[8]), .ZN(c[9]));
   AND2_X1 i_0_1 (.A1(in2[9]), .A2(in1[9]), .ZN(c[10]));
   AND2_X1 i_0_2 (.A1(in2[10]), .A2(in1[10]), .ZN(c[11]));
   AND2_X1 i_0_3 (.A1(in2[11]), .A2(in1[11]), .ZN(c[12]));
   AND2_X1 i_0_4 (.A1(in2[12]), .A2(in1[12]), .ZN(c[13]));
   AND2_X1 i_0_5 (.A1(in2[13]), .A2(in1[13]), .ZN(c[14]));
   AND2_X1 i_0_6 (.A1(in2[14]), .A2(in1[14]), .ZN(c[15]));
   AND2_X1 i_0_7 (.A1(in2[15]), .A2(in1[15]), .ZN(c[16]));
   AND2_X1 i_0_8 (.A1(in2[16]), .A2(in1[16]), .ZN(c[17]));
   AND2_X1 i_0_9 (.A1(in2[17]), .A2(in1[17]), .ZN(c[18]));
   AND2_X1 i_0_10 (.A1(in2[18]), .A2(in1[18]), .ZN(c[19]));
   AND2_X1 i_0_11 (.A1(in2[19]), .A2(in1[19]), .ZN(c[20]));
   AND2_X1 i_0_12 (.A1(in2[20]), .A2(in1[20]), .ZN(c[21]));
   AND2_X1 i_0_13 (.A1(in2[21]), .A2(in1[21]), .ZN(c[22]));
   AND2_X1 i_0_14 (.A1(in2[22]), .A2(in1[22]), .ZN(c[23]));
   AND2_X1 i_0_15 (.A1(in2[23]), .A2(in1[23]), .ZN(c[24]));
   AND2_X1 i_0_16 (.A1(in2[24]), .A2(in1[24]), .ZN(c[25]));
   AND2_X1 i_0_17 (.A1(in2[25]), .A2(in1[25]), .ZN(c[26]));
   AND2_X1 i_0_18 (.A1(in2[26]), .A2(in1[26]), .ZN(c[27]));
   AND2_X1 i_0_19 (.A1(in2[27]), .A2(in1[27]), .ZN(c[28]));
   AND2_X1 i_0_20 (.A1(in2[28]), .A2(in1[28]), .ZN(c[29]));
   AND2_X1 i_0_21 (.A1(in2[29]), .A2(in1[29]), .ZN(c[30]));
   AND2_X1 i_0_22 (.A1(in2[30]), .A2(in1[30]), .ZN(c[31]));
   NAND2_X1 i_0_23 (.A1(n_0_1), .A2(n_0_0), .ZN(c[32]));
   OAI21_X1 i_0_24 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_0));
   NAND2_X1 i_0_25 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_1));
   NAND2_X1 i_0_26 (.A1(n_0_3), .A2(n_0_2), .ZN(c[33]));
   OAI21_X1 i_0_27 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_2));
   NAND2_X1 i_0_28 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_3));
   NAND2_X1 i_0_29 (.A1(n_0_5), .A2(n_0_4), .ZN(c[34]));
   OAI21_X1 i_0_30 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_4));
   NAND2_X1 i_0_31 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_5));
   NAND2_X1 i_0_32 (.A1(n_0_7), .A2(n_0_6), .ZN(c[35]));
   OAI21_X1 i_0_33 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_6));
   NAND2_X1 i_0_34 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_7));
   NAND2_X1 i_0_35 (.A1(n_0_9), .A2(n_0_8), .ZN(c[36]));
   OAI21_X1 i_0_36 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_8));
   NAND2_X1 i_0_37 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_9));
   NAND2_X1 i_0_38 (.A1(n_0_11), .A2(n_0_10), .ZN(c[37]));
   OAI21_X1 i_0_39 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_10));
   NAND2_X1 i_0_40 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_11));
   NAND2_X1 i_0_41 (.A1(n_0_13), .A2(n_0_12), .ZN(c[38]));
   OAI21_X1 i_0_42 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_12));
   NAND2_X1 i_0_43 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_13));
   NAND2_X1 i_0_44 (.A1(n_0_15), .A2(n_0_14), .ZN(c[39]));
   OAI21_X1 i_0_45 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_14));
   NAND2_X1 i_0_46 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_15));
   NAND2_X1 i_0_47 (.A1(n_0_17), .A2(n_0_16), .ZN(c[40]));
   OAI21_X1 i_0_48 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_16));
   NAND2_X1 i_0_49 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_17));
   NAND2_X1 i_0_50 (.A1(n_0_19), .A2(n_0_18), .ZN(c[41]));
   OAI21_X1 i_0_51 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_18));
   NAND2_X1 i_0_52 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_19));
   NAND2_X1 i_0_53 (.A1(n_0_21), .A2(n_0_20), .ZN(c[42]));
   OAI21_X1 i_0_54 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_20));
   NAND2_X1 i_0_55 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_21));
   NAND2_X1 i_0_56 (.A1(n_0_23), .A2(n_0_22), .ZN(c[43]));
   OAI21_X1 i_0_57 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_22));
   NAND2_X1 i_0_58 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_23));
   NAND2_X1 i_0_59 (.A1(n_0_25), .A2(n_0_24), .ZN(c[44]));
   OAI21_X1 i_0_60 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_24));
   NAND2_X1 i_0_61 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_25));
   NAND2_X1 i_0_62 (.A1(n_0_27), .A2(n_0_26), .ZN(c[45]));
   OAI21_X1 i_0_63 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_26));
   NAND2_X1 i_0_64 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_27));
   NAND2_X1 i_0_65 (.A1(n_0_29), .A2(n_0_28), .ZN(c[46]));
   OAI21_X1 i_0_66 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_28));
   NAND2_X1 i_0_67 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_29));
   NAND2_X1 i_0_68 (.A1(n_0_31), .A2(n_0_30), .ZN(c[47]));
   OAI21_X1 i_0_69 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_30));
   NAND2_X1 i_0_70 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_31));
   NAND2_X1 i_0_71 (.A1(n_0_33), .A2(n_0_32), .ZN(c[48]));
   OAI21_X1 i_0_72 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_32));
   NAND2_X1 i_0_73 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_33));
   NAND2_X1 i_0_74 (.A1(n_0_35), .A2(n_0_34), .ZN(c[49]));
   OAI21_X1 i_0_75 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_34));
   NAND2_X1 i_0_76 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_35));
   NAND2_X1 i_0_77 (.A1(n_0_37), .A2(n_0_36), .ZN(c[50]));
   OAI21_X1 i_0_78 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_36));
   NAND2_X1 i_0_79 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_37));
   NAND2_X1 i_0_80 (.A1(n_0_39), .A2(n_0_38), .ZN(c[51]));
   OAI21_X1 i_0_81 (.A(in3[50]), .B1(in1[50]), .B2(in2[50]), .ZN(n_0_38));
   NAND2_X1 i_0_82 (.A1(in2[50]), .A2(in1[50]), .ZN(n_0_39));
   NAND2_X1 i_0_83 (.A1(n_0_41), .A2(n_0_40), .ZN(c[52]));
   OAI21_X1 i_0_84 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_40));
   NAND2_X1 i_0_85 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_41));
   NAND2_X1 i_0_86 (.A1(n_0_43), .A2(n_0_42), .ZN(c[53]));
   OAI21_X1 i_0_87 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_42));
   NAND2_X1 i_0_88 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_43));
   NAND2_X1 i_0_89 (.A1(n_0_45), .A2(n_0_44), .ZN(c[54]));
   OAI21_X1 i_0_90 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_44));
   NAND2_X1 i_0_91 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_45));
   NAND2_X1 i_0_92 (.A1(n_0_47), .A2(n_0_46), .ZN(c[55]));
   OAI21_X1 i_0_93 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_46));
   NAND2_X1 i_0_94 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_47));
   NAND2_X1 i_0_95 (.A1(n_0_49), .A2(n_0_48), .ZN(c[56]));
   OAI21_X1 i_0_96 (.A(in2[55]), .B1(in3[55]), .B2(in1[55]), .ZN(n_0_48));
   NAND2_X1 i_0_97 (.A1(in3[55]), .A2(in1[55]), .ZN(n_0_49));
   NAND2_X1 i_0_98 (.A1(n_0_51), .A2(n_0_50), .ZN(c[57]));
   OAI21_X1 i_0_99 (.A(in2[56]), .B1(in3[56]), .B2(in1[56]), .ZN(n_0_50));
   NAND2_X1 i_0_100 (.A1(in3[56]), .A2(in1[56]), .ZN(n_0_51));
   NAND2_X1 i_0_101 (.A1(n_0_53), .A2(n_0_52), .ZN(c[58]));
   OAI21_X1 i_0_102 (.A(in2[57]), .B1(in3[57]), .B2(in1[57]), .ZN(n_0_52));
   NAND2_X1 i_0_103 (.A1(in3[57]), .A2(in1[57]), .ZN(n_0_53));
   NAND2_X1 i_0_104 (.A1(n_0_55), .A2(n_0_54), .ZN(c[59]));
   OAI21_X1 i_0_105 (.A(in2[58]), .B1(in3[58]), .B2(in1[58]), .ZN(n_0_54));
   NAND2_X1 i_0_106 (.A1(in3[58]), .A2(in1[58]), .ZN(n_0_55));
   NAND2_X1 i_0_107 (.A1(n_0_57), .A2(n_0_56), .ZN(c[60]));
   OAI21_X1 i_0_108 (.A(in2[59]), .B1(in3[59]), .B2(in1[59]), .ZN(n_0_56));
   NAND2_X1 i_0_109 (.A1(in3[59]), .A2(in1[59]), .ZN(n_0_57));
   NAND2_X1 i_0_110 (.A1(n_0_59), .A2(n_0_58), .ZN(c[61]));
   OAI21_X1 i_0_111 (.A(in2[60]), .B1(in3[60]), .B2(in1[60]), .ZN(n_0_58));
   NAND2_X1 i_0_112 (.A1(in3[60]), .A2(in1[60]), .ZN(n_0_59));
   NAND2_X1 i_0_113 (.A1(n_0_61), .A2(n_0_60), .ZN(c[62]));
   OAI21_X1 i_0_114 (.A(in2[61]), .B1(in3[61]), .B2(in1[61]), .ZN(n_0_60));
   NAND2_X1 i_0_115 (.A1(in3[61]), .A2(in1[61]), .ZN(n_0_61));
   NAND2_X1 i_0_116 (.A1(n_0_63), .A2(n_0_62), .ZN(c[63]));
   OAI21_X1 i_0_117 (.A(in2[62]), .B1(in3[62]), .B2(in1[62]), .ZN(n_0_62));
   NAND2_X1 i_0_118 (.A1(in3[62]), .A2(in1[62]), .ZN(n_0_63));
   XOR2_X1 i_0_119 (.A(in2[8]), .B(in1[8]), .Z(sum[8]));
   XOR2_X1 i_0_120 (.A(in2[9]), .B(in1[9]), .Z(sum[9]));
   XOR2_X1 i_0_121 (.A(in2[10]), .B(in1[10]), .Z(sum[10]));
   XOR2_X1 i_0_122 (.A(in2[11]), .B(in1[11]), .Z(sum[11]));
   XOR2_X1 i_0_123 (.A(in2[12]), .B(in1[12]), .Z(sum[12]));
   XOR2_X1 i_0_124 (.A(in2[13]), .B(in1[13]), .Z(sum[13]));
   XOR2_X1 i_0_125 (.A(in2[14]), .B(in1[14]), .Z(sum[14]));
   XOR2_X1 i_0_126 (.A(in2[15]), .B(in1[15]), .Z(sum[15]));
   XOR2_X1 i_0_127 (.A(in2[16]), .B(in1[16]), .Z(sum[16]));
   XOR2_X1 i_0_128 (.A(in2[17]), .B(in1[17]), .Z(sum[17]));
   XOR2_X1 i_0_129 (.A(in2[18]), .B(in1[18]), .Z(sum[18]));
   XOR2_X1 i_0_130 (.A(in2[19]), .B(in1[19]), .Z(sum[19]));
   XOR2_X1 i_0_131 (.A(in2[20]), .B(in1[20]), .Z(sum[20]));
   XOR2_X1 i_0_132 (.A(in2[21]), .B(in1[21]), .Z(sum[21]));
   XOR2_X1 i_0_133 (.A(in2[22]), .B(in1[22]), .Z(sum[22]));
   XOR2_X1 i_0_134 (.A(in2[23]), .B(in1[23]), .Z(sum[23]));
   XOR2_X1 i_0_135 (.A(in2[24]), .B(in1[24]), .Z(sum[24]));
   XOR2_X1 i_0_136 (.A(in2[25]), .B(in1[25]), .Z(sum[25]));
   XOR2_X1 i_0_137 (.A(in2[26]), .B(in1[26]), .Z(sum[26]));
   XOR2_X1 i_0_138 (.A(in2[27]), .B(in1[27]), .Z(sum[27]));
   XOR2_X1 i_0_139 (.A(in2[28]), .B(in1[28]), .Z(sum[28]));
   XOR2_X1 i_0_140 (.A(in2[29]), .B(in1[29]), .Z(sum[29]));
   XOR2_X1 i_0_141 (.A(in2[30]), .B(in1[30]), .Z(sum[30]));
   XNOR2_X1 i_0_142 (.A(in2[31]), .B(n_0_64), .ZN(sum[31]));
   XNOR2_X1 i_0_143 (.A(in3[31]), .B(in1[31]), .ZN(n_0_64));
   XNOR2_X1 i_0_144 (.A(in2[32]), .B(n_0_65), .ZN(sum[32]));
   XNOR2_X1 i_0_145 (.A(in3[32]), .B(in1[32]), .ZN(n_0_65));
   XNOR2_X1 i_0_146 (.A(in2[33]), .B(n_0_66), .ZN(sum[33]));
   XNOR2_X1 i_0_147 (.A(in3[33]), .B(in1[33]), .ZN(n_0_66));
   XNOR2_X1 i_0_148 (.A(in2[34]), .B(n_0_67), .ZN(sum[34]));
   XNOR2_X1 i_0_149 (.A(in3[34]), .B(in1[34]), .ZN(n_0_67));
   XNOR2_X1 i_0_150 (.A(in2[35]), .B(n_0_68), .ZN(sum[35]));
   XNOR2_X1 i_0_151 (.A(in3[35]), .B(in1[35]), .ZN(n_0_68));
   XNOR2_X1 i_0_152 (.A(in2[36]), .B(n_0_69), .ZN(sum[36]));
   XNOR2_X1 i_0_153 (.A(in3[36]), .B(in1[36]), .ZN(n_0_69));
   XNOR2_X1 i_0_154 (.A(in2[37]), .B(n_0_70), .ZN(sum[37]));
   XNOR2_X1 i_0_155 (.A(in3[37]), .B(in1[37]), .ZN(n_0_70));
   XNOR2_X1 i_0_156 (.A(in2[38]), .B(n_0_71), .ZN(sum[38]));
   XNOR2_X1 i_0_157 (.A(in3[38]), .B(in1[38]), .ZN(n_0_71));
   XNOR2_X1 i_0_158 (.A(in2[39]), .B(n_0_72), .ZN(sum[39]));
   XNOR2_X1 i_0_159 (.A(in3[39]), .B(in1[39]), .ZN(n_0_72));
   XNOR2_X1 i_0_160 (.A(in2[40]), .B(n_0_73), .ZN(sum[40]));
   XNOR2_X1 i_0_161 (.A(in3[40]), .B(in1[40]), .ZN(n_0_73));
   XNOR2_X1 i_0_162 (.A(in2[41]), .B(n_0_74), .ZN(sum[41]));
   XNOR2_X1 i_0_163 (.A(in3[41]), .B(in1[41]), .ZN(n_0_74));
   XNOR2_X1 i_0_164 (.A(in2[42]), .B(n_0_75), .ZN(sum[42]));
   XNOR2_X1 i_0_165 (.A(in3[42]), .B(in1[42]), .ZN(n_0_75));
   XNOR2_X1 i_0_166 (.A(in2[43]), .B(n_0_76), .ZN(sum[43]));
   XNOR2_X1 i_0_167 (.A(in3[43]), .B(in1[43]), .ZN(n_0_76));
   XNOR2_X1 i_0_168 (.A(in2[44]), .B(n_0_77), .ZN(sum[44]));
   XNOR2_X1 i_0_169 (.A(in3[44]), .B(in1[44]), .ZN(n_0_77));
   XNOR2_X1 i_0_170 (.A(in2[45]), .B(n_0_78), .ZN(sum[45]));
   XNOR2_X1 i_0_171 (.A(in3[45]), .B(in1[45]), .ZN(n_0_78));
   XNOR2_X1 i_0_172 (.A(in2[46]), .B(n_0_79), .ZN(sum[46]));
   XNOR2_X1 i_0_173 (.A(in3[46]), .B(in1[46]), .ZN(n_0_79));
   XNOR2_X1 i_0_180 (.A(in2[50]), .B(n_0_83), .ZN(sum[50]));
   XNOR2_X1 i_0_181 (.A(in3[50]), .B(in1[50]), .ZN(n_0_83));
   XNOR2_X1 i_0_182 (.A(in2[51]), .B(n_0_84), .ZN(sum[51]));
   XNOR2_X1 i_0_183 (.A(in3[51]), .B(in1[51]), .ZN(n_0_84));
   XNOR2_X1 i_0_184 (.A(in2[52]), .B(n_0_85), .ZN(sum[52]));
   XNOR2_X1 i_0_185 (.A(in3[52]), .B(in1[52]), .ZN(n_0_85));
   XNOR2_X1 i_0_186 (.A(in2[53]), .B(n_0_86), .ZN(sum[53]));
   XNOR2_X1 i_0_187 (.A(in3[53]), .B(in1[53]), .ZN(n_0_86));
   XNOR2_X1 i_0_188 (.A(in2[54]), .B(n_0_87), .ZN(sum[54]));
   XNOR2_X1 i_0_189 (.A(in3[54]), .B(in1[54]), .ZN(n_0_87));
   XNOR2_X1 i_0_190 (.A(in2[55]), .B(n_0_88), .ZN(sum[55]));
   XNOR2_X1 i_0_191 (.A(in3[55]), .B(in1[55]), .ZN(n_0_88));
   XNOR2_X1 i_0_192 (.A(in2[56]), .B(n_0_89), .ZN(sum[56]));
   XNOR2_X1 i_0_193 (.A(in3[56]), .B(in1[56]), .ZN(n_0_89));
   XNOR2_X1 i_0_194 (.A(in2[57]), .B(n_0_90), .ZN(sum[57]));
   XNOR2_X1 i_0_195 (.A(in3[57]), .B(in1[57]), .ZN(n_0_90));
   XNOR2_X1 i_0_196 (.A(in2[58]), .B(n_0_91), .ZN(sum[58]));
   XNOR2_X1 i_0_197 (.A(in3[58]), .B(in1[58]), .ZN(n_0_91));
   XNOR2_X1 i_0_198 (.A(in2[59]), .B(n_0_92), .ZN(sum[59]));
   XNOR2_X1 i_0_199 (.A(in3[59]), .B(in1[59]), .ZN(n_0_92));
   XNOR2_X1 i_0_200 (.A(in2[60]), .B(n_0_93), .ZN(sum[60]));
   XNOR2_X1 i_0_201 (.A(in3[60]), .B(in1[60]), .ZN(n_0_93));
   XNOR2_X1 i_0_202 (.A(in2[61]), .B(n_0_94), .ZN(sum[61]));
   XNOR2_X1 i_0_203 (.A(in3[61]), .B(in1[61]), .ZN(n_0_94));
   XNOR2_X1 i_0_204 (.A(in2[62]), .B(n_0_95), .ZN(sum[62]));
   XNOR2_X1 i_0_205 (.A(in3[62]), .B(in1[62]), .ZN(n_0_95));
   XNOR2_X1 i_0_206 (.A(in2[63]), .B(n_0_96), .ZN(sum[63]));
   XNOR2_X1 i_0_207 (.A(in3[63]), .B(in1[63]), .ZN(n_0_96));
   XNOR2_X1 i_0_174 (.A(in2[47]), .B(in3[47]), .ZN(n_0_80));
   XNOR2_X1 i_0_175 (.A(in1[47]), .B(n_0_80), .ZN(sum[47]));
   XOR2_X1 i_0_176 (.A(in2[48]), .B(n_0_81), .Z(sum[48]));
   XOR2_X1 i_0_177 (.A(in3[48]), .B(in1[48]), .Z(n_0_81));
   XOR2_X1 i_0_178 (.A(in2[49]), .B(n_0_82), .Z(sum[49]));
   XOR2_X1 i_0_179 (.A(in3[49]), .B(in1[49]), .Z(n_0_82));
endmodule

module CSA__4_23(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   AND2_X1 i_0_0 (.A1(in2[9]), .A2(in1[9]), .ZN(c[10]));
   AND2_X1 i_0_1 (.A1(in2[10]), .A2(in1[10]), .ZN(c[11]));
   AND2_X1 i_0_2 (.A1(in2[11]), .A2(in1[11]), .ZN(c[12]));
   AND2_X1 i_0_3 (.A1(in2[12]), .A2(in1[12]), .ZN(c[13]));
   AND2_X1 i_0_4 (.A1(in2[13]), .A2(in1[13]), .ZN(c[14]));
   AND2_X1 i_0_5 (.A1(in2[14]), .A2(in1[14]), .ZN(c[15]));
   AND2_X1 i_0_6 (.A1(in2[15]), .A2(in1[15]), .ZN(c[16]));
   AND2_X1 i_0_7 (.A1(in2[16]), .A2(in1[16]), .ZN(c[17]));
   AND2_X1 i_0_8 (.A1(in2[17]), .A2(in1[17]), .ZN(c[18]));
   AND2_X1 i_0_9 (.A1(in2[18]), .A2(in1[18]), .ZN(c[19]));
   AND2_X1 i_0_10 (.A1(in2[19]), .A2(in1[19]), .ZN(c[20]));
   AND2_X1 i_0_11 (.A1(in2[20]), .A2(in1[20]), .ZN(c[21]));
   AND2_X1 i_0_12 (.A1(in2[21]), .A2(in1[21]), .ZN(c[22]));
   AND2_X1 i_0_13 (.A1(in2[22]), .A2(in1[22]), .ZN(c[23]));
   AND2_X1 i_0_14 (.A1(in2[23]), .A2(in1[23]), .ZN(c[24]));
   AND2_X1 i_0_15 (.A1(in2[24]), .A2(in1[24]), .ZN(c[25]));
   AND2_X1 i_0_16 (.A1(in2[25]), .A2(in1[25]), .ZN(c[26]));
   AND2_X1 i_0_17 (.A1(in2[26]), .A2(in1[26]), .ZN(c[27]));
   AND2_X1 i_0_18 (.A1(in2[27]), .A2(in1[27]), .ZN(c[28]));
   AND2_X1 i_0_19 (.A1(in2[28]), .A2(in1[28]), .ZN(c[29]));
   AND2_X1 i_0_20 (.A1(in2[29]), .A2(in1[29]), .ZN(c[30]));
   AND2_X1 i_0_21 (.A1(in2[30]), .A2(in1[30]), .ZN(c[31]));
   NAND2_X1 i_0_22 (.A1(n_0_1), .A2(n_0_0), .ZN(c[32]));
   OAI21_X1 i_0_23 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_0));
   NAND2_X1 i_0_24 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_1));
   AND2_X1 i_0_25 (.A1(in2[32]), .A2(in1[32]), .ZN(c[33]));
   AND2_X1 i_0_26 (.A1(in2[33]), .A2(in1[33]), .ZN(c[34]));
   AND2_X1 i_0_27 (.A1(in2[34]), .A2(in1[34]), .ZN(c[35]));
   AND2_X1 i_0_28 (.A1(in2[35]), .A2(in1[35]), .ZN(c[36]));
   AND2_X1 i_0_29 (.A1(in2[36]), .A2(in1[36]), .ZN(c[37]));
   AND2_X1 i_0_30 (.A1(in2[37]), .A2(in1[37]), .ZN(c[38]));
   AND2_X1 i_0_31 (.A1(in2[38]), .A2(in1[38]), .ZN(c[39]));
   AND2_X1 i_0_32 (.A1(in2[39]), .A2(in1[39]), .ZN(c[40]));
   AND2_X1 i_0_33 (.A1(in2[40]), .A2(in1[40]), .ZN(c[41]));
   AND2_X1 i_0_34 (.A1(in2[41]), .A2(in1[41]), .ZN(c[42]));
   AND2_X1 i_0_35 (.A1(in2[42]), .A2(in1[42]), .ZN(c[43]));
   AND2_X1 i_0_36 (.A1(in2[43]), .A2(in1[43]), .ZN(c[44]));
   AND2_X1 i_0_37 (.A1(in2[44]), .A2(in1[44]), .ZN(c[45]));
   AND2_X1 i_0_38 (.A1(in2[45]), .A2(in1[45]), .ZN(c[46]));
   AND2_X1 i_0_39 (.A1(in2[46]), .A2(in1[46]), .ZN(c[47]));
   AND2_X1 i_0_40 (.A1(in2[47]), .A2(in1[47]), .ZN(c[48]));
   AND2_X1 i_0_41 (.A1(in2[48]), .A2(in1[48]), .ZN(c[49]));
   AND2_X1 i_0_42 (.A1(in2[49]), .A2(in1[49]), .ZN(c[50]));
   AND2_X1 i_0_43 (.A1(in2[50]), .A2(in1[50]), .ZN(c[51]));
   AND2_X1 i_0_44 (.A1(in2[51]), .A2(in1[51]), .ZN(c[52]));
   AND2_X1 i_0_45 (.A1(in2[52]), .A2(in1[52]), .ZN(c[53]));
   AND2_X1 i_0_46 (.A1(in2[53]), .A2(in1[53]), .ZN(c[54]));
   AND2_X1 i_0_47 (.A1(in2[54]), .A2(in1[54]), .ZN(c[55]));
   AND2_X1 i_0_48 (.A1(in2[55]), .A2(in1[55]), .ZN(c[56]));
   AND2_X1 i_0_49 (.A1(in2[56]), .A2(in1[56]), .ZN(c[57]));
   AND2_X1 i_0_50 (.A1(in2[57]), .A2(in1[57]), .ZN(c[58]));
   AND2_X1 i_0_51 (.A1(in2[58]), .A2(in1[58]), .ZN(c[59]));
   AND2_X1 i_0_52 (.A1(in2[59]), .A2(in1[59]), .ZN(c[60]));
   AND2_X1 i_0_53 (.A1(in2[60]), .A2(in1[60]), .ZN(c[61]));
   AND2_X1 i_0_54 (.A1(in2[61]), .A2(in1[61]), .ZN(c[62]));
   AND2_X1 i_0_55 (.A1(in2[62]), .A2(in1[62]), .ZN(c[63]));
   XOR2_X1 i_0_56 (.A(in2[9]), .B(in1[9]), .Z(sum[9]));
   XOR2_X1 i_0_57 (.A(in2[10]), .B(in1[10]), .Z(sum[10]));
   XOR2_X1 i_0_58 (.A(in2[11]), .B(in1[11]), .Z(sum[11]));
   XOR2_X1 i_0_59 (.A(in2[12]), .B(in1[12]), .Z(sum[12]));
   XOR2_X1 i_0_60 (.A(in2[13]), .B(in1[13]), .Z(sum[13]));
   XOR2_X1 i_0_61 (.A(in2[14]), .B(in1[14]), .Z(sum[14]));
   XOR2_X1 i_0_62 (.A(in2[15]), .B(in1[15]), .Z(sum[15]));
   XOR2_X1 i_0_63 (.A(in2[16]), .B(in1[16]), .Z(sum[16]));
   XOR2_X1 i_0_64 (.A(in2[17]), .B(in1[17]), .Z(sum[17]));
   XOR2_X1 i_0_65 (.A(in2[18]), .B(in1[18]), .Z(sum[18]));
   XOR2_X1 i_0_66 (.A(in2[19]), .B(in1[19]), .Z(sum[19]));
   XOR2_X1 i_0_67 (.A(in2[20]), .B(in1[20]), .Z(sum[20]));
   XOR2_X1 i_0_68 (.A(in2[21]), .B(in1[21]), .Z(sum[21]));
   XOR2_X1 i_0_69 (.A(in2[22]), .B(in1[22]), .Z(sum[22]));
   XOR2_X1 i_0_70 (.A(in2[23]), .B(in1[23]), .Z(sum[23]));
   XOR2_X1 i_0_71 (.A(in2[24]), .B(in1[24]), .Z(sum[24]));
   XOR2_X1 i_0_72 (.A(in2[25]), .B(in1[25]), .Z(sum[25]));
   XOR2_X1 i_0_73 (.A(in2[26]), .B(in1[26]), .Z(sum[26]));
   XOR2_X1 i_0_74 (.A(in2[27]), .B(in1[27]), .Z(sum[27]));
   XOR2_X1 i_0_75 (.A(in2[28]), .B(in1[28]), .Z(sum[28]));
   XOR2_X1 i_0_76 (.A(in2[29]), .B(in1[29]), .Z(sum[29]));
   XOR2_X1 i_0_77 (.A(in2[30]), .B(in1[30]), .Z(sum[30]));
   XNOR2_X1 i_0_78 (.A(in2[31]), .B(n_0_2), .ZN(sum[31]));
   XNOR2_X1 i_0_79 (.A(in3[31]), .B(in1[31]), .ZN(n_0_2));
   XOR2_X1 i_0_80 (.A(in2[32]), .B(in1[32]), .Z(sum[32]));
   XOR2_X1 i_0_81 (.A(in2[33]), .B(in1[33]), .Z(sum[33]));
   XOR2_X1 i_0_82 (.A(in2[34]), .B(in1[34]), .Z(sum[34]));
   XOR2_X1 i_0_83 (.A(in2[35]), .B(in1[35]), .Z(sum[35]));
   XOR2_X1 i_0_84 (.A(in2[36]), .B(in1[36]), .Z(sum[36]));
   XOR2_X1 i_0_85 (.A(in2[37]), .B(in1[37]), .Z(sum[37]));
   XOR2_X1 i_0_86 (.A(in2[38]), .B(in1[38]), .Z(sum[38]));
   XOR2_X1 i_0_87 (.A(in2[39]), .B(in1[39]), .Z(sum[39]));
   XOR2_X1 i_0_88 (.A(in2[40]), .B(in1[40]), .Z(sum[40]));
   XOR2_X1 i_0_89 (.A(in2[41]), .B(in1[41]), .Z(sum[41]));
   XOR2_X1 i_0_90 (.A(in2[42]), .B(in1[42]), .Z(sum[42]));
   XOR2_X1 i_0_91 (.A(in2[43]), .B(in1[43]), .Z(sum[43]));
   XOR2_X1 i_0_92 (.A(in2[44]), .B(in1[44]), .Z(sum[44]));
   XOR2_X1 i_0_93 (.A(in2[45]), .B(in1[45]), .Z(sum[45]));
   XOR2_X1 i_0_94 (.A(in2[46]), .B(in1[46]), .Z(sum[46]));
   XOR2_X1 i_0_95 (.A(in2[47]), .B(in1[47]), .Z(sum[47]));
   XOR2_X1 i_0_96 (.A(in2[48]), .B(in1[48]), .Z(sum[48]));
   XOR2_X1 i_0_97 (.A(in2[49]), .B(in1[49]), .Z(sum[49]));
   XOR2_X1 i_0_98 (.A(in2[50]), .B(in1[50]), .Z(sum[50]));
   XOR2_X1 i_0_99 (.A(in2[51]), .B(in1[51]), .Z(sum[51]));
   XOR2_X1 i_0_100 (.A(in2[52]), .B(in1[52]), .Z(sum[52]));
   XOR2_X1 i_0_101 (.A(in2[53]), .B(in1[53]), .Z(sum[53]));
   XOR2_X1 i_0_102 (.A(in2[54]), .B(in1[54]), .Z(sum[54]));
   XOR2_X1 i_0_103 (.A(in2[55]), .B(in1[55]), .Z(sum[55]));
   XOR2_X1 i_0_104 (.A(in2[56]), .B(in1[56]), .Z(sum[56]));
   XOR2_X1 i_0_105 (.A(in2[57]), .B(in1[57]), .Z(sum[57]));
   XOR2_X1 i_0_106 (.A(in2[58]), .B(in1[58]), .Z(sum[58]));
   XOR2_X1 i_0_107 (.A(in2[59]), .B(in1[59]), .Z(sum[59]));
   XOR2_X1 i_0_108 (.A(in2[60]), .B(in1[60]), .Z(sum[60]));
   XOR2_X1 i_0_109 (.A(in2[61]), .B(in1[61]), .Z(sum[61]));
   XOR2_X1 i_0_110 (.A(in2[62]), .B(in1[62]), .Z(sum[62]));
   XOR2_X1 i_0_111 (.A(in2[63]), .B(in1[63]), .Z(sum[63]));
endmodule

module datapath(b, cin, a, sum);
   input [63:0]b;
   input cin;
   input [63:0]a;
   output [63:0]sum;

   INV_X1 i_0 (.A(n_0), .ZN(sum[10]));
   OAI21_X1 i_1 (.A(n_274), .B1(b[10]), .B2(a[10]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_274), .B(n_1), .Z(sum[11]));
   OAI21_X1 i_3 (.A(n_273), .B1(b[11]), .B2(a[11]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_272), .B(n_2), .ZN(sum[12]));
   OAI21_X1 i_5 (.A(n_276), .B1(b[12]), .B2(a[12]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_270), .B(n_3), .Z(sum[13]));
   XOR2_X1 i_7 (.A(b[13]), .B(a[13]), .Z(n_3));
   XOR2_X1 i_8 (.A(n_269), .B(n_10), .Z(sum[14]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(sum[15]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(sum[16]));
   NOR2_X1 i_11 (.A1(n_266), .A2(n_257), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(sum[17]));
   OAI22_X1 i_13 (.A1(b[16]), .A2(a[16]), .B1(n_257), .B2(n_7), .ZN(n_5));
   AOI21_X1 i_14 (.A(n_267), .B1(b[15]), .B2(a[15]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_267), .B1(n_261), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_264), .B1(n_269), .B2(n_262), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_262), .B1(b[14]), .B2(a[14]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_268), .A2(n_259), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_255), .B(n_18), .ZN(sum[18]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(sum[19]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(sum[20]));
   NOR2_X1 i_23 (.A1(n_252), .A2(n_243), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(sum[21]));
   OAI22_X1 i_25 (.A1(b[20]), .A2(a[20]), .B1(n_243), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_253), .B1(b[19]), .B2(a[19]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_253), .B1(n_247), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_250), .B1(n_255), .B2(n_248), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_250), .B1(b[18]), .B2(a[18]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_254), .A2(n_113), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_160), .B(n_26), .Z(sum[22]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(sum[23]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(sum[24]));
   NOR2_X1 i_35 (.A1(n_109), .A2(n_229), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(sum[25]));
   OAI22_X1 i_37 (.A1(b[24]), .A2(a[24]), .B1(n_229), .B2(n_23), .ZN(n_21));
   AOI21_X1 i_38 (.A(n_111), .B1(b[23]), .B2(a[23]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_111), .B1(n_162), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_161), .B1(n_160), .B2(n_163), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_163), .B1(b[22]), .B2(a[22]), .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_165), .A2(n_166), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_155), .B(n_34), .Z(sum[26]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(sum[27]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(sum[28]));
   NOR2_X1 i_47 (.A1(n_196), .A2(n_189), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(sum[29]));
   OAI21_X1 i_49 (.A(n_96), .B1(n_189), .B2(n_31), .ZN(n_29));
   NOR2_X1 i_50 (.A1(n_198), .A2(n_188), .ZN(n_30));
   INV_X1 i_51 (.A(n_32), .ZN(n_31));
   OAI21_X1 i_52 (.A(n_97), .B1(n_188), .B2(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_169), .B1(n_155), .B2(n_193), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_193), .B1(b[26]), .B2(a[26]), .ZN(n_34));
   AOI21_X1 i_55 (.A(n_191), .B1(b[29]), .B2(a[29]), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_63), .B(n_42), .Z(sum[30]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(sum[31]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(sum[32]));
   NOR2_X1 i_59 (.A1(n_221), .A2(n_173), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(sum[33]));
   OAI21_X1 i_61 (.A(n_106), .B1(n_173), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_223), .A2(n_181), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_108), .B1(n_181), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_204), .B1(n_175), .B2(n_63), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_175), .B1(b[30]), .B2(a[30]), .ZN(n_42));
   AOI21_X1 i_67 (.A(n_203), .B1(b[33]), .B2(a[33]), .ZN(n_43));
   XOR2_X1 i_68 (.A(n_61), .B(n_50), .Z(sum[34]));
   XOR2_X1 i_69 (.A(n_49), .B(n_46), .Z(sum[35]));
   XOR2_X1 i_70 (.A(n_47), .B(n_44), .Z(sum[36]));
   NOR2_X1 i_71 (.A1(n_207), .A2(n_179), .ZN(n_44));
   XNOR2_X1 i_72 (.A(n_51), .B(n_45), .ZN(sum[37]));
   OAI21_X1 i_73 (.A(n_100), .B1(n_179), .B2(n_47), .ZN(n_45));
   NOR2_X1 i_74 (.A1(n_209), .A2(n_167), .ZN(n_46));
   INV_X1 i_75 (.A(n_48), .ZN(n_47));
   OAI21_X1 i_76 (.A(n_101), .B1(n_167), .B2(n_49), .ZN(n_48));
   AOI21_X1 i_77 (.A(n_98), .B1(n_182), .B2(n_61), .ZN(n_49));
   OAI21_X1 i_78 (.A(n_182), .B1(b[34]), .B2(a[34]), .ZN(n_50));
   AOI21_X1 i_79 (.A(n_199), .B1(b[37]), .B2(a[37]), .ZN(n_51));
   XNOR2_X1 i_80 (.A(n_60), .B(n_59), .ZN(sum[38]));
   XOR2_X1 i_81 (.A(n_57), .B(n_56), .Z(sum[39]));
   XNOR2_X1 i_82 (.A(n_53), .B(n_52), .ZN(sum[40]));
   OAI22_X1 i_83 (.A1(b[39]), .A2(a[39]), .B1(n_94), .B2(n_57), .ZN(n_52));
   NOR2_X1 i_84 (.A1(n_215), .A2(n_172), .ZN(n_53));
   XNOR2_X1 i_85 (.A(n_65), .B(n_54), .ZN(sum[41]));
   OAI21_X1 i_86 (.A(n_55), .B1(n_214), .B2(n_172), .ZN(n_54));
   NAND3_X1 i_87 (.A1(n_183), .A2(n_56), .A3(n_58), .ZN(n_55));
   NOR2_X1 i_88 (.A1(n_216), .A2(n_94), .ZN(n_56));
   INV_X1 i_89 (.A(n_58), .ZN(n_57));
   OAI22_X1 i_90 (.A1(b[38]), .A2(a[38]), .B1(n_95), .B2(n_60), .ZN(n_58));
   OAI21_X1 i_91 (.A(n_177), .B1(b[38]), .B2(a[38]), .ZN(n_59));
   OAI21_X1 i_92 (.A(n_176), .B1(n_194), .B2(n_61), .ZN(n_60));
   INV_X1 i_93 (.A(n_62), .ZN(n_61));
   OAI21_X1 i_94 (.A(n_170), .B1(n_200), .B2(n_63), .ZN(n_62));
   INV_X1 i_95 (.A(n_64), .ZN(n_63));
   OAI21_X1 i_96 (.A(n_185), .B1(n_155), .B2(n_168), .ZN(n_64));
   AOI21_X1 i_97 (.A(n_184), .B1(b[41]), .B2(a[41]), .ZN(n_65));
   XOR2_X1 i_98 (.A(n_144), .B(n_72), .Z(sum[42]));
   XOR2_X1 i_99 (.A(n_71), .B(n_68), .Z(sum[43]));
   XOR2_X1 i_100 (.A(n_69), .B(n_66), .Z(sum[44]));
   NOR2_X1 i_101 (.A1(n_139), .A2(n_125), .ZN(n_66));
   XOR2_X1 i_102 (.A(n_73), .B(n_67), .Z(sum[45]));
   OAI21_X1 i_103 (.A(n_138), .B1(n_125), .B2(n_69), .ZN(n_67));
   NOR2_X1 i_104 (.A1(n_137), .A2(n_131), .ZN(n_68));
   INV_X1 i_105 (.A(n_70), .ZN(n_69));
   OAI21_X1 i_106 (.A(n_136), .B1(n_131), .B2(n_71), .ZN(n_70));
   AOI21_X1 i_107 (.A(n_135), .B1(n_144), .B2(n_129), .ZN(n_71));
   OAI21_X1 i_108 (.A(n_129), .B1(b[42]), .B2(a[42]), .ZN(n_72));
   OAI21_X1 i_109 (.A(n_140), .B1(n_249), .B2(n_246), .ZN(n_73));
   XOR2_X1 i_110 (.A(n_124), .B(n_80), .Z(sum[46]));
   XOR2_X1 i_111 (.A(n_79), .B(n_76), .Z(sum[47]));
   XOR2_X1 i_112 (.A(n_77), .B(n_74), .Z(sum[48]));
   NOR2_X1 i_113 (.A1(n_117), .A2(n_141), .ZN(n_74));
   XNOR2_X1 i_114 (.A(n_81), .B(n_75), .ZN(sum[49]));
   OAI21_X1 i_115 (.A(n_245), .B1(n_141), .B2(n_77), .ZN(n_75));
   NOR2_X1 i_116 (.A1(n_116), .A2(n_143), .ZN(n_76));
   INV_X1 i_117 (.A(n_78), .ZN(n_77));
   OAI21_X1 i_118 (.A(n_242), .B1(n_143), .B2(n_79), .ZN(n_78));
   AOI21_X1 i_119 (.A(n_208), .B1(n_237), .B2(n_124), .ZN(n_79));
   OAI21_X1 i_120 (.A(n_237), .B1(b[46]), .B2(a[46]), .ZN(n_80));
   AOI21_X1 i_121 (.A(n_239), .B1(b[49]), .B2(a[49]), .ZN(n_81));
   XNOR2_X1 i_122 (.A(n_90), .B(n_89), .ZN(sum[50]));
   XOR2_X1 i_123 (.A(n_87), .B(n_86), .Z(sum[51]));
   XNOR2_X1 i_124 (.A(n_83), .B(n_82), .ZN(sum[52]));
   OAI22_X1 i_125 (.A1(b[51]), .A2(a[51]), .B1(n_222), .B2(n_87), .ZN(n_82));
   NOR2_X1 i_126 (.A1(n_227), .A2(n_147), .ZN(n_83));
   XNOR2_X1 i_127 (.A(n_91), .B(n_84), .ZN(sum[53]));
   OAI21_X1 i_128 (.A(n_85), .B1(n_282), .B2(n_147), .ZN(n_84));
   NAND3_X1 i_129 (.A1(n_220), .A2(n_86), .A3(n_88), .ZN(n_85));
   NOR2_X1 i_130 (.A1(n_226), .A2(n_222), .ZN(n_86));
   INV_X1 i_131 (.A(n_88), .ZN(n_87));
   OAI22_X1 i_132 (.A1(b[50]), .A2(a[50]), .B1(n_224), .B2(n_90), .ZN(n_88));
   OAI21_X1 i_133 (.A(n_225), .B1(b[50]), .B2(a[50]), .ZN(n_89));
   OAI21_X1 i_134 (.A(n_230), .B1(n_206), .B2(n_124), .ZN(n_90));
   AOI21_X1 i_135 (.A(n_228), .B1(b[53]), .B2(a[53]), .ZN(n_91));
   XNOR2_X1 i_136 (.A(n_123), .B(n_99), .ZN(sum[54]));
   XNOR2_X1 i_137 (.A(n_93), .B(n_92), .ZN(sum[56]));
   OAI22_X1 i_138 (.A1(b[55]), .A2(a[55]), .B1(n_119), .B2(n_121), .ZN(n_92));
   NOR2_X1 i_139 (.A1(n_280), .A2(n_281), .ZN(n_93));
   OAI21_X1 i_140 (.A(n_241), .B1(b[54]), .B2(a[54]), .ZN(n_99));
   XNOR2_X1 i_141 (.A(n_104), .B(n_103), .ZN(sum[60]));
   NOR2_X1 i_142 (.A1(n_305), .A2(n_107), .ZN(n_103));
   OAI21_X1 i_143 (.A(n_320), .B1(b[60]), .B2(a[60]), .ZN(n_104));
   XNOR2_X1 i_144 (.A(n_110), .B(n_105), .ZN(sum[61]));
   OAI21_X1 i_145 (.A(n_320), .B1(n_315), .B2(n_107), .ZN(n_105));
   NOR2_X1 i_146 (.A1(n_306), .A2(n_317), .ZN(n_107));
   OAI22_X1 i_147 (.A1(b[61]), .A2(a[61]), .B1(n_321), .B2(n_323), .ZN(n_110));
   INV_X1 i_179 (.A(n_130), .ZN(n_125));
   NAND2_X1 i_183 (.A1(b[42]), .A2(a[42]), .ZN(n_129));
   INV_X1 i_197 (.A(n_235), .ZN(n_143));
   INV_X1 i_201 (.A(n_220), .ZN(n_147));
   INV_X1 i_221 (.A(n_180), .ZN(n_167));
   INV_X1 i_226 (.A(n_183), .ZN(n_172));
   AND2_X1 i_148 (.A1(b[39]), .A2(a[39]), .ZN(n_94));
   INV_X1 i_149 (.A(n_177), .ZN(n_95));
   NAND2_X1 i_150 (.A1(b[38]), .A2(a[38]), .ZN(n_177));
   INV_X1 i_235 (.A(n_174), .ZN(n_181));
   INV_X1 i_151 (.A(n_192), .ZN(n_188));
   INV_X1 i_152 (.A(n_196), .ZN(n_96));
   NOR2_X1 i_153 (.A1(b[28]), .A2(a[28]), .ZN(n_196));
   INV_X1 i_154 (.A(n_198), .ZN(n_97));
   NOR2_X1 i_155 (.A1(b[27]), .A2(a[27]), .ZN(n_198));
   NOR2_X1 i_156 (.A1(b[34]), .A2(a[34]), .ZN(n_98));
   INV_X1 i_157 (.A(n_207), .ZN(n_100));
   NOR2_X1 i_158 (.A1(b[36]), .A2(a[36]), .ZN(n_207));
   INV_X1 i_159 (.A(n_209), .ZN(n_101));
   NOR2_X1 i_160 (.A1(b[35]), .A2(a[35]), .ZN(n_209));
   NOR3_X1 i_161 (.A1(n_184), .A2(n_215), .A3(n_216), .ZN(n_102));
   NOR2_X1 i_162 (.A1(n_216), .A2(n_215), .ZN(n_214));
   NOR2_X1 i_163 (.A1(b[40]), .A2(a[40]), .ZN(n_215));
   NOR2_X1 i_164 (.A1(b[39]), .A2(a[39]), .ZN(n_216));
   INV_X1 i_166 (.A(n_221), .ZN(n_106));
   NOR2_X1 i_167 (.A1(b[32]), .A2(a[32]), .ZN(n_221));
   INV_X1 i_168 (.A(n_223), .ZN(n_108));
   NOR2_X1 i_169 (.A1(b[31]), .A2(a[31]), .ZN(n_223));
   INV_X1 i_170 (.A(n_164), .ZN(n_229));
   NOR2_X1 i_171 (.A1(b[24]), .A2(a[24]), .ZN(n_109));
   NOR2_X1 i_172 (.A1(b[23]), .A2(a[23]), .ZN(n_111));
   NOR2_X1 i_173 (.A1(n_254), .A2(n_244), .ZN(n_112));
   INV_X1 i_174 (.A(n_244), .ZN(n_243));
   NAND2_X1 i_175 (.A1(b[20]), .A2(a[20]), .ZN(n_244));
   AND2_X1 i_176 (.A1(b[21]), .A2(a[21]), .ZN(n_113));
   AOI21_X1 i_177 (.A(n_251), .B1(n_248), .B2(n_247), .ZN(n_114));
   NAND2_X1 i_178 (.A1(b[19]), .A2(a[19]), .ZN(n_247));
   NAND2_X1 i_180 (.A1(b[18]), .A2(a[18]), .ZN(n_248));
   NOR3_X1 i_181 (.A1(n_251), .A2(n_250), .A3(n_255), .ZN(n_115));
   NOR2_X1 i_182 (.A1(b[18]), .A2(a[18]), .ZN(n_250));
   OR3_X1 i_184 (.A1(n_254), .A2(n_252), .A3(n_253), .ZN(n_251));
   NOR2_X1 i_185 (.A1(b[20]), .A2(a[20]), .ZN(n_252));
   NOR2_X1 i_186 (.A1(b[19]), .A2(a[19]), .ZN(n_253));
   NOR2_X1 i_187 (.A1(b[21]), .A2(a[21]), .ZN(n_254));
   NOR4_X1 i_188 (.A1(n_259), .A2(n_256), .A3(n_260), .A4(n_263), .ZN(n_255));
   NOR2_X1 i_189 (.A1(n_268), .A2(n_258), .ZN(n_256));
   INV_X1 i_190 (.A(n_258), .ZN(n_257));
   NAND2_X1 i_191 (.A1(b[16]), .A2(a[16]), .ZN(n_258));
   AND2_X1 i_192 (.A1(b[17]), .A2(a[17]), .ZN(n_259));
   AOI21_X1 i_193 (.A(n_265), .B1(n_262), .B2(n_261), .ZN(n_260));
   NAND2_X1 i_194 (.A1(b[15]), .A2(a[15]), .ZN(n_261));
   NAND2_X1 i_195 (.A1(b[14]), .A2(a[14]), .ZN(n_262));
   NOR3_X1 i_196 (.A1(n_265), .A2(n_264), .A3(n_269), .ZN(n_263));
   NOR2_X1 i_198 (.A1(b[14]), .A2(a[14]), .ZN(n_264));
   OR3_X1 i_199 (.A1(n_268), .A2(n_266), .A3(n_267), .ZN(n_265));
   NOR2_X1 i_200 (.A1(b[16]), .A2(a[16]), .ZN(n_266));
   NOR2_X1 i_202 (.A1(b[15]), .A2(a[15]), .ZN(n_267));
   NOR2_X1 i_203 (.A1(b[17]), .A2(a[17]), .ZN(n_268));
   OAI22_X1 i_204 (.A1(b[13]), .A2(a[13]), .B1(n_277), .B2(n_270), .ZN(n_269));
   NAND2_X1 i_205 (.A1(n_276), .A2(n_271), .ZN(n_270));
   OAI21_X1 i_206 (.A(n_272), .B1(b[12]), .B2(a[12]), .ZN(n_271));
   AOI21_X1 i_207 (.A(n_275), .B1(n_274), .B2(n_273), .ZN(n_272));
   NAND2_X1 i_208 (.A1(b[11]), .A2(a[11]), .ZN(n_273));
   NAND2_X1 i_209 (.A1(b[10]), .A2(a[10]), .ZN(n_274));
   NOR2_X1 i_210 (.A1(b[11]), .A2(a[11]), .ZN(n_275));
   NAND2_X1 i_211 (.A1(b[12]), .A2(a[12]), .ZN(n_276));
   AND2_X1 i_212 (.A1(b[13]), .A2(a[13]), .ZN(n_277));
   NOR2_X1 i_336 (.A1(n_226), .A2(n_227), .ZN(n_282));
   INV_X1 i_165 (.A(n_238), .ZN(n_141));
   NOR2_X1 i_213 (.A1(a[47]), .A2(b[47]), .ZN(n_116));
   NOR2_X1 i_214 (.A1(a[48]), .A2(b[48]), .ZN(n_117));
   XOR2_X1 i_215 (.A(n_121), .B(n_118), .Z(sum[55]));
   NOR2_X1 i_216 (.A1(n_120), .A2(n_119), .ZN(n_118));
   AND2_X1 i_217 (.A1(b[55]), .A2(a[55]), .ZN(n_119));
   NOR2_X1 i_218 (.A1(b[55]), .A2(a[55]), .ZN(n_120));
   INV_X1 i_219 (.A(n_122), .ZN(n_121));
   OAI22_X1 i_220 (.A1(b[54]), .A2(a[54]), .B1(n_240), .B2(n_123), .ZN(n_122));
   OAI21_X1 i_222 (.A(n_210), .B1(n_205), .B2(n_124), .ZN(n_123));
   NOR2_X1 i_223 (.A1(n_127), .A2(n_126), .ZN(n_124));
   NOR2_X1 i_224 (.A1(n_144), .A2(n_132), .ZN(n_126));
   OAI222_X1 i_225 (.A1(n_133), .A2(n_128), .B1(n_142), .B2(n_130), .C1(n_249), 
      .C2(n_246), .ZN(n_127));
   AOI21_X1 i_227 (.A(n_131), .B1(b[42]), .B2(a[42]), .ZN(n_128));
   NAND2_X1 i_228 (.A1(b[44]), .A2(a[44]), .ZN(n_130));
   AND2_X1 i_229 (.A1(b[43]), .A2(a[43]), .ZN(n_131));
   OAI21_X1 i_230 (.A(n_134), .B1(b[42]), .B2(a[42]), .ZN(n_132));
   INV_X1 i_231 (.A(n_134), .ZN(n_133));
   NOR3_X1 i_232 (.A1(n_142), .A2(n_137), .A3(n_139), .ZN(n_134));
   NOR2_X1 i_233 (.A1(b[42]), .A2(a[42]), .ZN(n_135));
   INV_X1 i_234 (.A(n_137), .ZN(n_136));
   NOR2_X1 i_236 (.A1(b[43]), .A2(a[43]), .ZN(n_137));
   INV_X1 i_237 (.A(n_139), .ZN(n_138));
   NOR2_X1 i_238 (.A1(b[44]), .A2(a[44]), .ZN(n_139));
   INV_X1 i_239 (.A(n_142), .ZN(n_140));
   NOR2_X1 i_240 (.A1(b[45]), .A2(a[45]), .ZN(n_142));
   NOR3_X1 i_241 (.A1(n_151), .A2(n_146), .A3(n_145), .ZN(n_144));
   NOR3_X1 i_242 (.A1(n_168), .A2(n_152), .A3(n_155), .ZN(n_145));
   OAI221_X1 i_243 (.A(n_148), .B1(n_176), .B2(n_154), .C1(n_170), .C2(n_153), 
      .ZN(n_146));
   AOI21_X1 i_244 (.A(n_149), .B1(b[41]), .B2(a[41]), .ZN(n_148));
   OAI21_X1 i_245 (.A(n_150), .B1(n_184), .B2(n_183), .ZN(n_149));
   OAI21_X1 i_246 (.A(n_102), .B1(n_95), .B2(n_94), .ZN(n_150));
   NOR2_X1 i_247 (.A1(n_185), .A2(n_152), .ZN(n_151));
   OR2_X1 i_248 (.A1(n_200), .A2(n_153), .ZN(n_152));
   OR2_X1 i_249 (.A1(n_194), .A2(n_154), .ZN(n_153));
   OAI21_X1 i_250 (.A(n_102), .B1(b[38]), .B2(a[38]), .ZN(n_154));
   NOR4_X1 i_251 (.A1(n_166), .A2(n_156), .A3(n_157), .A4(n_158), .ZN(n_155));
   NOR2_X1 i_252 (.A1(n_165), .A2(n_164), .ZN(n_156));
   AOI21_X1 i_253 (.A(n_159), .B1(n_163), .B2(n_162), .ZN(n_157));
   NOR3_X1 i_254 (.A1(n_161), .A2(n_159), .A3(n_160), .ZN(n_158));
   OR3_X1 i_255 (.A1(n_109), .A2(n_165), .A3(n_111), .ZN(n_159));
   NOR4_X1 i_256 (.A1(n_113), .A2(n_112), .A3(n_114), .A4(n_115), .ZN(n_160));
   NOR2_X1 i_257 (.A1(b[22]), .A2(a[22]), .ZN(n_161));
   NAND2_X1 i_258 (.A1(b[23]), .A2(a[23]), .ZN(n_162));
   NAND2_X1 i_259 (.A1(b[22]), .A2(a[22]), .ZN(n_163));
   NAND2_X1 i_260 (.A1(b[24]), .A2(a[24]), .ZN(n_164));
   NOR2_X1 i_261 (.A1(b[25]), .A2(a[25]), .ZN(n_165));
   AND2_X1 i_262 (.A1(b[25]), .A2(a[25]), .ZN(n_166));
   OR2_X1 i_263 (.A1(n_187), .A2(n_169), .ZN(n_168));
   NOR2_X1 i_264 (.A1(b[26]), .A2(a[26]), .ZN(n_169));
   AOI221_X1 i_265 (.A(n_171), .B1(n_202), .B2(n_173), .C1(b[33]), .C2(a[33]), 
      .ZN(n_170));
   AOI21_X1 i_266 (.A(n_201), .B1(n_175), .B2(n_174), .ZN(n_171));
   AND2_X1 i_267 (.A1(b[32]), .A2(a[32]), .ZN(n_173));
   NAND2_X1 i_268 (.A1(b[31]), .A2(a[31]), .ZN(n_174));
   NAND2_X1 i_269 (.A1(b[30]), .A2(a[30]), .ZN(n_175));
   AOI221_X1 i_270 (.A(n_178), .B1(b[37]), .B2(a[37]), .C1(n_197), .C2(n_179), 
      .ZN(n_176));
   AOI21_X1 i_271 (.A(n_195), .B1(n_182), .B2(n_180), .ZN(n_178));
   AND2_X1 i_272 (.A1(b[36]), .A2(a[36]), .ZN(n_179));
   NAND2_X1 i_273 (.A1(b[35]), .A2(a[35]), .ZN(n_180));
   NAND2_X1 i_274 (.A1(b[34]), .A2(a[34]), .ZN(n_182));
   NAND2_X1 i_275 (.A1(b[40]), .A2(a[40]), .ZN(n_183));
   NOR2_X1 i_276 (.A1(b[41]), .A2(a[41]), .ZN(n_184));
   AOI221_X1 i_277 (.A(n_186), .B1(n_190), .B2(n_189), .C1(b[29]), .C2(a[29]), 
      .ZN(n_185));
   AOI21_X1 i_278 (.A(n_187), .B1(n_193), .B2(n_192), .ZN(n_186));
   NAND3_X1 i_279 (.A1(n_96), .A2(n_190), .A3(n_97), .ZN(n_187));
   AND2_X1 i_280 (.A1(b[28]), .A2(a[28]), .ZN(n_189));
   INV_X1 i_281 (.A(n_191), .ZN(n_190));
   NOR2_X1 i_282 (.A1(b[29]), .A2(a[29]), .ZN(n_191));
   NAND2_X1 i_283 (.A1(b[27]), .A2(a[27]), .ZN(n_192));
   NAND2_X1 i_284 (.A1(b[26]), .A2(a[26]), .ZN(n_193));
   OR2_X1 i_285 (.A1(n_98), .A2(n_195), .ZN(n_194));
   NAND3_X1 i_286 (.A1(n_100), .A2(n_197), .A3(n_101), .ZN(n_195));
   INV_X1 i_287 (.A(n_199), .ZN(n_197));
   NOR2_X1 i_288 (.A1(b[37]), .A2(a[37]), .ZN(n_199));
   OR2_X1 i_289 (.A1(n_204), .A2(n_201), .ZN(n_200));
   NAND3_X1 i_290 (.A1(n_106), .A2(n_202), .A3(n_108), .ZN(n_201));
   INV_X1 i_291 (.A(n_203), .ZN(n_202));
   NOR2_X1 i_292 (.A1(b[33]), .A2(a[33]), .ZN(n_203));
   NOR2_X1 i_293 (.A1(b[30]), .A2(a[30]), .ZN(n_204));
   OR2_X1 i_294 (.A1(n_218), .A2(n_206), .ZN(n_205));
   OAI21_X1 i_295 (.A(n_233), .B1(b[46]), .B2(a[46]), .ZN(n_206));
   NOR2_X1 i_296 (.A1(b[46]), .A2(a[46]), .ZN(n_208));
   INV_X1 i_297 (.A(n_211), .ZN(n_210));
   OAI211_X1 i_298 (.A(n_212), .B(n_213), .C1(n_230), .C2(n_218), .ZN(n_211));
   OAI21_X1 i_299 (.A(n_219), .B1(n_224), .B2(n_222), .ZN(n_212));
   AOI21_X1 i_300 (.A(n_217), .B1(b[53]), .B2(a[53]), .ZN(n_213));
   NOR2_X1 i_301 (.A1(n_228), .A2(n_220), .ZN(n_217));
   OAI21_X1 i_302 (.A(n_219), .B1(b[50]), .B2(a[50]), .ZN(n_218));
   NOR3_X1 i_303 (.A1(n_228), .A2(n_226), .A3(n_227), .ZN(n_219));
   NAND2_X1 i_304 (.A1(b[52]), .A2(a[52]), .ZN(n_220));
   AND2_X1 i_305 (.A1(b[51]), .A2(a[51]), .ZN(n_222));
   INV_X1 i_306 (.A(n_225), .ZN(n_224));
   NAND2_X1 i_307 (.A1(b[50]), .A2(a[50]), .ZN(n_225));
   NOR2_X1 i_308 (.A1(b[51]), .A2(a[51]), .ZN(n_226));
   NOR2_X1 i_309 (.A1(b[52]), .A2(a[52]), .ZN(n_227));
   NOR2_X1 i_310 (.A1(b[53]), .A2(a[53]), .ZN(n_228));
   AOI21_X1 i_311 (.A(n_231), .B1(b[49]), .B2(a[49]), .ZN(n_230));
   OAI21_X1 i_312 (.A(n_232), .B1(n_239), .B2(n_238), .ZN(n_231));
   OAI21_X1 i_313 (.A(n_233), .B1(n_236), .B2(n_234), .ZN(n_232));
   NOR3_X1 i_314 (.A1(n_116), .A2(n_239), .A3(n_117), .ZN(n_233));
   INV_X1 i_315 (.A(n_235), .ZN(n_234));
   NAND2_X1 i_316 (.A1(b[47]), .A2(a[47]), .ZN(n_235));
   INV_X1 i_317 (.A(n_237), .ZN(n_236));
   NAND2_X1 i_318 (.A1(b[46]), .A2(a[46]), .ZN(n_237));
   NAND2_X1 i_319 (.A1(b[48]), .A2(a[48]), .ZN(n_238));
   NOR2_X1 i_320 (.A1(b[49]), .A2(a[49]), .ZN(n_239));
   INV_X1 i_321 (.A(n_241), .ZN(n_240));
   NAND2_X1 i_322 (.A1(b[54]), .A2(a[54]), .ZN(n_241));
   INV_X1 i_323 (.A(n_116), .ZN(n_242));
   INV_X1 i_324 (.A(n_117), .ZN(n_245));
   INV_X1 i_325 (.A(a[45]), .ZN(n_246));
   INV_X1 i_326 (.A(b[45]), .ZN(n_249));
   NOR2_X1 i_327 (.A1(a[57]), .A2(b[57]), .ZN(n_278));
   NAND2_X1 i_328 (.A1(a[56]), .A2(b[56]), .ZN(n_279));
   NOR2_X1 i_329 (.A1(a[56]), .A2(b[56]), .ZN(n_280));
   INV_X1 i_330 (.A(n_279), .ZN(n_281));
   NOR2_X1 i_331 (.A1(n_280), .A2(n_120), .ZN(n_283));
   NAND2_X1 i_332 (.A1(n_118), .A2(n_122), .ZN(n_284));
   AOI21_X1 i_333 (.A(n_281), .B1(n_283), .B2(n_284), .ZN(n_285));
   AOI21_X1 i_334 (.A(n_278), .B1(a[57]), .B2(b[57]), .ZN(n_286));
   XNOR2_X1 i_335 (.A(n_285), .B(n_286), .ZN(sum[57]));
   INV_X1 i_337 (.A(n_278), .ZN(n_287));
   XOR2_X1 i_338 (.A(n_290), .B(n_288), .Z(sum[58]));
   OAI21_X1 i_339 (.A(n_289), .B1(b[58]), .B2(a[58]), .ZN(n_288));
   NAND2_X1 i_340 (.A1(b[58]), .A2(a[58]), .ZN(n_289));
   AOI21_X1 i_341 (.A(n_293), .B1(n_292), .B2(n_291), .ZN(n_290));
   NOR2_X1 i_342 (.A1(n_205), .A2(n_297), .ZN(n_291));
   OAI21_X1 i_343 (.A(n_299), .B1(n_144), .B2(n_132), .ZN(n_292));
   OAI211_X1 i_344 (.A(n_294), .B(n_295), .C1(n_300), .C2(n_297), .ZN(n_293));
   OAI21_X1 i_345 (.A(n_298), .B1(n_240), .B2(n_119), .ZN(n_294));
   AOI21_X1 i_346 (.A(n_296), .B1(b[57]), .B2(a[57]), .ZN(n_295));
   NOR2_X1 i_347 (.A1(n_278), .A2(n_279), .ZN(n_296));
   OAI21_X1 i_348 (.A(n_298), .B1(b[54]), .B2(a[54]), .ZN(n_297));
   NOR3_X1 i_349 (.A1(n_120), .A2(n_301), .A3(n_280), .ZN(n_298));
   INV_X1 i_350 (.A(n_127), .ZN(n_299));
   INV_X1 i_351 (.A(n_211), .ZN(n_300));
   INV_X1 i_352 (.A(n_287), .ZN(n_301));
   XNOR2_X1 i_353 (.A(n_303), .B(n_302), .ZN(sum[59]));
   AOI21_X1 i_354 (.A(n_305), .B1(a[59]), .B2(b[59]), .ZN(n_302));
   AOI21_X1 i_355 (.A(n_306), .B1(a[58]), .B2(b[58]), .ZN(n_303));
   INV_X1 i_356 (.A(n_305), .ZN(n_304));
   NOR2_X1 i_357 (.A1(a[59]), .A2(b[59]), .ZN(n_305));
   NOR2_X1 i_358 (.A1(n_308), .A2(n_307), .ZN(n_306));
   AOI21_X1 i_359 (.A(n_293), .B1(n_292), .B2(n_291), .ZN(n_307));
   NOR2_X1 i_360 (.A1(a[58]), .A2(b[58]), .ZN(n_308));
   INV_X1 i_361 (.A(b[59]), .ZN(n_309));
   INV_X1 i_362 (.A(a[59]), .ZN(n_310));
   XNOR2_X1 i_363 (.A(n_312), .B(n_311), .ZN(sum[62]));
   OAI22_X1 i_364 (.A1(n_324), .A2(b[62]), .B1(a[62]), .B2(n_322), .ZN(n_311));
   AOI21_X1 i_365 (.A(n_318), .B1(n_314), .B2(n_313), .ZN(n_312));
   OAI21_X1 i_366 (.A(n_316), .B1(n_290), .B2(n_308), .ZN(n_313));
   NOR2_X1 i_367 (.A1(n_319), .A2(n_315), .ZN(n_314));
   OAI21_X1 i_368 (.A(n_304), .B1(a[60]), .B2(b[60]), .ZN(n_315));
   INV_X1 i_369 (.A(n_317), .ZN(n_316));
   OAI21_X1 i_370 (.A(n_289), .B1(n_310), .B2(n_309), .ZN(n_317));
   OAI22_X1 i_371 (.A1(n_323), .A2(n_321), .B1(n_320), .B2(n_319), .ZN(n_318));
   NOR2_X1 i_372 (.A1(a[61]), .A2(b[61]), .ZN(n_319));
   NAND2_X1 i_373 (.A1(a[60]), .A2(b[60]), .ZN(n_320));
   INV_X1 i_374 (.A(b[61]), .ZN(n_321));
   INV_X1 i_375 (.A(b[62]), .ZN(n_322));
   INV_X1 i_376 (.A(a[61]), .ZN(n_323));
   INV_X1 i_377 (.A(a[62]), .ZN(n_324));
   NAND2_X1 i_378 (.A1(n_328), .A2(n_325), .ZN(sum[63]));
   OR3_X1 i_379 (.A1(n_331), .A2(n_330), .A3(n_326), .ZN(n_325));
   AOI22_X1 i_380 (.A1(n_324), .A2(n_322), .B1(n_332), .B2(n_327), .ZN(n_326));
   OAI21_X1 i_381 (.A(n_314), .B1(n_306), .B2(n_317), .ZN(n_327));
   OAI21_X1 i_382 (.A(n_331), .B1(n_330), .B2(n_329), .ZN(n_328));
   AOI21_X1 i_383 (.A(n_312), .B1(n_324), .B2(n_322), .ZN(n_329));
   AND2_X1 i_384 (.A1(a[62]), .A2(b[62]), .ZN(n_330));
   XNOR2_X1 i_385 (.A(a[63]), .B(b[63]), .ZN(n_331));
   INV_X1 i_386 (.A(n_318), .ZN(n_332));
endmodule

module simple_Adder(a, b, cin, S);
   input [63:0]a;
   input [63:0]b;
   input cin;
   output [63:0]S;

   datapath i_0 (.b({b[63], b[62], b[61], b[60], b[59], b[58], b[57], b[56], 
      b[55], b[54], b[53], b[52], b[51], b[50], b[49], b[48], b[47], b[46], 
      b[45], b[44], b[43], b[42], b[41], b[40], b[39], b[38], b[37], b[36], 
      b[35], b[34], b[33], b[32], b[31], b[30], b[29], b[28], b[27], b[26], 
      b[25], b[24], b[23], b[22], b[21], b[20], b[19], b[18], b[17], b[16], 
      b[15], b[14], b[13], b[12], b[11], b[10], uc_0, uc_1, uc_2, uc_3, uc_4, 
      uc_5, uc_6, uc_7, uc_8, uc_9}), .cin(), .a({a[63], a[62], a[61], a[60], 
      a[59], a[58], a[57], a[56], a[55], a[54], a[53], a[52], a[51], a[50], 
      a[49], a[48], a[47], a[46], a[45], a[44], a[43], a[42], a[41], a[40], 
      a[39], a[38], a[37], a[36], a[35], a[34], a[33], a[32], a[31], a[30], 
      a[29], a[28], a[27], a[26], a[25], a[24], a[23], a[22], a[21], a[20], 
      a[19], a[18], a[17], a[16], a[15], a[14], a[13], a[12], a[11], a[10], 
      uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19}), 
      .sum({S[63], S[62], S[61], S[60], S[59], S[58], S[57], S[56], S[55], S[54], 
      S[53], S[52], S[51], S[50], S[49], S[48], S[47], S[46], S[45], S[44], 
      S[43], S[42], S[41], S[40], S[39], S[38], S[37], S[36], S[35], S[34], 
      S[33], S[32], S[31], S[30], S[29], S[28], S[27], S[26], S[25], S[24], 
      S[23], S[22], S[21], S[20], S[19], S[18], S[17], S[16], S[15], S[14], 
      S[13], S[12], S[11], S[10], uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, 
      uc_26, uc_27, uc_28, uc_29}));
endmodule

module CSA(in1, in2, in3, sum, c);
   input [63:0]in1;
   input [63:0]in2;
   input [63:0]in3;
   output [63:0]sum;
   output [63:0]c;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;

   AND2_X1 i_0_0 (.A1(in2[28]), .A2(in1[28]), .ZN(c[29]));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(c[30]));
   OAI21_X1 i_0_2 (.A(in2[29]), .B1(in3[29]), .B2(in1[29]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in3[29]), .A2(in1[29]), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_2), .ZN(c[31]));
   OAI21_X1 i_0_5 (.A(in2[30]), .B1(in3[30]), .B2(in1[30]), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(in3[30]), .A2(in1[30]), .ZN(n_0_3));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4), .ZN(c[32]));
   OAI21_X1 i_0_8 (.A(in2[31]), .B1(in3[31]), .B2(in1[31]), .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(in3[31]), .A2(in1[31]), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_7), .A2(n_0_6), .ZN(c[33]));
   OAI21_X1 i_0_11 (.A(in2[32]), .B1(in3[32]), .B2(in1[32]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in3[32]), .A2(in1[32]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_9), .A2(n_0_8), .ZN(c[34]));
   OAI21_X1 i_0_14 (.A(in2[33]), .B1(in3[33]), .B2(in1[33]), .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(in3[33]), .A2(in1[33]), .ZN(n_0_9));
   NAND2_X1 i_0_16 (.A1(n_0_11), .A2(n_0_10), .ZN(c[35]));
   OAI21_X1 i_0_17 (.A(in2[34]), .B1(in3[34]), .B2(in1[34]), .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(in3[34]), .A2(in1[34]), .ZN(n_0_11));
   NAND2_X1 i_0_19 (.A1(n_0_13), .A2(n_0_12), .ZN(c[36]));
   OAI21_X1 i_0_20 (.A(in2[35]), .B1(in3[35]), .B2(in1[35]), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(in3[35]), .A2(in1[35]), .ZN(n_0_13));
   NAND2_X1 i_0_22 (.A1(n_0_15), .A2(n_0_14), .ZN(c[37]));
   OAI21_X1 i_0_23 (.A(in2[36]), .B1(in3[36]), .B2(in1[36]), .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(in3[36]), .A2(in1[36]), .ZN(n_0_15));
   NAND2_X1 i_0_25 (.A1(n_0_17), .A2(n_0_16), .ZN(c[38]));
   OAI21_X1 i_0_26 (.A(in2[37]), .B1(in3[37]), .B2(in1[37]), .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(in3[37]), .A2(in1[37]), .ZN(n_0_17));
   NAND2_X1 i_0_28 (.A1(n_0_19), .A2(n_0_18), .ZN(c[39]));
   OAI21_X1 i_0_29 (.A(in2[38]), .B1(in3[38]), .B2(in1[38]), .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(in3[38]), .A2(in1[38]), .ZN(n_0_19));
   NAND2_X1 i_0_31 (.A1(n_0_21), .A2(n_0_20), .ZN(c[40]));
   OAI21_X1 i_0_32 (.A(in2[39]), .B1(in3[39]), .B2(in1[39]), .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(in3[39]), .A2(in1[39]), .ZN(n_0_21));
   NAND2_X1 i_0_34 (.A1(n_0_23), .A2(n_0_22), .ZN(c[41]));
   OAI21_X1 i_0_35 (.A(in2[40]), .B1(in3[40]), .B2(in1[40]), .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(in3[40]), .A2(in1[40]), .ZN(n_0_23));
   NAND2_X1 i_0_37 (.A1(n_0_25), .A2(n_0_24), .ZN(c[42]));
   OAI21_X1 i_0_38 (.A(in2[41]), .B1(in3[41]), .B2(in1[41]), .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(in3[41]), .A2(in1[41]), .ZN(n_0_25));
   NAND2_X1 i_0_40 (.A1(n_0_27), .A2(n_0_26), .ZN(c[43]));
   OAI21_X1 i_0_41 (.A(in2[42]), .B1(in3[42]), .B2(in1[42]), .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(in3[42]), .A2(in1[42]), .ZN(n_0_27));
   NAND2_X1 i_0_43 (.A1(n_0_29), .A2(n_0_28), .ZN(c[44]));
   OAI21_X1 i_0_44 (.A(in2[43]), .B1(in3[43]), .B2(in1[43]), .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(in3[43]), .A2(in1[43]), .ZN(n_0_29));
   NAND2_X1 i_0_46 (.A1(n_0_31), .A2(n_0_30), .ZN(c[45]));
   OAI21_X1 i_0_47 (.A(in2[44]), .B1(in3[44]), .B2(in1[44]), .ZN(n_0_30));
   NAND2_X1 i_0_48 (.A1(in3[44]), .A2(in1[44]), .ZN(n_0_31));
   NAND2_X1 i_0_49 (.A1(n_0_33), .A2(n_0_32), .ZN(c[46]));
   OAI21_X1 i_0_50 (.A(in2[45]), .B1(in3[45]), .B2(in1[45]), .ZN(n_0_32));
   NAND2_X1 i_0_51 (.A1(in3[45]), .A2(in1[45]), .ZN(n_0_33));
   NAND2_X1 i_0_52 (.A1(n_0_35), .A2(n_0_34), .ZN(c[47]));
   OAI21_X1 i_0_53 (.A(in2[46]), .B1(in3[46]), .B2(in1[46]), .ZN(n_0_34));
   NAND2_X1 i_0_54 (.A1(in3[46]), .A2(in1[46]), .ZN(n_0_35));
   NAND2_X1 i_0_55 (.A1(n_0_37), .A2(n_0_36), .ZN(c[48]));
   OAI21_X1 i_0_56 (.A(in2[47]), .B1(in3[47]), .B2(in1[47]), .ZN(n_0_36));
   NAND2_X1 i_0_57 (.A1(in3[47]), .A2(in1[47]), .ZN(n_0_37));
   NAND2_X1 i_0_58 (.A1(n_0_39), .A2(n_0_38), .ZN(c[49]));
   OAI21_X1 i_0_59 (.A(in2[48]), .B1(in3[48]), .B2(in1[48]), .ZN(n_0_38));
   NAND2_X1 i_0_60 (.A1(in3[48]), .A2(in1[48]), .ZN(n_0_39));
   NAND2_X1 i_0_61 (.A1(n_0_41), .A2(n_0_40), .ZN(c[50]));
   OAI21_X1 i_0_62 (.A(in2[49]), .B1(in3[49]), .B2(in1[49]), .ZN(n_0_40));
   NAND2_X1 i_0_63 (.A1(in3[49]), .A2(in1[49]), .ZN(n_0_41));
   NAND2_X1 i_0_64 (.A1(n_0_43), .A2(n_0_42), .ZN(c[51]));
   OAI21_X1 i_0_65 (.A(in2[50]), .B1(in3[50]), .B2(in1[50]), .ZN(n_0_42));
   NAND2_X1 i_0_66 (.A1(in3[50]), .A2(in1[50]), .ZN(n_0_43));
   NAND2_X1 i_0_67 (.A1(n_0_45), .A2(n_0_44), .ZN(c[52]));
   OAI21_X1 i_0_68 (.A(in2[51]), .B1(in3[51]), .B2(in1[51]), .ZN(n_0_44));
   NAND2_X1 i_0_69 (.A1(in3[51]), .A2(in1[51]), .ZN(n_0_45));
   NAND2_X1 i_0_70 (.A1(n_0_47), .A2(n_0_46), .ZN(c[53]));
   OAI21_X1 i_0_71 (.A(in2[52]), .B1(in3[52]), .B2(in1[52]), .ZN(n_0_46));
   NAND2_X1 i_0_72 (.A1(in3[52]), .A2(in1[52]), .ZN(n_0_47));
   NAND2_X1 i_0_73 (.A1(n_0_49), .A2(n_0_48), .ZN(c[54]));
   OAI21_X1 i_0_74 (.A(in2[53]), .B1(in3[53]), .B2(in1[53]), .ZN(n_0_48));
   NAND2_X1 i_0_75 (.A1(in3[53]), .A2(in1[53]), .ZN(n_0_49));
   NAND2_X1 i_0_76 (.A1(n_0_51), .A2(n_0_50), .ZN(c[55]));
   OAI21_X1 i_0_77 (.A(in2[54]), .B1(in3[54]), .B2(in1[54]), .ZN(n_0_50));
   NAND2_X1 i_0_78 (.A1(in3[54]), .A2(in1[54]), .ZN(n_0_51));
   NAND2_X1 i_0_79 (.A1(n_0_53), .A2(n_0_52), .ZN(c[56]));
   OAI21_X1 i_0_80 (.A(in2[55]), .B1(in3[55]), .B2(in1[55]), .ZN(n_0_52));
   NAND2_X1 i_0_81 (.A1(in3[55]), .A2(in1[55]), .ZN(n_0_53));
   NAND2_X1 i_0_82 (.A1(n_0_55), .A2(n_0_54), .ZN(c[57]));
   OAI21_X1 i_0_83 (.A(in2[56]), .B1(in3[56]), .B2(in1[56]), .ZN(n_0_54));
   NAND2_X1 i_0_84 (.A1(in3[56]), .A2(in1[56]), .ZN(n_0_55));
   NAND2_X1 i_0_85 (.A1(n_0_57), .A2(n_0_56), .ZN(c[58]));
   OAI21_X1 i_0_86 (.A(in2[57]), .B1(in3[57]), .B2(in1[57]), .ZN(n_0_56));
   NAND2_X1 i_0_87 (.A1(in3[57]), .A2(in1[57]), .ZN(n_0_57));
   NAND2_X1 i_0_88 (.A1(n_0_59), .A2(n_0_58), .ZN(c[59]));
   OAI21_X1 i_0_89 (.A(in2[58]), .B1(in3[58]), .B2(in1[63]), .ZN(n_0_58));
   NAND2_X1 i_0_90 (.A1(in3[58]), .A2(in1[63]), .ZN(n_0_59));
   NAND2_X1 i_0_91 (.A1(n_0_62), .A2(n_0_60), .ZN(c[60]));
   OAI21_X1 i_0_92 (.A(in3[59]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_60));
   NAND2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(c[63]));
   OAI21_X1 i_0_94 (.A(in3[63]), .B1(in1[63]), .B2(in2[63]), .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(in2[63]), .A2(in1[63]), .ZN(n_0_62));
   XOR2_X1 i_0_96 (.A(in2[28]), .B(in1[28]), .Z(sum[28]));
   XNOR2_X1 i_0_97 (.A(in2[29]), .B(n_0_63), .ZN(sum[29]));
   XNOR2_X1 i_0_98 (.A(in3[29]), .B(in1[29]), .ZN(n_0_63));
   XNOR2_X1 i_0_99 (.A(in2[30]), .B(n_0_64), .ZN(sum[30]));
   XNOR2_X1 i_0_100 (.A(in3[30]), .B(in1[30]), .ZN(n_0_64));
   XNOR2_X1 i_0_101 (.A(in2[31]), .B(n_0_65), .ZN(sum[31]));
   XNOR2_X1 i_0_102 (.A(in3[31]), .B(in1[31]), .ZN(n_0_65));
   XNOR2_X1 i_0_103 (.A(in2[32]), .B(n_0_66), .ZN(sum[32]));
   XNOR2_X1 i_0_104 (.A(in3[32]), .B(in1[32]), .ZN(n_0_66));
   XNOR2_X1 i_0_105 (.A(in2[33]), .B(n_0_67), .ZN(sum[33]));
   XNOR2_X1 i_0_106 (.A(in3[33]), .B(in1[33]), .ZN(n_0_67));
   XNOR2_X1 i_0_107 (.A(in2[34]), .B(n_0_68), .ZN(sum[34]));
   XNOR2_X1 i_0_108 (.A(in3[34]), .B(in1[34]), .ZN(n_0_68));
   XNOR2_X1 i_0_109 (.A(in2[35]), .B(n_0_69), .ZN(sum[35]));
   XNOR2_X1 i_0_110 (.A(in3[35]), .B(in1[35]), .ZN(n_0_69));
   XNOR2_X1 i_0_111 (.A(in2[36]), .B(n_0_70), .ZN(sum[36]));
   XNOR2_X1 i_0_112 (.A(in3[36]), .B(in1[36]), .ZN(n_0_70));
   XNOR2_X1 i_0_113 (.A(in2[37]), .B(n_0_71), .ZN(sum[37]));
   XNOR2_X1 i_0_114 (.A(in3[37]), .B(in1[37]), .ZN(n_0_71));
   XNOR2_X1 i_0_115 (.A(in2[38]), .B(n_0_72), .ZN(sum[38]));
   XNOR2_X1 i_0_116 (.A(in3[38]), .B(in1[38]), .ZN(n_0_72));
   XNOR2_X1 i_0_117 (.A(in2[39]), .B(n_0_73), .ZN(sum[39]));
   XNOR2_X1 i_0_118 (.A(in3[39]), .B(in1[39]), .ZN(n_0_73));
   XNOR2_X1 i_0_119 (.A(in2[40]), .B(n_0_74), .ZN(sum[40]));
   XNOR2_X1 i_0_120 (.A(in3[40]), .B(in1[40]), .ZN(n_0_74));
   XNOR2_X1 i_0_121 (.A(in2[41]), .B(n_0_75), .ZN(sum[41]));
   XNOR2_X1 i_0_122 (.A(in3[41]), .B(in1[41]), .ZN(n_0_75));
   XNOR2_X1 i_0_123 (.A(in2[42]), .B(n_0_76), .ZN(sum[42]));
   XNOR2_X1 i_0_124 (.A(in3[42]), .B(in1[42]), .ZN(n_0_76));
   XNOR2_X1 i_0_125 (.A(in2[43]), .B(n_0_77), .ZN(sum[43]));
   XNOR2_X1 i_0_126 (.A(in3[43]), .B(in1[43]), .ZN(n_0_77));
   XNOR2_X1 i_0_127 (.A(in2[44]), .B(n_0_78), .ZN(sum[44]));
   XNOR2_X1 i_0_128 (.A(in3[44]), .B(in1[44]), .ZN(n_0_78));
   XNOR2_X1 i_0_129 (.A(in2[45]), .B(n_0_79), .ZN(sum[45]));
   XNOR2_X1 i_0_130 (.A(in3[45]), .B(in1[45]), .ZN(n_0_79));
   XNOR2_X1 i_0_131 (.A(in2[46]), .B(n_0_80), .ZN(sum[46]));
   XNOR2_X1 i_0_132 (.A(in3[46]), .B(in1[46]), .ZN(n_0_80));
   XNOR2_X1 i_0_133 (.A(in2[47]), .B(n_0_81), .ZN(sum[47]));
   XNOR2_X1 i_0_134 (.A(in3[47]), .B(in1[47]), .ZN(n_0_81));
   XNOR2_X1 i_0_135 (.A(in2[48]), .B(n_0_82), .ZN(sum[48]));
   XNOR2_X1 i_0_136 (.A(in3[48]), .B(in1[48]), .ZN(n_0_82));
   XNOR2_X1 i_0_137 (.A(in2[49]), .B(n_0_83), .ZN(sum[49]));
   XNOR2_X1 i_0_138 (.A(in3[49]), .B(in1[49]), .ZN(n_0_83));
   XNOR2_X1 i_0_139 (.A(in2[50]), .B(n_0_84), .ZN(sum[50]));
   XNOR2_X1 i_0_140 (.A(in3[50]), .B(in1[50]), .ZN(n_0_84));
   XNOR2_X1 i_0_141 (.A(in2[51]), .B(n_0_85), .ZN(sum[51]));
   XNOR2_X1 i_0_142 (.A(in3[51]), .B(in1[51]), .ZN(n_0_85));
   XNOR2_X1 i_0_143 (.A(in2[52]), .B(n_0_86), .ZN(sum[52]));
   XNOR2_X1 i_0_144 (.A(in3[52]), .B(in1[52]), .ZN(n_0_86));
   XNOR2_X1 i_0_145 (.A(in2[53]), .B(n_0_87), .ZN(sum[53]));
   XNOR2_X1 i_0_146 (.A(in3[53]), .B(in1[53]), .ZN(n_0_87));
   XNOR2_X1 i_0_147 (.A(in2[54]), .B(n_0_88), .ZN(sum[54]));
   XNOR2_X1 i_0_148 (.A(in3[54]), .B(in1[54]), .ZN(n_0_88));
   XNOR2_X1 i_0_149 (.A(in2[55]), .B(n_0_89), .ZN(sum[55]));
   XNOR2_X1 i_0_150 (.A(in3[55]), .B(in1[55]), .ZN(n_0_89));
   XNOR2_X1 i_0_151 (.A(in2[56]), .B(n_0_90), .ZN(sum[56]));
   XNOR2_X1 i_0_152 (.A(in3[56]), .B(in1[56]), .ZN(n_0_90));
   XNOR2_X1 i_0_153 (.A(in2[57]), .B(n_0_91), .ZN(sum[57]));
   XNOR2_X1 i_0_154 (.A(in3[57]), .B(in1[57]), .ZN(n_0_91));
   XNOR2_X1 i_0_155 (.A(in2[58]), .B(n_0_92), .ZN(sum[58]));
   XNOR2_X1 i_0_156 (.A(in3[58]), .B(in1[63]), .ZN(n_0_92));
   XOR2_X1 i_0_157 (.A(in3[59]), .B(n_0_93), .Z(sum[59]));
   XOR2_X1 i_0_158 (.A(in3[63]), .B(n_0_93), .Z(sum[63]));
   XOR2_X1 i_0_159 (.A(in2[63]), .B(in1[63]), .Z(n_0_93));
endmodule

module wallace(a, b, c);
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   wire [63:0]\c1[0] ;
   wire [63:0]\s1[0] ;
   wire [63:0]\c1[1] ;
   wire [63:0]\s1[1] ;
   wire [63:0]\c2[0] ;
   wire [63:0]\s2[0] ;
   wire [63:0]\c1[2] ;
   wire [63:0]\s1[2] ;
   wire [63:0]\c2[1] ;
   wire [63:0]\s2[1] ;
   wire [63:0]\c3[0] ;
   wire [63:0]\s3[0] ;
   wire [63:0]\c1[3] ;
   wire [63:0]\s1[3] ;
   wire [63:0]\c1[8] ;
   wire [63:0]\s1[8] ;
   wire [63:0]\c2[2] ;
   wire [63:0]\s2[2] ;
   wire [63:0]\c3[1] ;
   wire [63:0]\s3[1] ;
   wire [63:0]\c4[0] ;
   wire [63:0]\s4[0] ;
   wire [63:0]\c2[5] ;
   wire [63:0]\s2[5] ;
   wire [63:0]\c3[3] ;
   wire [63:0]\s3[3] ;
   wire [63:0]\c1[7] ;
   wire [63:0]\s1[7] ;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0;
   wire n_0_0_3;
   wire n_0_1;
   wire n_0_0_4;
   wire n_0_2;
   wire n_0_0_5;
   wire n_0_3;
   wire n_0_0_6;
   wire n_0_4;
   wire n_0_0_7;
   wire n_0_5;
   wire n_0_0_8;
   wire n_0_6;
   wire n_0_0_9;
   wire n_0_7;
   wire n_0_0_10;
   wire n_0_8;
   wire n_0_0_11;
   wire n_0_9;
   wire n_0_0_12;
   wire n_0_10;
   wire n_0_0_13;
   wire n_0_11;
   wire n_0_0_14;
   wire n_0_12;
   wire n_0_0_15;
   wire n_0_13;
   wire n_0_0_16;
   wire n_0_14;
   wire n_0_0_17;
   wire n_0_15;
   wire n_0_0_18;
   wire n_0_16;
   wire n_0_0_19;
   wire n_0_17;
   wire n_0_0_20;
   wire n_0_18;
   wire n_0_0_21;
   wire n_0_19;
   wire n_0_0_22;
   wire n_0_20;
   wire n_0_0_23;
   wire n_0_21;
   wire n_0_0_24;
   wire n_0_22;
   wire n_0_0_25;
   wire n_0_23;
   wire n_0_0_26;
   wire n_0_24;
   wire n_0_0_27;
   wire n_0_25;
   wire n_0_0_28;
   wire n_0_26;
   wire n_0_0_29;
   wire n_0_27;
   wire n_0_0_30;
   wire n_0_28;
   wire n_0_0_31;
   wire n_0_29;
   wire n_0_544;
   wire n_0_545;
   wire n_0_546;
   wire n_0_547;
   wire n_0_548;
   wire n_0_549;
   wire n_0_550;
   wire n_0_551;
   wire n_0_552;
   wire n_0_553;
   wire n_0_554;
   wire n_0_555;
   wire n_0_556;
   wire n_0_557;
   wire n_0_558;
   wire n_0_559;
   wire n_0_560;
   wire n_0_561;
   wire n_0_562;
   wire n_0_563;
   wire n_0_564;
   wire n_0_565;
   wire n_0_566;
   wire n_0_567;
   wire n_0_568;
   wire n_0_569;
   wire n_0_570;
   wire n_0_571;
   wire n_0_572;
   wire n_0_573;
   wire n_0_31;
   wire n_0_0_34;
   wire n_0_512;
   wire n_0_513;
   wire n_0_514;
   wire n_0_515;
   wire n_0_516;
   wire n_0_517;
   wire n_0_518;
   wire n_0_519;
   wire n_0_520;
   wire n_0_521;
   wire n_0_522;
   wire n_0_523;
   wire n_0_524;
   wire n_0_525;
   wire n_0_526;
   wire n_0_527;
   wire n_0_528;
   wire n_0_529;
   wire n_0_530;
   wire n_0_531;
   wire n_0_532;
   wire n_0_533;
   wire n_0_534;
   wire n_0_535;
   wire n_0_536;
   wire n_0_537;
   wire n_0_538;
   wire n_0_539;
   wire n_0_540;
   wire n_0_541;
   wire n_0_542;
   wire n_0_543;
   wire n_0_0_35;
   wire n_0_480;
   wire n_0_481;
   wire n_0_482;
   wire n_0_483;
   wire n_0_484;
   wire n_0_485;
   wire n_0_486;
   wire n_0_487;
   wire n_0_488;
   wire n_0_489;
   wire n_0_490;
   wire n_0_491;
   wire n_0_492;
   wire n_0_493;
   wire n_0_494;
   wire n_0_495;
   wire n_0_496;
   wire n_0_497;
   wire n_0_498;
   wire n_0_499;
   wire n_0_500;
   wire n_0_501;
   wire n_0_502;
   wire n_0_503;
   wire n_0_504;
   wire n_0_505;
   wire n_0_506;
   wire n_0_507;
   wire n_0_508;
   wire n_0_509;
   wire n_0_510;
   wire n_0_511;
   wire n_0_0_36;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_0_37;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_0_38;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_0_39;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_0_40;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_0_41;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_0_42;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_0_43;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_0_44;
   wire n_0_574;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_0_54;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_0_55;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_0_56;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_0_57;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_0_58;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_192;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_33;
   wire n_0_0_32;
   wire n_0_0_0;
   wire n_0_30;
   wire n_0_0_64;
   wire n_0_32;
   wire n_0_0_65;
   wire [63:0]\c2[3] ;
   wire [63:0]\s2[3] ;
   wire [63:0]\c1[5] ;
   wire [63:0]\s1[5] ;
   wire [63:0]\c1[4] ;
   wire [63:0]\s1[4] ;
   wire [63:0]\c5[0] ;
   wire [63:0]\s5[0] ;
   wire [63:0]\c4[1] ;
   wire [63:0]\s4[1] ;
   wire [63:0]\c3[2] ;
   wire [63:0]\s3[2] ;
   wire [63:0]\c2[4] ;
   wire [63:0]\s2[4] ;
   wire [63:0]\c1[6] ;
   wire [63:0]\s1[6] ;
   wire [63:0]\c2[6] ;
   wire [63:0]\s2[6] ;
   wire [63:0]\c3[4] ;
   wire [63:0]\s3[4] ;
   wire [63:0]\c4[2] ;
   wire [63:0]\s4[2] ;
   wire [63:0]\c5[1] ;
   wire [63:0]\s5[1] ;
   wire [63:0]c6;
   wire [63:0]s6;
   wire [63:0]c7;
   wire [63:0]s7;
   wire [63:0]c8;
   wire [63:0]s8;
   wire [63:0]c9;
   wire [63:0]s9;
   wire [63:0]\c1[9] ;
   wire [63:0]\s1[9] ;

   CSA__1_2 A1_1 (.in1({n_0_30, uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, 
      uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, 
      uc_29, uc_30, uc_31, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, 
      n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, 
      n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, 
      n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_32}), .in2({n_0_32, uc_33, uc_34, 
      uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, 
      uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, uc_51, uc_52, uc_53, uc_54, 
      uc_55, uc_56, uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, uc_63, n_0_31, 
      n_0_573, n_0_572, n_0_571, n_0_570, n_0_569, n_0_568, n_0_567, n_0_566, 
      n_0_565, n_0_564, n_0_563, n_0_562, n_0_561, n_0_560, n_0_559, n_0_558, 
      n_0_557, n_0_556, n_0_555, n_0_554, n_0_553, n_0_552, n_0_551, n_0_550, 
      n_0_549, n_0_548, n_0_547, n_0_546, n_0_545, n_0_544, uc_64}), .in3({
      n_0_543, uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, uc_72, uc_73, 
      uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, uc_82, uc_83, 
      uc_84, uc_85, uc_86, uc_87, uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, 
      uc_94, n_0_542, n_0_541, n_0_540, n_0_539, n_0_538, n_0_537, n_0_536, 
      n_0_535, n_0_534, n_0_533, n_0_532, n_0_531, n_0_530, n_0_529, n_0_528, 
      n_0_527, n_0_526, n_0_525, n_0_524, n_0_523, n_0_522, n_0_521, n_0_520, 
      n_0_519, n_0_518, n_0_517, n_0_516, n_0_515, n_0_514, n_0_513, n_0_512, 
      uc_95, uc_96}), .sum({\s1[0] [33], uc_97, uc_98, uc_99, uc_100, uc_101, 
      uc_102, uc_103, uc_104, uc_105, uc_106, uc_107, uc_108, uc_109, uc_110, 
      uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, uc_117, uc_118, uc_119, 
      uc_120, uc_121, uc_122, uc_123, uc_124, uc_125, uc_126, \s1[0] [32], 
      \s1[0] [31], \s1[0] [30], \s1[0] [29], \s1[0] [28], \s1[0] [27], 
      \s1[0] [26], \s1[0] [25], \s1[0] [24], \s1[0] [23], \s1[0] [22], 
      \s1[0] [21], \s1[0] [20], \s1[0] [19], \s1[0] [18], \s1[0] [17], 
      \s1[0] [16], \s1[0] [15], \s1[0] [14], \s1[0] [13], \s1[0] [12], 
      \s1[0] [11], \s1[0] [10], \s1[0] [9], \s1[0] [8], \s1[0] [7], \s1[0] [6], 
      \s1[0] [5], \s1[0] [4], \s1[0] [3], \s1[0] [2], c[1], uc_127}), .c({
      \c1[0] [34], uc_128, uc_129, uc_130, uc_131, uc_132, uc_133, uc_134, 
      uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, uc_142, uc_143, 
      uc_144, uc_145, uc_146, uc_147, uc_148, uc_149, uc_150, uc_151, uc_152, 
      uc_153, uc_154, uc_155, uc_156, \c1[0] [33], \c1[0] [32], \c1[0] [31], 
      \c1[0] [30], \c1[0] [29], \c1[0] [28], \c1[0] [27], \c1[0] [26], 
      \c1[0] [25], \c1[0] [24], \c1[0] [23], \c1[0] [22], \c1[0] [21], 
      \c1[0] [20], \c1[0] [19], \c1[0] [18], \c1[0] [17], \c1[0] [16], 
      \c1[0] [15], \c1[0] [14], \c1[0] [13], \c1[0] [12], \c1[0] [11], 
      \c1[0] [10], \c1[0] [9], \c1[0] [8], \c1[0] [7], \c1[0] [6], \c1[0] [5], 
      \c1[0] [4], \c1[0] [3], \c1[0] [2], uc_157, uc_158}));
   CSA__1_5 A1_2 (.in1({n_0_511, uc_159, uc_160, uc_161, uc_162, uc_163, uc_164, 
      uc_165, uc_166, uc_167, uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, 
      uc_174, uc_175, uc_176, uc_177, uc_178, uc_179, uc_180, uc_181, uc_182, 
      uc_183, uc_184, uc_185, uc_186, uc_187, n_0_510, n_0_509, n_0_508, n_0_507, 
      n_0_506, n_0_505, n_0_504, n_0_503, n_0_502, n_0_501, n_0_500, n_0_499, 
      n_0_498, n_0_497, n_0_496, n_0_495, n_0_494, n_0_493, n_0_492, n_0_491, 
      n_0_490, n_0_489, n_0_488, n_0_487, n_0_486, n_0_485, n_0_484, n_0_483, 
      n_0_482, n_0_481, uc_188, uc_189, uc_190, uc_191}), .in2({n_0_479, uc_192, 
      uc_193, uc_194, uc_195, uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, 
      uc_202, uc_203, uc_204, uc_205, uc_206, uc_207, uc_208, uc_209, uc_210, 
      uc_211, uc_212, uc_213, uc_214, uc_215, uc_216, uc_217, uc_218, uc_219, 
      n_0_478, n_0_477, n_0_476, n_0_475, n_0_474, n_0_473, n_0_472, n_0_471, 
      n_0_470, n_0_469, n_0_468, n_0_467, n_0_466, n_0_465, n_0_464, n_0_463, 
      n_0_462, n_0_461, n_0_460, n_0_459, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, uc_220, 
      uc_221, uc_222, uc_223}), .in3({n_0_447, uc_224, uc_225, uc_226, uc_227, 
      uc_228, uc_229, uc_230, uc_231, uc_232, uc_233, uc_234, uc_235, uc_236, 
      uc_237, uc_238, uc_239, uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, 
      uc_246, uc_247, uc_248, uc_249, uc_250, n_0_446, n_0_445, n_0_444, n_0_443, 
      n_0_442, n_0_441, n_0_440, n_0_439, n_0_438, n_0_437, n_0_436, n_0_435, 
      n_0_434, n_0_433, n_0_432, n_0_431, n_0_430, n_0_429, n_0_428, n_0_427, 
      n_0_426, n_0_425, n_0_424, n_0_423, n_0_422, n_0_421, n_0_420, n_0_419, 
      n_0_418, n_0_417, n_0_416, uc_251, uc_252, uc_253, uc_254, uc_255}), 
      .sum({\s1[1] [36], uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, uc_262, 
      uc_263, uc_264, uc_265, uc_266, uc_267, uc_268, uc_269, uc_270, uc_271, 
      uc_272, uc_273, uc_274, uc_275, uc_276, uc_277, uc_278, uc_279, uc_280, 
      uc_281, uc_282, \s1[1] [35], \s1[1] [34], \s1[1] [33], \s1[1] [32], 
      \s1[1] [31], \s1[1] [30], \s1[1] [29], \s1[1] [28], \s1[1] [27], 
      \s1[1] [26], \s1[1] [25], \s1[1] [24], \s1[1] [23], \s1[1] [22], 
      \s1[1] [21], \s1[1] [20], \s1[1] [19], \s1[1] [18], \s1[1] [17], 
      \s1[1] [16], \s1[1] [15], \s1[1] [14], \s1[1] [13], \s1[1] [12], 
      \s1[1] [11], \s1[1] [10], \s1[1] [9], \s1[1] [8], \s1[1] [7], \s1[1] [6], 
      \s1[1] [5], \s1[1] [4], uc_283, uc_284, uc_285, uc_286}), .c({\c1[1] [37], 
      uc_287, uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, uc_294, uc_295, 
      uc_296, uc_297, uc_298, uc_299, uc_300, uc_301, uc_302, uc_303, uc_304, 
      uc_305, uc_306, uc_307, uc_308, uc_309, uc_310, uc_311, uc_312, 
      \c1[1] [36], \c1[1] [35], \c1[1] [34], \c1[1] [33], \c1[1] [32], 
      \c1[1] [31], \c1[1] [30], \c1[1] [29], \c1[1] [28], \c1[1] [27], 
      \c1[1] [26], \c1[1] [25], \c1[1] [24], \c1[1] [23], \c1[1] [22], 
      \c1[1] [21], \c1[1] [20], \c1[1] [19], \c1[1] [18], \c1[1] [17], 
      \c1[1] [16], \c1[1] [15], \c1[1] [14], \c1[1] [13], \c1[1] [12], 
      \c1[1] [11], \c1[1] [10], \c1[1] [9], \c1[1] [8], \c1[1] [7], \c1[1] [6], 
      \c1[1] [5], uc_313, uc_314, uc_315, uc_316, uc_317}));
   CSA__1_8 A2_1 (.in1({\s1[0] [33], uc_318, uc_319, uc_320, uc_321, uc_322, 
      uc_323, uc_324, uc_325, uc_326, uc_327, uc_328, uc_329, uc_330, uc_331, 
      uc_332, uc_333, uc_334, uc_335, uc_336, uc_337, uc_338, uc_339, uc_340, 
      uc_341, uc_342, uc_343, uc_344, uc_345, uc_346, uc_347, \s1[0] [32], 
      \s1[0] [31], \s1[0] [30], \s1[0] [29], \s1[0] [28], \s1[0] [27], 
      \s1[0] [26], \s1[0] [25], \s1[0] [24], \s1[0] [23], \s1[0] [22], 
      \s1[0] [21], \s1[0] [20], \s1[0] [19], \s1[0] [18], \s1[0] [17], 
      \s1[0] [16], \s1[0] [15], \s1[0] [14], \s1[0] [13], \s1[0] [12], 
      \s1[0] [11], \s1[0] [10], \s1[0] [9], \s1[0] [8], \s1[0] [7], \s1[0] [6], 
      \s1[0] [5], \s1[0] [4], \s1[0] [3], \s1[0] [2], uc_348, uc_349}), .in2({
      \c1[0] [34], uc_350, uc_351, uc_352, uc_353, uc_354, uc_355, uc_356, 
      uc_357, uc_358, uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, 
      uc_366, uc_367, uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, uc_374, 
      uc_375, uc_376, uc_377, uc_378, \c1[0] [33], \c1[0] [32], \c1[0] [31], 
      \c1[0] [30], \c1[0] [29], \c1[0] [28], \c1[0] [27], \c1[0] [26], 
      \c1[0] [25], \c1[0] [24], \c1[0] [23], \c1[0] [22], \c1[0] [21], 
      \c1[0] [20], \c1[0] [19], \c1[0] [18], \c1[0] [17], \c1[0] [16], 
      \c1[0] [15], \c1[0] [14], \c1[0] [13], \c1[0] [12], \c1[0] [11], 
      \c1[0] [10], \c1[0] [9], \c1[0] [8], \c1[0] [7], \c1[0] [6], \c1[0] [5], 
      \c1[0] [4], \c1[0] [3], \c1[0] [2], uc_379, uc_380}), .in3({\s1[1] [36], 
      uc_381, uc_382, uc_383, uc_384, uc_385, uc_386, uc_387, uc_388, uc_389, 
      uc_390, uc_391, uc_392, uc_393, uc_394, uc_395, uc_396, uc_397, uc_398, 
      uc_399, uc_400, uc_401, uc_402, uc_403, uc_404, uc_405, uc_406, uc_407, 
      \s1[1] [35], \s1[1] [34], \s1[1] [33], \s1[1] [32], \s1[1] [31], 
      \s1[1] [30], \s1[1] [29], \s1[1] [28], \s1[1] [27], \s1[1] [26], 
      \s1[1] [25], \s1[1] [24], \s1[1] [23], \s1[1] [22], \s1[1] [21], 
      \s1[1] [20], \s1[1] [19], \s1[1] [18], \s1[1] [17], \s1[1] [16], 
      \s1[1] [15], \s1[1] [14], \s1[1] [13], \s1[1] [12], \s1[1] [11], 
      \s1[1] [10], \s1[1] [9], \s1[1] [8], \s1[1] [7], \s1[1] [6], \s1[1] [5], 
      \s1[1] [4], n_0_480, uc_408, uc_409, uc_410}), .sum({\s2[0] [36], uc_411, 
      uc_412, uc_413, uc_414, uc_415, uc_416, uc_417, uc_418, uc_419, uc_420, 
      uc_421, uc_422, uc_423, uc_424, uc_425, uc_426, uc_427, uc_428, uc_429, 
      uc_430, uc_431, uc_432, uc_433, uc_434, uc_435, uc_436, uc_437, 
      \s2[0] [35], \s2[0] [34], \s2[0] [33], \s2[0] [32], \s2[0] [31], 
      \s2[0] [30], \s2[0] [29], \s2[0] [28], \s2[0] [27], \s2[0] [26], 
      \s2[0] [25], \s2[0] [24], \s2[0] [23], \s2[0] [22], \s2[0] [21], 
      \s2[0] [20], \s2[0] [19], \s2[0] [18], \s2[0] [17], \s2[0] [16], 
      \s2[0] [15], \s2[0] [14], \s2[0] [13], \s2[0] [12], \s2[0] [11], 
      \s2[0] [10], \s2[0] [9], \s2[0] [8], \s2[0] [7], \s2[0] [6], \s2[0] [5], 
      \s2[0] [4], \s2[0] [3], c[2], uc_438, uc_439}), .c({\c2[0] [37], uc_440, 
      uc_441, uc_442, uc_443, uc_444, uc_445, uc_446, uc_447, uc_448, uc_449, 
      uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, 
      uc_459, uc_460, uc_461, uc_462, uc_463, uc_464, uc_465, \c2[0] [36], 
      \c2[0] [35], \c2[0] [34], \c2[0] [33], \c2[0] [32], \c2[0] [31], 
      \c2[0] [30], \c2[0] [29], \c2[0] [28], \c2[0] [27], \c2[0] [26], 
      \c2[0] [25], \c2[0] [24], \c2[0] [23], \c2[0] [22], \c2[0] [21], 
      \c2[0] [20], \c2[0] [19], \c2[0] [18], \c2[0] [17], \c2[0] [16], 
      \c2[0] [15], \c2[0] [14], \c2[0] [13], \c2[0] [12], \c2[0] [11], 
      \c2[0] [10], \c2[0] [9], \c2[0] [8], \c2[0] [7], \c2[0] [6], \c2[0] [5], 
      \c2[0] [4], \c2[0] [3], uc_466, uc_467, uc_468}));
   CSA__1_11 A1_3 (.in1({n_0_415, uc_469, uc_470, uc_471, uc_472, uc_473, uc_474, 
      uc_475, uc_476, uc_477, uc_478, uc_479, uc_480, uc_481, uc_482, uc_483, 
      uc_484, uc_485, uc_486, uc_487, uc_488, uc_489, uc_490, uc_491, uc_492, 
      uc_493, uc_494, n_0_414, n_0_413, n_0_412, n_0_411, n_0_410, n_0_409, 
      n_0_408, n_0_407, n_0_406, n_0_405, n_0_404, n_0_403, n_0_402, n_0_401, 
      n_0_400, n_0_399, n_0_398, n_0_397, n_0_396, n_0_395, n_0_394, n_0_393, 
      n_0_392, n_0_391, n_0_390, n_0_389, n_0_388, n_0_387, n_0_386, n_0_385, 
      uc_495, uc_496, uc_497, uc_498, uc_499, uc_500, uc_501}), .in2({n_0_383, 
      uc_502, uc_503, uc_504, uc_505, uc_506, uc_507, uc_508, uc_509, uc_510, 
      uc_511, uc_512, uc_513, uc_514, uc_515, uc_516, uc_517, uc_518, uc_519, 
      uc_520, uc_521, uc_522, uc_523, uc_524, uc_525, uc_526, n_0_382, n_0_381, 
      n_0_380, n_0_379, n_0_378, n_0_377, n_0_376, n_0_375, n_0_374, n_0_373, 
      n_0_372, n_0_371, n_0_370, n_0_369, n_0_368, n_0_367, n_0_366, n_0_365, 
      n_0_364, n_0_363, n_0_362, n_0_361, n_0_360, n_0_359, n_0_358, n_0_357, 
      n_0_356, n_0_355, n_0_354, n_0_353, n_0_352, uc_527, uc_528, uc_529, 
      uc_530, uc_531, uc_532, uc_533}), .in3({n_0_351, uc_534, uc_535, uc_536, 
      uc_537, uc_538, uc_539, uc_540, uc_541, uc_542, uc_543, uc_544, uc_545, 
      uc_546, uc_547, uc_548, uc_549, uc_550, uc_551, uc_552, uc_553, uc_554, 
      uc_555, uc_556, uc_557, n_0_350, n_0_349, n_0_348, n_0_347, n_0_346, 
      n_0_345, n_0_344, n_0_343, n_0_342, n_0_341, n_0_340, n_0_339, n_0_338, 
      n_0_337, n_0_336, n_0_335, n_0_334, n_0_333, n_0_332, n_0_331, n_0_330, 
      n_0_329, n_0_328, n_0_327, n_0_326, n_0_325, n_0_324, n_0_323, n_0_322, 
      n_0_321, n_0_320, uc_558, uc_559, uc_560, uc_561, uc_562, uc_563, uc_564, 
      uc_565}), .sum({\s1[2] [39], uc_566, uc_567, uc_568, uc_569, uc_570, 
      uc_571, uc_572, uc_573, uc_574, uc_575, uc_576, uc_577, uc_578, uc_579, 
      uc_580, uc_581, uc_582, uc_583, uc_584, uc_585, uc_586, uc_587, uc_588, 
      uc_589, \s1[2] [38], \s1[2] [37], \s1[2] [36], \s1[2] [35], \s1[2] [34], 
      \s1[2] [33], \s1[2] [32], \s1[2] [31], \s1[2] [30], \s1[2] [29], 
      \s1[2] [28], \s1[2] [27], \s1[2] [26], \s1[2] [25], \s1[2] [24], 
      \s1[2] [23], \s1[2] [22], \s1[2] [21], \s1[2] [20], \s1[2] [19], 
      \s1[2] [18], \s1[2] [17], \s1[2] [16], \s1[2] [15], \s1[2] [14], 
      \s1[2] [13], \s1[2] [12], \s1[2] [11], \s1[2] [10], \s1[2] [9], \s1[2] [8], 
      \s1[2] [7], uc_590, uc_591, uc_592, uc_593, uc_594, uc_595, uc_596}), 
      .c({\c1[2] [40], uc_597, uc_598, uc_599, uc_600, uc_601, uc_602, uc_603, 
      uc_604, uc_605, uc_606, uc_607, uc_608, uc_609, uc_610, uc_611, uc_612, 
      uc_613, uc_614, uc_615, uc_616, uc_617, uc_618, uc_619, \c1[2] [39], 
      \c1[2] [38], \c1[2] [37], \c1[2] [36], \c1[2] [35], \c1[2] [34], 
      \c1[2] [33], \c1[2] [32], \c1[2] [31], \c1[2] [30], \c1[2] [29], 
      \c1[2] [28], \c1[2] [27], \c1[2] [26], \c1[2] [25], \c1[2] [24], 
      \c1[2] [23], \c1[2] [22], \c1[2] [21], \c1[2] [20], \c1[2] [19], 
      \c1[2] [18], \c1[2] [17], \c1[2] [16], \c1[2] [15], \c1[2] [14], 
      \c1[2] [13], \c1[2] [12], \c1[2] [11], \c1[2] [10], \c1[2] [9], \c1[2] [8], 
      uc_620, uc_621, uc_622, uc_623, uc_624, uc_625, uc_626, uc_627}));
   CSA__1_14 A2_2 (.in1({\c1[1] [37], uc_628, uc_629, uc_630, uc_631, uc_632, 
      uc_633, uc_634, uc_635, uc_636, uc_637, uc_638, uc_639, uc_640, uc_641, 
      uc_642, uc_643, uc_644, uc_645, uc_646, uc_647, uc_648, uc_649, uc_650, 
      uc_651, uc_652, uc_653, \c1[1] [36], \c1[1] [35], \c1[1] [34], \c1[1] [33], 
      \c1[1] [32], \c1[1] [31], \c1[1] [30], \c1[1] [29], \c1[1] [28], 
      \c1[1] [27], \c1[1] [26], \c1[1] [25], \c1[1] [24], \c1[1] [23], 
      \c1[1] [22], \c1[1] [21], \c1[1] [20], \c1[1] [19], \c1[1] [18], 
      \c1[1] [17], \c1[1] [16], \c1[1] [15], \c1[1] [14], \c1[1] [13], 
      \c1[1] [12], \c1[1] [11], \c1[1] [10], \c1[1] [9], \c1[1] [8], \c1[1] [7], 
      \c1[1] [6], uc_654, uc_655, uc_656, uc_657, uc_658, uc_659}), .in2({
      \s1[2] [39], uc_660, uc_661, uc_662, uc_663, uc_664, uc_665, uc_666, 
      uc_667, uc_668, uc_669, uc_670, uc_671, uc_672, uc_673, uc_674, uc_675, 
      uc_676, uc_677, uc_678, uc_679, uc_680, uc_681, uc_682, uc_683, 
      \s1[2] [38], \s1[2] [37], \s1[2] [36], \s1[2] [35], \s1[2] [34], 
      \s1[2] [33], \s1[2] [32], \s1[2] [31], \s1[2] [30], \s1[2] [29], 
      \s1[2] [28], \s1[2] [27], \s1[2] [26], \s1[2] [25], \s1[2] [24], 
      \s1[2] [23], \s1[2] [22], \s1[2] [21], \s1[2] [20], \s1[2] [19], 
      \s1[2] [18], \s1[2] [17], \s1[2] [16], \s1[2] [15], \s1[2] [14], 
      \s1[2] [13], \s1[2] [12], \s1[2] [11], \s1[2] [10], \s1[2] [9], \s1[2] [8], 
      \s1[2] [7], n_0_384, uc_684, uc_685, uc_686, uc_687, uc_688, uc_689}), 
      .in3({\c1[2] [40], uc_690, uc_691, uc_692, uc_693, uc_694, uc_695, uc_696, 
      uc_697, uc_698, uc_699, uc_700, uc_701, uc_702, uc_703, uc_704, uc_705, 
      uc_706, uc_707, uc_708, uc_709, uc_710, uc_711, uc_712, \c1[2] [39], 
      \c1[2] [38], \c1[2] [37], \c1[2] [36], \c1[2] [35], \c1[2] [34], 
      \c1[2] [33], \c1[2] [32], \c1[2] [31], \c1[2] [30], \c1[2] [29], 
      \c1[2] [28], \c1[2] [27], \c1[2] [26], \c1[2] [25], \c1[2] [24], 
      \c1[2] [23], \c1[2] [22], \c1[2] [21], \c1[2] [20], \c1[2] [19], 
      \c1[2] [18], \c1[2] [17], \c1[2] [16], \c1[2] [15], \c1[2] [14], 
      \c1[2] [13], \c1[2] [12], \c1[2] [11], \c1[2] [10], \c1[2] [9], \c1[2] [8], 
      uc_713, uc_714, uc_715, uc_716, uc_717, uc_718, uc_719, uc_720}), .sum({
      \s2[1] [40], uc_721, uc_722, uc_723, uc_724, uc_725, uc_726, uc_727, 
      uc_728, uc_729, uc_730, uc_731, uc_732, uc_733, uc_734, uc_735, uc_736, 
      uc_737, uc_738, uc_739, uc_740, uc_741, uc_742, uc_743, \s2[1] [39], 
      \s2[1] [38], \s2[1] [37], \s2[1] [36], \s2[1] [35], \s2[1] [34], 
      \s2[1] [33], \s2[1] [32], \s2[1] [31], \s2[1] [30], \s2[1] [29], 
      \s2[1] [28], \s2[1] [27], \s2[1] [26], \s2[1] [25], \s2[1] [24], 
      \s2[1] [23], \s2[1] [22], \s2[1] [21], \s2[1] [20], \s2[1] [19], 
      \s2[1] [18], \s2[1] [17], \s2[1] [16], \s2[1] [15], \s2[1] [14], 
      \s2[1] [13], \s2[1] [12], \s2[1] [11], \s2[1] [10], \s2[1] [9], \s2[1] [8], 
      \s2[1] [7], \s2[1] [6], uc_744, uc_745, uc_746, uc_747, uc_748, uc_749}), 
      .c({\c2[1] [41], uc_750, uc_751, uc_752, uc_753, uc_754, uc_755, uc_756, 
      uc_757, uc_758, uc_759, uc_760, uc_761, uc_762, uc_763, uc_764, uc_765, 
      uc_766, uc_767, uc_768, uc_769, uc_770, uc_771, \c2[1] [40], \c2[1] [39], 
      \c2[1] [38], \c2[1] [37], \c2[1] [36], \c2[1] [35], \c2[1] [34], 
      \c2[1] [33], \c2[1] [32], \c2[1] [31], \c2[1] [30], \c2[1] [29], 
      \c2[1] [28], \c2[1] [27], \c2[1] [26], \c2[1] [25], \c2[1] [24], 
      \c2[1] [23], \c2[1] [22], \c2[1] [21], \c2[1] [20], \c2[1] [19], 
      \c2[1] [18], \c2[1] [17], \c2[1] [16], \c2[1] [15], \c2[1] [14], 
      \c2[1] [13], \c2[1] [12], \c2[1] [11], \c2[1] [10], \c2[1] [9], \c2[1] [8], 
      \c2[1] [7], uc_772, uc_773, uc_774, uc_775, uc_776, uc_777, uc_778}));
   CSA__1_17 A3_1 (.in1({\s2[0] [36], uc_779, uc_780, uc_781, uc_782, uc_783, 
      uc_784, uc_785, uc_786, uc_787, uc_788, uc_789, uc_790, uc_791, uc_792, 
      uc_793, uc_794, uc_795, uc_796, uc_797, uc_798, uc_799, uc_800, uc_801, 
      uc_802, uc_803, uc_804, uc_805, \s2[0] [35], \s2[0] [34], \s2[0] [33], 
      \s2[0] [32], \s2[0] [31], \s2[0] [30], \s2[0] [29], \s2[0] [28], 
      \s2[0] [27], \s2[0] [26], \s2[0] [25], \s2[0] [24], \s2[0] [23], 
      \s2[0] [22], \s2[0] [21], \s2[0] [20], \s2[0] [19], \s2[0] [18], 
      \s2[0] [17], \s2[0] [16], \s2[0] [15], \s2[0] [14], \s2[0] [13], 
      \s2[0] [12], \s2[0] [11], \s2[0] [10], \s2[0] [9], \s2[0] [8], \s2[0] [7], 
      \s2[0] [6], \s2[0] [5], \s2[0] [4], \s2[0] [3], uc_806, uc_807, uc_808}), 
      .in2({\c2[0] [37], uc_809, uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, 
      uc_816, uc_817, uc_818, uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, 
      uc_825, uc_826, uc_827, uc_828, uc_829, uc_830, uc_831, uc_832, uc_833, 
      uc_834, \c2[0] [36], \c2[0] [35], \c2[0] [34], \c2[0] [33], \c2[0] [32], 
      \c2[0] [31], \c2[0] [30], \c2[0] [29], \c2[0] [28], \c2[0] [27], 
      \c2[0] [26], \c2[0] [25], \c2[0] [24], \c2[0] [23], \c2[0] [22], 
      \c2[0] [21], \c2[0] [20], \c2[0] [19], \c2[0] [18], \c2[0] [17], 
      \c2[0] [16], \c2[0] [15], \c2[0] [14], \c2[0] [13], \c2[0] [12], 
      \c2[0] [11], \c2[0] [10], \c2[0] [9], \c2[0] [8], \c2[0] [7], \c2[0] [6], 
      \c2[0] [5], \c2[0] [4], \c2[0] [3], uc_835, uc_836, uc_837}), .in3({
      \s2[1] [40], uc_838, uc_839, uc_840, uc_841, uc_842, uc_843, uc_844, 
      uc_845, uc_846, uc_847, uc_848, uc_849, uc_850, uc_851, uc_852, uc_853, 
      uc_854, uc_855, uc_856, uc_857, uc_858, uc_859, uc_860, \s2[1] [39], 
      \s2[1] [38], \s2[1] [37], \s2[1] [36], \s2[1] [35], \s2[1] [34], 
      \s2[1] [33], \s2[1] [32], \s2[1] [31], \s2[1] [30], \s2[1] [29], 
      \s2[1] [28], \s2[1] [27], \s2[1] [26], \s2[1] [25], \s2[1] [24], 
      \s2[1] [23], \s2[1] [22], \s2[1] [21], \s2[1] [20], \s2[1] [19], 
      \s2[1] [18], \s2[1] [17], \s2[1] [16], \s2[1] [15], \s2[1] [14], 
      \s2[1] [13], \s2[1] [12], \s2[1] [11], \s2[1] [10], \s2[1] [9], \s2[1] [8], 
      \s2[1] [7], \s2[1] [6], \c1[1] [5], uc_861, uc_862, uc_863, uc_864, uc_865}), 
      .sum({\s3[0] [40], uc_866, uc_867, uc_868, uc_869, uc_870, uc_871, uc_872, 
      uc_873, uc_874, uc_875, uc_876, uc_877, uc_878, uc_879, uc_880, uc_881, 
      uc_882, uc_883, uc_884, uc_885, uc_886, uc_887, uc_888, \s3[0] [39], 
      \s3[0] [38], \s3[0] [37], \s3[0] [36], \s3[0] [35], \s3[0] [34], 
      \s3[0] [33], \s3[0] [32], \s3[0] [31], \s3[0] [30], \s3[0] [29], 
      \s3[0] [28], \s3[0] [27], \s3[0] [26], \s3[0] [25], \s3[0] [24], 
      \s3[0] [23], \s3[0] [22], \s3[0] [21], \s3[0] [20], \s3[0] [19], 
      \s3[0] [18], \s3[0] [17], \s3[0] [16], \s3[0] [15], \s3[0] [14], 
      \s3[0] [13], \s3[0] [12], \s3[0] [11], \s3[0] [10], \s3[0] [9], \s3[0] [8], 
      \s3[0] [7], \s3[0] [6], \s3[0] [5], \s3[0] [4], c[3], uc_889, uc_890, 
      uc_891}), .c({\c3[0] [41], uc_892, uc_893, uc_894, uc_895, uc_896, uc_897, 
      uc_898, uc_899, uc_900, uc_901, uc_902, uc_903, uc_904, uc_905, uc_906, 
      uc_907, uc_908, uc_909, uc_910, uc_911, uc_912, uc_913, \c3[0] [40], 
      \c3[0] [39], \c3[0] [38], \c3[0] [37], \c3[0] [36], \c3[0] [35], 
      \c3[0] [34], \c3[0] [33], \c3[0] [32], \c3[0] [31], \c3[0] [30], 
      \c3[0] [29], \c3[0] [28], \c3[0] [27], \c3[0] [26], \c3[0] [25], 
      \c3[0] [24], \c3[0] [23], \c3[0] [22], \c3[0] [21], \c3[0] [20], 
      \c3[0] [19], \c3[0] [18], \c3[0] [17], \c3[0] [16], \c3[0] [15], 
      \c3[0] [14], \c3[0] [13], \c3[0] [12], \c3[0] [11], \c3[0] [10], 
      \c3[0] [9], \c3[0] [8], \c3[0] [7], \c3[0] [6], \c3[0] [5], \c3[0] [4], 
      uc_914, uc_915, uc_916, uc_917}));
   CSA__1_20 A1_4 (.in1({n_0_319, uc_918, uc_919, uc_920, uc_921, uc_922, uc_923, 
      uc_924, uc_925, uc_926, uc_927, uc_928, uc_929, uc_930, uc_931, uc_932, 
      uc_933, uc_934, uc_935, uc_936, uc_937, uc_938, uc_939, uc_940, n_0_318, 
      n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, n_0_312, n_0_311, n_0_310, 
      n_0_309, n_0_308, n_0_307, n_0_306, n_0_305, n_0_304, n_0_303, n_0_302, 
      n_0_301, n_0_300, n_0_299, n_0_298, n_0_297, n_0_296, n_0_295, n_0_294, 
      n_0_293, n_0_292, n_0_291, n_0_290, n_0_289, uc_941, uc_942, uc_943, 
      uc_944, uc_945, uc_946, uc_947, uc_948, uc_949, uc_950}), .in2({n_0_287, 
      uc_951, uc_952, uc_953, uc_954, uc_955, uc_956, uc_957, uc_958, uc_959, 
      uc_960, uc_961, uc_962, uc_963, uc_964, uc_965, uc_966, uc_967, uc_968, 
      uc_969, uc_970, uc_971, uc_972, n_0_286, n_0_285, n_0_284, n_0_283, 
      n_0_282, n_0_281, n_0_280, n_0_279, n_0_278, n_0_277, n_0_276, n_0_275, 
      n_0_274, n_0_273, n_0_272, n_0_271, n_0_270, n_0_269, n_0_268, n_0_267, 
      n_0_266, n_0_265, n_0_264, n_0_263, n_0_262, n_0_261, n_0_260, n_0_259, 
      n_0_258, n_0_257, n_0_256, uc_973, uc_974, uc_975, uc_976, uc_977, uc_978, 
      uc_979, uc_980, uc_981, uc_982}), .in3({n_0_255, uc_983, uc_984, uc_985, 
      uc_986, uc_987, uc_988, uc_989, uc_990, uc_991, uc_992, uc_993, uc_994, 
      uc_995, uc_996, uc_997, uc_998, uc_999, uc_1000, uc_1001, uc_1002, uc_1003, 
      n_0_254, n_0_253, n_0_252, n_0_251, n_0_250, n_0_249, n_0_248, n_0_247, 
      n_0_246, n_0_245, n_0_244, n_0_243, n_0_242, n_0_241, n_0_240, n_0_239, 
      n_0_238, n_0_237, n_0_236, n_0_235, n_0_234, n_0_233, n_0_232, n_0_231, 
      n_0_230, n_0_229, n_0_228, n_0_227, n_0_226, n_0_225, n_0_224, uc_1004, 
      uc_1005, uc_1006, uc_1007, uc_1008, uc_1009, uc_1010, uc_1011, uc_1012, 
      uc_1013, uc_1014}), .sum({\s1[3] [42], uc_1015, uc_1016, uc_1017, uc_1018, 
      uc_1019, uc_1020, uc_1021, uc_1022, uc_1023, uc_1024, uc_1025, uc_1026, 
      uc_1027, uc_1028, uc_1029, uc_1030, uc_1031, uc_1032, uc_1033, uc_1034, 
      uc_1035, \s1[3] [41], \s1[3] [40], \s1[3] [39], \s1[3] [38], \s1[3] [37], 
      \s1[3] [36], \s1[3] [35], \s1[3] [34], \s1[3] [33], \s1[3] [32], 
      \s1[3] [31], \s1[3] [30], \s1[3] [29], \s1[3] [28], \s1[3] [27], 
      \s1[3] [26], \s1[3] [25], \s1[3] [24], \s1[3] [23], \s1[3] [22], 
      \s1[3] [21], \s1[3] [20], \s1[3] [19], \s1[3] [18], \s1[3] [17], 
      \s1[3] [16], \s1[3] [15], \s1[3] [14], \s1[3] [13], \s1[3] [12], 
      \s1[3] [11], \s1[3] [10], uc_1036, uc_1037, uc_1038, uc_1039, uc_1040, 
      uc_1041, uc_1042, uc_1043, uc_1044, uc_1045}), .c({\c1[3] [43], uc_1046, 
      uc_1047, uc_1048, uc_1049, uc_1050, uc_1051, uc_1052, uc_1053, uc_1054, 
      uc_1055, uc_1056, uc_1057, uc_1058, uc_1059, uc_1060, uc_1061, uc_1062, 
      uc_1063, uc_1064, uc_1065, \c1[3] [42], \c1[3] [41], \c1[3] [40], 
      \c1[3] [39], \c1[3] [38], \c1[3] [37], \c1[3] [36], \c1[3] [35], 
      \c1[3] [34], \c1[3] [33], \c1[3] [32], \c1[3] [31], \c1[3] [30], 
      \c1[3] [29], \c1[3] [28], \c1[3] [27], \c1[3] [26], \c1[3] [25], 
      \c1[3] [24], \c1[3] [23], \c1[3] [22], \c1[3] [21], \c1[3] [20], 
      \c1[3] [19], \c1[3] [18], \c1[3] [17], \c1[3] [16], \c1[3] [15], 
      \c1[3] [14], \c1[3] [13], \c1[3] [12], \c1[3] [11], uc_1066, uc_1067, 
      uc_1068, uc_1069, uc_1070, uc_1071, uc_1072, uc_1073, uc_1074, uc_1075, 
      uc_1076}));
   CSA__1_23 A1_9 (.in1({n_0_127, uc_1077, uc_1078, uc_1079, uc_1080, uc_1081, 
      uc_1082, uc_1083, uc_1084, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, 
      n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, 
      n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, 
      n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, 
      n_0_97, uc_1085, uc_1086, uc_1087, uc_1088, uc_1089, uc_1090, uc_1091, 
      uc_1092, uc_1093, uc_1094, uc_1095, uc_1096, uc_1097, uc_1098, uc_1099, 
      uc_1100, uc_1101, uc_1102, uc_1103, uc_1104, uc_1105, uc_1106, uc_1107, 
      uc_1108, uc_1109}), .in2({n_0_95, uc_1110, uc_1111, uc_1112, uc_1113, 
      uc_1114, uc_1115, uc_1116, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, 
      n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, 
      n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, 
      n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, uc_1117, uc_1118, 
      uc_1119, uc_1120, uc_1121, uc_1122, uc_1123, uc_1124, uc_1125, uc_1126, 
      uc_1127, uc_1128, uc_1129, uc_1130, uc_1131, uc_1132, uc_1133, uc_1134, 
      uc_1135, uc_1136, uc_1137, uc_1138, uc_1139, uc_1140, uc_1141}), .in3({
      n_0_192, uc_1142, uc_1143, uc_1144, uc_1145, uc_1146, uc_1147, n_0_63, 
      n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, 
      n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, 
      n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, 
      n_0_35, n_0_34, n_0_33, uc_1148, uc_1149, uc_1150, uc_1151, uc_1152, 
      uc_1153, uc_1154, uc_1155, uc_1156, uc_1157, uc_1158, uc_1159, uc_1160, 
      uc_1161, uc_1162, uc_1163, uc_1164, uc_1165, uc_1166, uc_1167, uc_1168, 
      uc_1169, uc_1170, uc_1171, uc_1172, uc_1173}), .sum({\s1[8] [57], uc_1174, 
      uc_1175, uc_1176, uc_1177, uc_1178, uc_1179, \s1[8] [56], \s1[8] [55], 
      \s1[8] [54], \s1[8] [53], \s1[8] [52], \s1[8] [51], \s1[8] [50], 
      \s1[8] [49], \s1[8] [48], \s1[8] [47], \s1[8] [46], \s1[8] [45], 
      \s1[8] [44], \s1[8] [43], \s1[8] [42], \s1[8] [41], \s1[8] [40], 
      \s1[8] [39], \s1[8] [38], \s1[8] [37], \s1[8] [36], \s1[8] [35], 
      \s1[8] [34], \s1[8] [33], \s1[8] [32], \s1[8] [31], \s1[8] [30], 
      \s1[8] [29], \s1[8] [28], \s1[8] [27], \s1[8] [26], \s1[8] [25], uc_1180, 
      uc_1181, uc_1182, uc_1183, uc_1184, uc_1185, uc_1186, uc_1187, uc_1188, 
      uc_1189, uc_1190, uc_1191, uc_1192, uc_1193, uc_1194, uc_1195, uc_1196, 
      uc_1197, uc_1198, uc_1199, uc_1200, uc_1201, uc_1202, uc_1203, uc_1204}), 
      .c({\c1[8] [58], uc_1205, uc_1206, uc_1207, uc_1208, uc_1209, \c1[8] [57], 
      \c1[8] [56], \c1[8] [55], \c1[8] [54], \c1[8] [53], \c1[8] [52], 
      \c1[8] [51], \c1[8] [50], \c1[8] [49], \c1[8] [48], \c1[8] [47], 
      \c1[8] [46], \c1[8] [45], \c1[8] [44], \c1[8] [43], \c1[8] [42], 
      \c1[8] [41], \c1[8] [40], \c1[8] [39], \c1[8] [38], \c1[8] [37], 
      \c1[8] [36], \c1[8] [35], \c1[8] [34], \c1[8] [33], \c1[8] [32], 
      \c1[8] [31], \c1[8] [30], \c1[8] [29], \c1[8] [28], \c1[8] [27], 
      \c1[8] [26], uc_1210, uc_1211, uc_1212, uc_1213, uc_1214, uc_1215, uc_1216, 
      uc_1217, uc_1218, uc_1219, uc_1220, uc_1221, uc_1222, uc_1223, uc_1224, 
      uc_1225, uc_1226, uc_1227, uc_1228, uc_1229, uc_1230, uc_1231, uc_1232, 
      uc_1233, uc_1234, uc_1235}));
   CSA__1_26 A2_3 (.in1({\s1[3] [42], uc_1236, uc_1237, uc_1238, uc_1239, 
      uc_1240, uc_1241, uc_1242, uc_1243, uc_1244, uc_1245, uc_1246, uc_1247, 
      uc_1248, uc_1249, uc_1250, uc_1251, uc_1252, uc_1253, uc_1254, uc_1255, 
      uc_1256, \s1[3] [41], \s1[3] [40], \s1[3] [39], \s1[3] [38], \s1[3] [37], 
      \s1[3] [36], \s1[3] [35], \s1[3] [34], \s1[3] [33], \s1[3] [32], 
      \s1[3] [31], \s1[3] [30], \s1[3] [29], \s1[3] [28], \s1[3] [27], 
      \s1[3] [26], \s1[3] [25], \s1[3] [24], \s1[3] [23], \s1[3] [22], 
      \s1[3] [21], \s1[3] [20], \s1[3] [19], \s1[3] [18], \s1[3] [17], 
      \s1[3] [16], \s1[3] [15], \s1[3] [14], \s1[3] [13], \s1[3] [12], 
      \s1[3] [11], uc_1257, uc_1258, uc_1259, uc_1260, uc_1261, uc_1262, uc_1263, 
      uc_1264, uc_1265, uc_1266, uc_1267}), .in2({\c1[3] [43], uc_1268, uc_1269, 
      uc_1270, uc_1271, uc_1272, uc_1273, uc_1274, uc_1275, uc_1276, uc_1277, 
      uc_1278, uc_1279, uc_1280, uc_1281, uc_1282, uc_1283, uc_1284, uc_1285, 
      uc_1286, uc_1287, \c1[3] [42], \c1[3] [41], \c1[3] [40], \c1[3] [39], 
      \c1[3] [38], \c1[3] [37], \c1[3] [36], \c1[3] [35], \c1[3] [34], 
      \c1[3] [33], \c1[3] [32], \c1[3] [31], \c1[3] [30], \c1[3] [29], 
      \c1[3] [28], \c1[3] [27], \c1[3] [26], \c1[3] [25], \c1[3] [24], 
      \c1[3] [23], \c1[3] [22], \c1[3] [21], \c1[3] [20], \c1[3] [19], 
      \c1[3] [18], \c1[3] [17], \c1[3] [16], \c1[3] [15], \c1[3] [14], 
      \c1[3] [13], \c1[3] [12], \c1[3] [11], uc_1288, uc_1289, uc_1290, uc_1291, 
      uc_1292, uc_1293, uc_1294, uc_1295, uc_1296, uc_1297, uc_1298}), .in3({
      \s1[4] [45], uc_1299, uc_1300, uc_1301, uc_1302, uc_1303, uc_1304, uc_1305, 
      uc_1306, uc_1307, uc_1308, uc_1309, uc_1310, uc_1311, uc_1312, uc_1313, 
      uc_1314, uc_1315, uc_1316, \s1[4] [44], \s1[4] [43], \s1[4] [42], 
      \s1[4] [41], \s1[4] [40], \s1[4] [39], \s1[4] [38], \s1[4] [37], 
      \s1[4] [36], \s1[4] [35], \s1[4] [34], \s1[4] [33], \s1[4] [32], 
      \s1[4] [31], \s1[4] [30], \s1[4] [29], \s1[4] [28], \s1[4] [27], 
      \s1[4] [26], \s1[4] [25], \s1[4] [24], \s1[4] [23], \s1[4] [22], 
      \s1[4] [21], \s1[4] [20], \s1[4] [19], \s1[4] [18], \s1[4] [17], 
      \s1[4] [16], \s1[4] [15], \s1[4] [14], \s1[4] [13], n_0_574, uc_1317, 
      uc_1318, uc_1319, uc_1320, uc_1321, uc_1322, uc_1323, uc_1324, uc_1325, 
      uc_1326, uc_1327, uc_1328}), .sum({\s2[2] [45], uc_1329, uc_1330, uc_1331, 
      uc_1332, uc_1333, uc_1334, uc_1335, uc_1336, uc_1337, uc_1338, uc_1339, 
      uc_1340, uc_1341, uc_1342, uc_1343, uc_1344, uc_1345, uc_1346, \s2[2] [44], 
      \s2[2] [43], \s2[2] [42], \s2[2] [41], \s2[2] [40], \s2[2] [39], 
      \s2[2] [38], \s2[2] [37], \s2[2] [36], \s2[2] [35], \s2[2] [34], 
      \s2[2] [33], \s2[2] [32], \s2[2] [31], \s2[2] [30], \s2[2] [29], 
      \s2[2] [28], \s2[2] [27], \s2[2] [26], \s2[2] [25], \s2[2] [24], 
      \s2[2] [23], \s2[2] [22], \s2[2] [21], \s2[2] [20], \s2[2] [19], 
      \s2[2] [18], \s2[2] [17], \s2[2] [16], \s2[2] [15], \s2[2] [14], 
      \s2[2] [13], \s2[2] [12], \s2[2] [11], uc_1347, uc_1348, uc_1349, uc_1350, 
      uc_1351, uc_1352, uc_1353, uc_1354, uc_1355, uc_1356, uc_1357}), .c({
      \c2[2] [46], uc_1358, uc_1359, uc_1360, uc_1361, uc_1362, uc_1363, uc_1364, 
      uc_1365, uc_1366, uc_1367, uc_1368, uc_1369, uc_1370, uc_1371, uc_1372, 
      uc_1373, uc_1374, \c2[2] [45], \c2[2] [44], \c2[2] [43], \c2[2] [42], 
      \c2[2] [41], \c2[2] [40], \c2[2] [39], \c2[2] [38], \c2[2] [37], 
      \c2[2] [36], \c2[2] [35], \c2[2] [34], \c2[2] [33], \c2[2] [32], 
      \c2[2] [31], \c2[2] [30], \c2[2] [29], \c2[2] [28], \c2[2] [27], 
      \c2[2] [26], \c2[2] [25], \c2[2] [24], \c2[2] [23], \c2[2] [22], 
      \c2[2] [21], \c2[2] [20], \c2[2] [19], \c2[2] [18], \c2[2] [17], 
      \c2[2] [16], \c2[2] [15], \c2[2] [14], \c2[2] [13], \c2[2] [12], uc_1375, 
      uc_1376, uc_1377, uc_1378, uc_1379, uc_1380, uc_1381, uc_1382, uc_1383, 
      uc_1384, uc_1385, uc_1386}));
   CSA__1_29 A3_2 (.in1({\c2[1] [41], uc_1387, uc_1388, uc_1389, uc_1390, 
      uc_1391, uc_1392, uc_1393, uc_1394, uc_1395, uc_1396, uc_1397, uc_1398, 
      uc_1399, uc_1400, uc_1401, uc_1402, uc_1403, uc_1404, uc_1405, uc_1406, 
      uc_1407, uc_1408, \c2[1] [40], \c2[1] [39], \c2[1] [38], \c2[1] [37], 
      \c2[1] [36], \c2[1] [35], \c2[1] [34], \c2[1] [33], \c2[1] [32], 
      \c2[1] [31], \c2[1] [30], \c2[1] [29], \c2[1] [28], \c2[1] [27], 
      \c2[1] [26], \c2[1] [25], \c2[1] [24], \c2[1] [23], \c2[1] [22], 
      \c2[1] [21], \c2[1] [20], \c2[1] [19], \c2[1] [18], \c2[1] [17], 
      \c2[1] [16], \c2[1] [15], \c2[1] [14], \c2[1] [13], \c2[1] [12], 
      \c2[1] [11], \c2[1] [10], \c2[1] [9], uc_1409, uc_1410, uc_1411, uc_1412, 
      uc_1413, uc_1414, uc_1415, uc_1416, uc_1417}), .in2({\s2[2] [45], uc_1418, 
      uc_1419, uc_1420, uc_1421, uc_1422, uc_1423, uc_1424, uc_1425, uc_1426, 
      uc_1427, uc_1428, uc_1429, uc_1430, uc_1431, uc_1432, uc_1433, uc_1434, 
      uc_1435, \s2[2] [44], \s2[2] [43], \s2[2] [42], \s2[2] [41], \s2[2] [40], 
      \s2[2] [39], \s2[2] [38], \s2[2] [37], \s2[2] [36], \s2[2] [35], 
      \s2[2] [34], \s2[2] [33], \s2[2] [32], \s2[2] [31], \s2[2] [30], 
      \s2[2] [29], \s2[2] [28], \s2[2] [27], \s2[2] [26], \s2[2] [25], 
      \s2[2] [24], \s2[2] [23], \s2[2] [22], \s2[2] [21], \s2[2] [20], 
      \s2[2] [19], \s2[2] [18], \s2[2] [17], \s2[2] [16], \s2[2] [15], 
      \s2[2] [14], \s2[2] [13], \s2[2] [12], \s2[2] [11], \s1[3] [10], n_0_288, 
      uc_1436, uc_1437, uc_1438, uc_1439, uc_1440, uc_1441, uc_1442, uc_1443, 
      uc_1444}), .in3({\c2[2] [46], uc_1445, uc_1446, uc_1447, uc_1448, uc_1449, 
      uc_1450, uc_1451, uc_1452, uc_1453, uc_1454, uc_1455, uc_1456, uc_1457, 
      uc_1458, uc_1459, uc_1460, uc_1461, \c2[2] [45], \c2[2] [44], \c2[2] [43], 
      \c2[2] [42], \c2[2] [41], \c2[2] [40], \c2[2] [39], \c2[2] [38], 
      \c2[2] [37], \c2[2] [36], \c2[2] [35], \c2[2] [34], \c2[2] [33], 
      \c2[2] [32], \c2[2] [31], \c2[2] [30], \c2[2] [29], \c2[2] [28], 
      \c2[2] [27], \c2[2] [26], \c2[2] [25], \c2[2] [24], \c2[2] [23], 
      \c2[2] [22], \c2[2] [21], \c2[2] [20], \c2[2] [19], \c2[2] [18], 
      \c2[2] [17], \c2[2] [16], \c2[2] [15], \c2[2] [14], \c2[2] [13], 
      \c2[2] [12], uc_1462, uc_1463, uc_1464, uc_1465, uc_1466, uc_1467, uc_1468, 
      uc_1469, uc_1470, uc_1471, uc_1472, uc_1473}), .sum({\s3[1] [46], uc_1474, 
      uc_1475, uc_1476, uc_1477, uc_1478, uc_1479, uc_1480, uc_1481, uc_1482, 
      uc_1483, uc_1484, uc_1485, uc_1486, uc_1487, uc_1488, uc_1489, uc_1490, 
      \s3[1] [45], \s3[1] [44], \s3[1] [43], \s3[1] [42], \s3[1] [41], 
      \s3[1] [40], \s3[1] [39], \s3[1] [38], \s3[1] [37], \s3[1] [36], 
      \s3[1] [35], \s3[1] [34], \s3[1] [33], \s3[1] [32], \s3[1] [31], 
      \s3[1] [30], \s3[1] [29], \s3[1] [28], \s3[1] [27], \s3[1] [26], 
      \s3[1] [25], \s3[1] [24], \s3[1] [23], \s3[1] [22], \s3[1] [21], 
      \s3[1] [20], \s3[1] [19], \s3[1] [18], \s3[1] [17], \s3[1] [16], 
      \s3[1] [15], \s3[1] [14], \s3[1] [13], \s3[1] [12], \s3[1] [11], 
      \s3[1] [10], \s3[1] [9], uc_1491, uc_1492, uc_1493, uc_1494, uc_1495, 
      uc_1496, uc_1497, uc_1498, uc_1499}), .c({\c3[1] [47], uc_1500, uc_1501, 
      uc_1502, uc_1503, uc_1504, uc_1505, uc_1506, uc_1507, uc_1508, uc_1509, 
      uc_1510, uc_1511, uc_1512, uc_1513, uc_1514, uc_1515, \c3[1] [46], 
      \c3[1] [45], \c3[1] [44], \c3[1] [43], \c3[1] [42], \c3[1] [41], 
      \c3[1] [40], \c3[1] [39], \c3[1] [38], \c3[1] [37], \c3[1] [36], 
      \c3[1] [35], \c3[1] [34], \c3[1] [33], \c3[1] [32], \c3[1] [31], 
      \c3[1] [30], \c3[1] [29], \c3[1] [28], \c3[1] [27], \c3[1] [26], 
      \c3[1] [25], \c3[1] [24], \c3[1] [23], \c3[1] [22], \c3[1] [21], 
      \c3[1] [20], \c3[1] [19], \c3[1] [18], \c3[1] [17], \c3[1] [16], 
      \c3[1] [15], \c3[1] [14], \c3[1] [13], \c3[1] [12], \c3[1] [11], 
      \c3[1] [10], uc_1516, uc_1517, uc_1518, uc_1519, uc_1520, uc_1521, uc_1522, 
      uc_1523, uc_1524, uc_1525}));
   CSA__1_32 A4_1 (.in1({\s3[0] [40], uc_1526, uc_1527, uc_1528, uc_1529, 
      uc_1530, uc_1531, uc_1532, uc_1533, uc_1534, uc_1535, uc_1536, uc_1537, 
      uc_1538, uc_1539, uc_1540, uc_1541, uc_1542, uc_1543, uc_1544, uc_1545, 
      uc_1546, uc_1547, uc_1548, \s3[0] [39], \s3[0] [38], \s3[0] [37], 
      \s3[0] [36], \s3[0] [35], \s3[0] [34], \s3[0] [33], \s3[0] [32], 
      \s3[0] [31], \s3[0] [30], \s3[0] [29], \s3[0] [28], \s3[0] [27], 
      \s3[0] [26], \s3[0] [25], \s3[0] [24], \s3[0] [23], \s3[0] [22], 
      \s3[0] [21], \s3[0] [20], \s3[0] [19], \s3[0] [18], \s3[0] [17], 
      \s3[0] [16], \s3[0] [15], \s3[0] [14], \s3[0] [13], \s3[0] [12], 
      \s3[0] [11], \s3[0] [10], \s3[0] [9], \s3[0] [8], \s3[0] [7], \s3[0] [6], 
      \s3[0] [5], \s3[0] [4], uc_1549, uc_1550, uc_1551, uc_1552}), .in2({
      \c3[0] [41], uc_1553, uc_1554, uc_1555, uc_1556, uc_1557, uc_1558, uc_1559, 
      uc_1560, uc_1561, uc_1562, uc_1563, uc_1564, uc_1565, uc_1566, uc_1567, 
      uc_1568, uc_1569, uc_1570, uc_1571, uc_1572, uc_1573, uc_1574, \c3[0] [40], 
      \c3[0] [39], \c3[0] [38], \c3[0] [37], \c3[0] [36], \c3[0] [35], 
      \c3[0] [34], \c3[0] [33], \c3[0] [32], \c3[0] [31], \c3[0] [30], 
      \c3[0] [29], \c3[0] [28], \c3[0] [27], \c3[0] [26], \c3[0] [25], 
      \c3[0] [24], \c3[0] [23], \c3[0] [22], \c3[0] [21], \c3[0] [20], 
      \c3[0] [19], \c3[0] [18], \c3[0] [17], \c3[0] [16], \c3[0] [15], 
      \c3[0] [14], \c3[0] [13], \c3[0] [12], \c3[0] [11], \c3[0] [10], 
      \c3[0] [9], \c3[0] [8], \c3[0] [7], \c3[0] [6], \c3[0] [5], \c3[0] [4], 
      uc_1575, uc_1576, uc_1577, uc_1578}), .in3({\s3[1] [46], uc_1579, uc_1580, 
      uc_1581, uc_1582, uc_1583, uc_1584, uc_1585, uc_1586, uc_1587, uc_1588, 
      uc_1589, uc_1590, uc_1591, uc_1592, uc_1593, uc_1594, uc_1595, \s3[1] [45], 
      \s3[1] [44], \s3[1] [43], \s3[1] [42], \s3[1] [41], \s3[1] [40], 
      \s3[1] [39], \s3[1] [38], \s3[1] [37], \s3[1] [36], \s3[1] [35], 
      \s3[1] [34], \s3[1] [33], \s3[1] [32], \s3[1] [31], \s3[1] [30], 
      \s3[1] [29], \s3[1] [28], \s3[1] [27], \s3[1] [26], \s3[1] [25], 
      \s3[1] [24], \s3[1] [23], \s3[1] [22], \s3[1] [21], \s3[1] [20], 
      \s3[1] [19], \s3[1] [18], \s3[1] [17], \s3[1] [16], \s3[1] [15], 
      \s3[1] [14], \s3[1] [13], \s3[1] [12], \s3[1] [11], \s3[1] [10], 
      \s3[1] [9], \c2[1] [8], \c2[1] [7], uc_1596, uc_1597, uc_1598, uc_1599, 
      uc_1600, uc_1601, uc_1602}), .sum({\s4[0] [46], uc_1603, uc_1604, uc_1605, 
      uc_1606, uc_1607, uc_1608, uc_1609, uc_1610, uc_1611, uc_1612, uc_1613, 
      uc_1614, uc_1615, uc_1616, uc_1617, uc_1618, uc_1619, \s4[0] [45], 
      \s4[0] [44], \s4[0] [43], \s4[0] [42], \s4[0] [41], \s4[0] [40], 
      \s4[0] [39], \s4[0] [38], \s4[0] [37], \s4[0] [36], \s4[0] [35], 
      \s4[0] [34], \s4[0] [33], \s4[0] [32], \s4[0] [31], \s4[0] [30], 
      \s4[0] [29], \s4[0] [28], \s4[0] [27], \s4[0] [26], \s4[0] [25], 
      \s4[0] [24], \s4[0] [23], \s4[0] [22], \s4[0] [21], \s4[0] [20], 
      \s4[0] [19], \s4[0] [18], \s4[0] [17], \s4[0] [16], \s4[0] [15], 
      \s4[0] [14], \s4[0] [13], \s4[0] [12], \s4[0] [11], \s4[0] [10], 
      \s4[0] [9], \s4[0] [8], \s4[0] [7], \s4[0] [6], \s4[0] [5], c[4], uc_1620, 
      uc_1621, uc_1622, uc_1623}), .c({\c4[0] [47], uc_1624, uc_1625, uc_1626, 
      uc_1627, uc_1628, uc_1629, uc_1630, uc_1631, uc_1632, uc_1633, uc_1634, 
      uc_1635, uc_1636, uc_1637, uc_1638, uc_1639, \c4[0] [46], \c4[0] [45], 
      \c4[0] [44], \c4[0] [43], \c4[0] [42], \c4[0] [41], \c4[0] [40], 
      \c4[0] [39], \c4[0] [38], \c4[0] [37], \c4[0] [36], \c4[0] [35], 
      \c4[0] [34], \c4[0] [33], \c4[0] [32], \c4[0] [31], \c4[0] [30], 
      \c4[0] [29], \c4[0] [28], \c4[0] [27], \c4[0] [26], \c4[0] [25], 
      \c4[0] [24], \c4[0] [23], \c4[0] [22], \c4[0] [21], \c4[0] [20], 
      \c4[0] [19], \c4[0] [18], \c4[0] [17], \c4[0] [16], \c4[0] [15], 
      \c4[0] [14], \c4[0] [13], \c4[0] [12], \c4[0] [11], \c4[0] [10], 
      \c4[0] [9], \c4[0] [8], \c4[0] [7], \c4[0] [6], \c4[0] [5], uc_1640, 
      uc_1641, uc_1642, uc_1643, uc_1644}));
   CSA__1_35 A2_6 (.in1({\c1[7] [55], uc_1645, uc_1646, uc_1647, uc_1648, 
      uc_1649, uc_1650, uc_1651, uc_1652, \c1[7] [54], \c1[7] [53], \c1[7] [52], 
      \c1[7] [51], \c1[7] [50], \c1[7] [49], \c1[7] [48], \c1[7] [47], 
      \c1[7] [46], \c1[7] [45], \c1[7] [44], \c1[7] [43], \c1[7] [42], 
      \c1[7] [41], \c1[7] [40], \c1[7] [39], \c1[7] [38], \c1[7] [37], 
      \c1[7] [36], \c1[7] [35], \c1[7] [34], \c1[7] [33], \c1[7] [32], 
      \c1[7] [31], \c1[7] [30], \c1[7] [29], \c1[7] [28], \c1[7] [27], 
      \c1[7] [26], \c1[7] [25], \c1[7] [24], uc_1653, uc_1654, uc_1655, uc_1656, 
      uc_1657, uc_1658, uc_1659, uc_1660, uc_1661, uc_1662, uc_1663, uc_1664, 
      uc_1665, uc_1666, uc_1667, uc_1668, uc_1669, uc_1670, uc_1671, uc_1672, 
      uc_1673, uc_1674, uc_1675, uc_1676}), .in2({\s1[8] [57], uc_1677, uc_1678, 
      uc_1679, uc_1680, uc_1681, uc_1682, \s1[8] [56], \s1[8] [55], \s1[8] [54], 
      \s1[8] [53], \s1[8] [52], \s1[8] [51], \s1[8] [50], \s1[8] [49], 
      \s1[8] [48], \s1[8] [47], \s1[8] [46], \s1[8] [45], \s1[8] [44], 
      \s1[8] [43], \s1[8] [42], \s1[8] [41], \s1[8] [40], \s1[8] [39], 
      \s1[8] [38], \s1[8] [37], \s1[8] [36], \s1[8] [35], \s1[8] [34], 
      \s1[8] [33], \s1[8] [32], \s1[8] [31], \s1[8] [30], \s1[8] [29], 
      \s1[8] [28], \s1[8] [27], \s1[8] [26], \s1[8] [25], n_0_96, uc_1683, 
      uc_1684, uc_1685, uc_1686, uc_1687, uc_1688, uc_1689, uc_1690, uc_1691, 
      uc_1692, uc_1693, uc_1694, uc_1695, uc_1696, uc_1697, uc_1698, uc_1699, 
      uc_1700, uc_1701, uc_1702, uc_1703, uc_1704, uc_1705, uc_1706}), .in3({
      \c1[8] [58], uc_1707, uc_1708, uc_1709, uc_1710, uc_1711, \c1[8] [57], 
      \c1[8] [56], \c1[8] [55], \c1[8] [54], \c1[8] [53], \c1[8] [52], 
      \c1[8] [51], \c1[8] [50], \c1[8] [49], \c1[8] [48], \c1[8] [47], 
      \c1[8] [46], \c1[8] [45], \c1[8] [44], \c1[8] [43], \c1[8] [42], 
      \c1[8] [41], \c1[8] [40], \c1[8] [39], \c1[8] [38], \c1[8] [37], 
      \c1[8] [36], \c1[8] [35], \c1[8] [34], \c1[8] [33], \c1[8] [32], 
      \c1[8] [31], \c1[8] [30], \c1[8] [29], \c1[8] [28], \c1[8] [27], 
      \c1[8] [26], uc_1712, uc_1713, uc_1714, uc_1715, uc_1716, uc_1717, uc_1718, 
      uc_1719, uc_1720, uc_1721, uc_1722, uc_1723, uc_1724, uc_1725, uc_1726, 
      uc_1727, uc_1728, uc_1729, uc_1730, uc_1731, uc_1732, uc_1733, uc_1734, 
      uc_1735, uc_1736, uc_1737}), .sum({\s2[5] [58], uc_1738, uc_1739, uc_1740, 
      uc_1741, uc_1742, \s2[5] [57], \s2[5] [56], \s2[5] [55], \s2[5] [54], 
      \s2[5] [53], \s2[5] [52], \s2[5] [51], \s2[5] [50], \s2[5] [49], 
      \s2[5] [48], \s2[5] [47], \s2[5] [46], \s2[5] [45], \s2[5] [44], 
      \s2[5] [43], \s2[5] [42], \s2[5] [41], \s2[5] [40], \s2[5] [39], 
      \s2[5] [38], \s2[5] [37], \s2[5] [36], \s2[5] [35], \s2[5] [34], 
      \s2[5] [33], \s2[5] [32], \s2[5] [31], \s2[5] [30], \s2[5] [29], 
      \s2[5] [28], \s2[5] [27], \s2[5] [26], \s2[5] [25], \s2[5] [24], uc_1743, 
      uc_1744, uc_1745, uc_1746, uc_1747, uc_1748, uc_1749, uc_1750, uc_1751, 
      uc_1752, uc_1753, uc_1754, uc_1755, uc_1756, uc_1757, uc_1758, uc_1759, 
      uc_1760, uc_1761, uc_1762, uc_1763, uc_1764, uc_1765, uc_1766}), .c({
      \c2[5] [59], uc_1767, uc_1768, uc_1769, uc_1770, \c2[5] [58], \c2[5] [57], 
      \c2[5] [56], \c2[5] [55], \c2[5] [54], \c2[5] [53], \c2[5] [52], 
      \c2[5] [51], \c2[5] [50], \c2[5] [49], \c2[5] [48], \c2[5] [47], 
      \c2[5] [46], \c2[5] [45], \c2[5] [44], \c2[5] [43], \c2[5] [42], 
      \c2[5] [41], \c2[5] [40], \c2[5] [39], \c2[5] [38], \c2[5] [37], 
      \c2[5] [36], \c2[5] [35], \c2[5] [34], \c2[5] [33], \c2[5] [32], 
      \c2[5] [31], \c2[5] [30], \c2[5] [29], \c2[5] [28], \c2[5] [27], 
      \c2[5] [26], \c2[5] [25], uc_1771, uc_1772, uc_1773, uc_1774, uc_1775, 
      uc_1776, uc_1777, uc_1778, uc_1779, uc_1780, uc_1781, uc_1782, uc_1783, 
      uc_1784, uc_1785, uc_1786, uc_1787, uc_1788, uc_1789, uc_1790, uc_1791, 
      uc_1792, uc_1793, uc_1794, uc_1795}));
   CSA__1_38 A3_4 (.in1({\c2[4] [55], uc_1796, uc_1797, uc_1798, uc_1799, 
      uc_1800, uc_1801, uc_1802, uc_1803, \c2[4] [54], \c2[4] [53], \c2[4] [52], 
      \c2[4] [51], \c2[4] [50], \c2[4] [49], \c2[4] [48], \c2[4] [47], 
      \c2[4] [46], \c2[4] [45], \c2[4] [44], \c2[4] [43], \c2[4] [42], 
      \c2[4] [41], \c2[4] [40], \c2[4] [39], \c2[4] [38], \c2[4] [37], 
      \c2[4] [36], \c2[4] [35], \c2[4] [34], \c2[4] [33], \c2[4] [32], 
      \c2[4] [31], \c2[4] [30], \c2[4] [29], \c2[4] [28], \c2[4] [27], 
      \c2[4] [26], \c2[4] [25], \c2[4] [24], \c2[4] [23], uc_1804, uc_1805, 
      uc_1806, uc_1807, uc_1808, uc_1809, uc_1810, uc_1811, uc_1812, uc_1813, 
      uc_1814, uc_1815, uc_1816, uc_1817, uc_1818, uc_1819, uc_1820, uc_1821, 
      uc_1822, uc_1823, uc_1824, uc_1825, uc_1826}), .in2({\s2[5] [58], uc_1827, 
      uc_1828, uc_1829, uc_1830, uc_1831, \s2[5] [57], \s2[5] [56], \s2[5] [55], 
      \s2[5] [54], \s2[5] [53], \s2[5] [52], \s2[5] [51], \s2[5] [50], 
      \s2[5] [49], \s2[5] [48], \s2[5] [47], \s2[5] [46], \s2[5] [45], 
      \s2[5] [44], \s2[5] [43], \s2[5] [42], \s2[5] [41], \s2[5] [40], 
      \s2[5] [39], \s2[5] [38], \s2[5] [37], \s2[5] [36], \s2[5] [35], 
      \s2[5] [34], \s2[5] [33], \s2[5] [32], \s2[5] [31], \s2[5] [30], 
      \s2[5] [29], \s2[5] [28], \s2[5] [27], \s2[5] [26], \s2[5] [25], 
      \s2[5] [24], \c1[7] [23], uc_1832, uc_1833, uc_1834, uc_1835, uc_1836, 
      uc_1837, uc_1838, uc_1839, uc_1840, uc_1841, uc_1842, uc_1843, uc_1844, 
      uc_1845, uc_1846, uc_1847, uc_1848, uc_1849, uc_1850, uc_1851, uc_1852, 
      uc_1853, uc_1854}), .in3({\c2[5] [59], uc_1855, uc_1856, uc_1857, uc_1858, 
      \c2[5] [58], \c2[5] [57], \c2[5] [56], \c2[5] [55], \c2[5] [54], 
      \c2[5] [53], \c2[5] [52], \c2[5] [51], \c2[5] [50], \c2[5] [49], 
      \c2[5] [48], \c2[5] [47], \c2[5] [46], \c2[5] [45], \c2[5] [44], 
      \c2[5] [43], \c2[5] [42], \c2[5] [41], \c2[5] [40], \c2[5] [39], 
      \c2[5] [38], \c2[5] [37], \c2[5] [36], \c2[5] [35], \c2[5] [34], 
      \c2[5] [33], \c2[5] [32], \c2[5] [31], \c2[5] [30], \c2[5] [29], 
      \c2[5] [28], \c2[5] [27], \c2[5] [26], \c2[5] [25], uc_1859, uc_1860, 
      uc_1861, uc_1862, uc_1863, uc_1864, uc_1865, uc_1866, uc_1867, uc_1868, 
      uc_1869, uc_1870, uc_1871, uc_1872, uc_1873, uc_1874, uc_1875, uc_1876, 
      uc_1877, uc_1878, uc_1879, uc_1880, uc_1881, uc_1882, uc_1883}), .sum({
      \s3[3] [59], uc_1884, uc_1885, uc_1886, uc_1887, \s3[3] [58], \s3[3] [57], 
      \s3[3] [56], \s3[3] [55], \s3[3] [54], \s3[3] [53], \s3[3] [52], 
      \s3[3] [51], \s3[3] [50], \s3[3] [49], \s3[3] [48], \s3[3] [47], 
      \s3[3] [46], \s3[3] [45], \s3[3] [44], \s3[3] [43], \s3[3] [42], 
      \s3[3] [41], \s3[3] [40], \s3[3] [39], \s3[3] [38], \s3[3] [37], 
      \s3[3] [36], \s3[3] [35], \s3[3] [34], \s3[3] [33], \s3[3] [32], 
      \s3[3] [31], \s3[3] [30], \s3[3] [29], \s3[3] [28], \s3[3] [27], 
      \s3[3] [26], \s3[3] [25], \s3[3] [24], \s3[3] [23], uc_1888, uc_1889, 
      uc_1890, uc_1891, uc_1892, uc_1893, uc_1894, uc_1895, uc_1896, uc_1897, 
      uc_1898, uc_1899, uc_1900, uc_1901, uc_1902, uc_1903, uc_1904, uc_1905, 
      uc_1906, uc_1907, uc_1908, uc_1909, uc_1910}), .c({\c3[3] [60], uc_1911, 
      uc_1912, uc_1913, \c3[3] [59], \c3[3] [58], \c3[3] [57], \c3[3] [56], 
      \c3[3] [55], \c3[3] [54], \c3[3] [53], \c3[3] [52], \c3[3] [51], 
      \c3[3] [50], \c3[3] [49], \c3[3] [48], \c3[3] [47], \c3[3] [46], 
      \c3[3] [45], \c3[3] [44], \c3[3] [43], \c3[3] [42], \c3[3] [41], 
      \c3[3] [40], \c3[3] [39], \c3[3] [38], \c3[3] [37], \c3[3] [36], 
      \c3[3] [35], \c3[3] [34], \c3[3] [33], \c3[3] [32], \c3[3] [31], 
      \c3[3] [30], \c3[3] [29], \c3[3] [28], \c3[3] [27], \c3[3] [26], 
      \c3[3] [25], \c3[3] [24], uc_1914, uc_1915, uc_1916, uc_1917, uc_1918, 
      uc_1919, uc_1920, uc_1921, uc_1922, uc_1923, uc_1924, uc_1925, uc_1926, 
      uc_1927, uc_1928, uc_1929, uc_1930, uc_1931, uc_1932, uc_1933, uc_1934, 
      uc_1935, uc_1936, uc_1937}));
   CSA__0_68 A1_8 (.in1({n_0_223, uc_1938, uc_1939, uc_1940, uc_1941, uc_1942, 
      uc_1943, uc_1944, uc_1945, uc_1946, uc_1947, uc_1948, n_0_222, n_0_221, 
      n_0_220, n_0_219, n_0_218, n_0_217, n_0_216, n_0_215, n_0_214, n_0_213, 
      n_0_212, n_0_211, n_0_210, n_0_209, n_0_208, n_0_207, n_0_206, n_0_205, 
      n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, n_0_199, n_0_198, n_0_197, 
      n_0_196, n_0_195, n_0_194, n_0_193, uc_1949, uc_1950, uc_1951, uc_1952, 
      uc_1953, uc_1954, uc_1955, uc_1956, uc_1957, uc_1958, uc_1959, uc_1960, 
      uc_1961, uc_1962, uc_1963, uc_1964, uc_1965, uc_1966, uc_1967, uc_1968, 
      uc_1969, uc_1970}), .in2({n_0_191, uc_1971, uc_1972, uc_1973, uc_1974, 
      uc_1975, uc_1976, uc_1977, uc_1978, uc_1979, uc_1980, n_0_190, n_0_189, 
      n_0_188, n_0_187, n_0_186, n_0_185, n_0_184, n_0_183, n_0_182, n_0_181, 
      n_0_180, n_0_179, n_0_178, n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, 
      n_0_172, n_0_171, n_0_170, n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, 
      n_0_164, n_0_163, n_0_162, n_0_161, n_0_160, uc_1981, uc_1982, uc_1983, 
      uc_1984, uc_1985, uc_1986, uc_1987, uc_1988, uc_1989, uc_1990, uc_1991, 
      uc_1992, uc_1993, uc_1994, uc_1995, uc_1996, uc_1997, uc_1998, uc_1999, 
      uc_2000, uc_2001, uc_2002}), .in3({n_0_159, uc_2003, uc_2004, uc_2005, 
      uc_2006, uc_2007, uc_2008, uc_2009, uc_2010, uc_2011, n_0_158, n_0_157, 
      n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, n_0_149, 
      n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, n_0_141, 
      n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, n_0_133, 
      n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, uc_2012, uc_2013, uc_2014, 
      uc_2015, uc_2016, uc_2017, uc_2018, uc_2019, uc_2020, uc_2021, uc_2022, 
      uc_2023, uc_2024, uc_2025, uc_2026, uc_2027, uc_2028, uc_2029, uc_2030, 
      uc_2031, uc_2032, uc_2033, uc_2034}), .sum({\s1[7] [54], uc_2035, uc_2036, 
      uc_2037, uc_2038, uc_2039, uc_2040, uc_2041, uc_2042, uc_2043, \s1[7] [53], 
      \s1[7] [52], \s1[7] [51], \s1[7] [50], \s1[7] [49], \s1[7] [48], 
      \s1[7] [47], \s1[7] [46], \s1[7] [45], \s1[7] [44], \s1[7] [43], 
      \s1[7] [42], \s1[7] [41], \s1[7] [40], \s1[7] [39], \s1[7] [38], 
      \s1[7] [37], \s1[7] [36], \s1[7] [35], \s1[7] [34], \s1[7] [33], 
      \s1[7] [32], \s1[7] [31], \s1[7] [30], \s1[7] [29], \s1[7] [28], 
      \s1[7] [27], \s1[7] [26], \s1[7] [25], \s1[7] [24], \s1[7] [23], 
      \s1[7] [22], uc_2044, uc_2045, uc_2046, uc_2047, uc_2048, uc_2049, uc_2050, 
      uc_2051, uc_2052, uc_2053, uc_2054, uc_2055, uc_2056, uc_2057, uc_2058, 
      uc_2059, uc_2060, uc_2061, uc_2062, uc_2063, uc_2064, uc_2065}), .c({
      \c1[7] [55], uc_2066, uc_2067, uc_2068, uc_2069, uc_2070, uc_2071, uc_2072, 
      uc_2073, \c1[7] [54], \c1[7] [53], \c1[7] [52], \c1[7] [51], \c1[7] [50], 
      \c1[7] [49], \c1[7] [48], \c1[7] [47], \c1[7] [46], \c1[7] [45], 
      \c1[7] [44], \c1[7] [43], \c1[7] [42], \c1[7] [41], \c1[7] [40], 
      \c1[7] [39], \c1[7] [38], \c1[7] [37], \c1[7] [36], \c1[7] [35], 
      \c1[7] [34], \c1[7] [33], \c1[7] [32], \c1[7] [31], \c1[7] [30], 
      \c1[7] [29], \c1[7] [28], \c1[7] [27], \c1[7] [26], \c1[7] [25], 
      \c1[7] [24], \c1[7] [23], uc_2074, uc_2075, uc_2076, uc_2077, uc_2078, 
      uc_2079, uc_2080, uc_2081, uc_2082, uc_2083, uc_2084, uc_2085, uc_2086, 
      uc_2087, uc_2088, uc_2089, uc_2090, uc_2091, uc_2092, uc_2093, uc_2094, 
      uc_2095, uc_2096}));
   INV_X1 i_0_0_1 (.A(a[0]), .ZN(n_0_0_1));
   NOR2_X1 i_0_0_2 (.A1(n_0_0_0), .A2(n_0_0_1), .ZN(c[0]));
   INV_X1 i_0_0_3 (.A(a[1]), .ZN(n_0_0_2));
   NOR2_X1 i_0_0_4 (.A1(n_0_0_0), .A2(n_0_0_2), .ZN(n_0_0));
   INV_X1 i_0_0_5 (.A(a[2]), .ZN(n_0_0_3));
   NOR2_X1 i_0_0_6 (.A1(n_0_0_0), .A2(n_0_0_3), .ZN(n_0_1));
   INV_X1 i_0_0_7 (.A(a[3]), .ZN(n_0_0_4));
   NOR2_X1 i_0_0_8 (.A1(n_0_0_0), .A2(n_0_0_4), .ZN(n_0_2));
   INV_X1 i_0_0_9 (.A(a[4]), .ZN(n_0_0_5));
   NOR2_X1 i_0_0_10 (.A1(n_0_0_0), .A2(n_0_0_5), .ZN(n_0_3));
   INV_X1 i_0_0_11 (.A(a[5]), .ZN(n_0_0_6));
   NOR2_X1 i_0_0_12 (.A1(n_0_0_0), .A2(n_0_0_6), .ZN(n_0_4));
   INV_X1 i_0_0_13 (.A(a[6]), .ZN(n_0_0_7));
   NOR2_X1 i_0_0_14 (.A1(n_0_0_0), .A2(n_0_0_7), .ZN(n_0_5));
   INV_X1 i_0_0_15 (.A(a[7]), .ZN(n_0_0_8));
   NOR2_X1 i_0_0_16 (.A1(n_0_0_0), .A2(n_0_0_8), .ZN(n_0_6));
   INV_X1 i_0_0_17 (.A(a[8]), .ZN(n_0_0_9));
   NOR2_X1 i_0_0_18 (.A1(n_0_0_0), .A2(n_0_0_9), .ZN(n_0_7));
   INV_X1 i_0_0_19 (.A(a[9]), .ZN(n_0_0_10));
   NOR2_X1 i_0_0_20 (.A1(n_0_0_0), .A2(n_0_0_10), .ZN(n_0_8));
   INV_X1 i_0_0_21 (.A(a[10]), .ZN(n_0_0_11));
   NOR2_X1 i_0_0_22 (.A1(n_0_0_0), .A2(n_0_0_11), .ZN(n_0_9));
   INV_X1 i_0_0_23 (.A(a[11]), .ZN(n_0_0_12));
   NOR2_X1 i_0_0_24 (.A1(n_0_0_0), .A2(n_0_0_12), .ZN(n_0_10));
   INV_X1 i_0_0_25 (.A(a[12]), .ZN(n_0_0_13));
   NOR2_X1 i_0_0_26 (.A1(n_0_0_0), .A2(n_0_0_13), .ZN(n_0_11));
   INV_X1 i_0_0_27 (.A(a[13]), .ZN(n_0_0_14));
   NOR2_X1 i_0_0_28 (.A1(n_0_0_0), .A2(n_0_0_14), .ZN(n_0_12));
   INV_X1 i_0_0_29 (.A(a[14]), .ZN(n_0_0_15));
   NOR2_X1 i_0_0_30 (.A1(n_0_0_0), .A2(n_0_0_15), .ZN(n_0_13));
   INV_X1 i_0_0_31 (.A(a[15]), .ZN(n_0_0_16));
   NOR2_X1 i_0_0_32 (.A1(n_0_0_0), .A2(n_0_0_16), .ZN(n_0_14));
   INV_X1 i_0_0_33 (.A(a[16]), .ZN(n_0_0_17));
   NOR2_X1 i_0_0_34 (.A1(n_0_0_0), .A2(n_0_0_17), .ZN(n_0_15));
   INV_X1 i_0_0_35 (.A(a[17]), .ZN(n_0_0_18));
   NOR2_X1 i_0_0_36 (.A1(n_0_0_0), .A2(n_0_0_18), .ZN(n_0_16));
   INV_X1 i_0_0_37 (.A(a[18]), .ZN(n_0_0_19));
   NOR2_X1 i_0_0_38 (.A1(n_0_0_0), .A2(n_0_0_19), .ZN(n_0_17));
   INV_X1 i_0_0_39 (.A(a[19]), .ZN(n_0_0_20));
   NOR2_X1 i_0_0_40 (.A1(n_0_0_0), .A2(n_0_0_20), .ZN(n_0_18));
   INV_X1 i_0_0_41 (.A(a[20]), .ZN(n_0_0_21));
   NOR2_X1 i_0_0_42 (.A1(n_0_0_0), .A2(n_0_0_21), .ZN(n_0_19));
   INV_X1 i_0_0_43 (.A(a[21]), .ZN(n_0_0_22));
   NOR2_X1 i_0_0_44 (.A1(n_0_0_0), .A2(n_0_0_22), .ZN(n_0_20));
   INV_X1 i_0_0_45 (.A(a[22]), .ZN(n_0_0_23));
   NOR2_X1 i_0_0_46 (.A1(n_0_0_0), .A2(n_0_0_23), .ZN(n_0_21));
   INV_X1 i_0_0_47 (.A(a[23]), .ZN(n_0_0_24));
   NOR2_X1 i_0_0_48 (.A1(n_0_0_0), .A2(n_0_0_24), .ZN(n_0_22));
   INV_X1 i_0_0_49 (.A(a[24]), .ZN(n_0_0_25));
   NOR2_X1 i_0_0_50 (.A1(n_0_0_0), .A2(n_0_0_25), .ZN(n_0_23));
   INV_X1 i_0_0_51 (.A(a[25]), .ZN(n_0_0_26));
   NOR2_X1 i_0_0_52 (.A1(n_0_0_0), .A2(n_0_0_26), .ZN(n_0_24));
   INV_X1 i_0_0_53 (.A(a[26]), .ZN(n_0_0_27));
   NOR2_X1 i_0_0_54 (.A1(n_0_0_0), .A2(n_0_0_27), .ZN(n_0_25));
   INV_X1 i_0_0_55 (.A(a[27]), .ZN(n_0_0_28));
   NOR2_X1 i_0_0_56 (.A1(n_0_0_0), .A2(n_0_0_28), .ZN(n_0_26));
   INV_X1 i_0_0_57 (.A(a[28]), .ZN(n_0_0_29));
   NOR2_X1 i_0_0_58 (.A1(n_0_0_0), .A2(n_0_0_29), .ZN(n_0_27));
   INV_X1 i_0_0_59 (.A(a[29]), .ZN(n_0_0_30));
   NOR2_X1 i_0_0_60 (.A1(n_0_0_0), .A2(n_0_0_30), .ZN(n_0_28));
   INV_X1 i_0_0_61 (.A(a[30]), .ZN(n_0_0_31));
   NOR2_X1 i_0_0_62 (.A1(n_0_0_0), .A2(n_0_0_31), .ZN(n_0_29));
   NOR2_X1 i_0_0_66 (.A1(n_0_0_33), .A2(n_0_0_1), .ZN(n_0_544));
   NOR2_X1 i_0_0_67 (.A1(n_0_0_33), .A2(n_0_0_2), .ZN(n_0_545));
   NOR2_X1 i_0_0_68 (.A1(n_0_0_33), .A2(n_0_0_3), .ZN(n_0_546));
   NOR2_X1 i_0_0_69 (.A1(n_0_0_33), .A2(n_0_0_4), .ZN(n_0_547));
   NOR2_X1 i_0_0_70 (.A1(n_0_0_33), .A2(n_0_0_5), .ZN(n_0_548));
   NOR2_X1 i_0_0_71 (.A1(n_0_0_33), .A2(n_0_0_6), .ZN(n_0_549));
   NOR2_X1 i_0_0_72 (.A1(n_0_0_33), .A2(n_0_0_7), .ZN(n_0_550));
   NOR2_X1 i_0_0_73 (.A1(n_0_0_33), .A2(n_0_0_8), .ZN(n_0_551));
   NOR2_X1 i_0_0_74 (.A1(n_0_0_33), .A2(n_0_0_9), .ZN(n_0_552));
   NOR2_X1 i_0_0_75 (.A1(n_0_0_33), .A2(n_0_0_10), .ZN(n_0_553));
   NOR2_X1 i_0_0_76 (.A1(n_0_0_33), .A2(n_0_0_11), .ZN(n_0_554));
   NOR2_X1 i_0_0_77 (.A1(n_0_0_33), .A2(n_0_0_12), .ZN(n_0_555));
   NOR2_X1 i_0_0_78 (.A1(n_0_0_33), .A2(n_0_0_13), .ZN(n_0_556));
   NOR2_X1 i_0_0_79 (.A1(n_0_0_33), .A2(n_0_0_14), .ZN(n_0_557));
   NOR2_X1 i_0_0_80 (.A1(n_0_0_33), .A2(n_0_0_15), .ZN(n_0_558));
   NOR2_X1 i_0_0_81 (.A1(n_0_0_33), .A2(n_0_0_16), .ZN(n_0_559));
   NOR2_X1 i_0_0_82 (.A1(n_0_0_33), .A2(n_0_0_17), .ZN(n_0_560));
   NOR2_X1 i_0_0_83 (.A1(n_0_0_33), .A2(n_0_0_18), .ZN(n_0_561));
   NOR2_X1 i_0_0_84 (.A1(n_0_0_33), .A2(n_0_0_19), .ZN(n_0_562));
   NOR2_X1 i_0_0_85 (.A1(n_0_0_33), .A2(n_0_0_20), .ZN(n_0_563));
   NOR2_X1 i_0_0_86 (.A1(n_0_0_33), .A2(n_0_0_21), .ZN(n_0_564));
   NOR2_X1 i_0_0_87 (.A1(n_0_0_33), .A2(n_0_0_22), .ZN(n_0_565));
   NOR2_X1 i_0_0_88 (.A1(n_0_0_33), .A2(n_0_0_23), .ZN(n_0_566));
   NOR2_X1 i_0_0_89 (.A1(n_0_0_33), .A2(n_0_0_24), .ZN(n_0_567));
   NOR2_X1 i_0_0_90 (.A1(n_0_0_33), .A2(n_0_0_25), .ZN(n_0_568));
   NOR2_X1 i_0_0_91 (.A1(n_0_0_33), .A2(n_0_0_26), .ZN(n_0_569));
   NOR2_X1 i_0_0_92 (.A1(n_0_0_33), .A2(n_0_0_27), .ZN(n_0_570));
   NOR2_X1 i_0_0_93 (.A1(n_0_0_33), .A2(n_0_0_28), .ZN(n_0_571));
   NOR2_X1 i_0_0_94 (.A1(n_0_0_33), .A2(n_0_0_29), .ZN(n_0_572));
   NOR2_X1 i_0_0_95 (.A1(n_0_0_33), .A2(n_0_0_30), .ZN(n_0_573));
   NOR2_X1 i_0_0_96 (.A1(n_0_0_33), .A2(n_0_0_31), .ZN(n_0_31));
   INV_X1 i_0_0_98 (.A(b[2]), .ZN(n_0_0_34));
   NOR2_X1 i_0_0_99 (.A1(n_0_0_34), .A2(n_0_0_1), .ZN(n_0_512));
   NOR2_X1 i_0_0_100 (.A1(n_0_0_34), .A2(n_0_0_2), .ZN(n_0_513));
   NOR2_X1 i_0_0_101 (.A1(n_0_0_34), .A2(n_0_0_3), .ZN(n_0_514));
   NOR2_X1 i_0_0_102 (.A1(n_0_0_34), .A2(n_0_0_4), .ZN(n_0_515));
   NOR2_X1 i_0_0_103 (.A1(n_0_0_34), .A2(n_0_0_5), .ZN(n_0_516));
   NOR2_X1 i_0_0_104 (.A1(n_0_0_34), .A2(n_0_0_6), .ZN(n_0_517));
   NOR2_X1 i_0_0_105 (.A1(n_0_0_34), .A2(n_0_0_7), .ZN(n_0_518));
   NOR2_X1 i_0_0_106 (.A1(n_0_0_34), .A2(n_0_0_8), .ZN(n_0_519));
   NOR2_X1 i_0_0_107 (.A1(n_0_0_34), .A2(n_0_0_9), .ZN(n_0_520));
   NOR2_X1 i_0_0_108 (.A1(n_0_0_34), .A2(n_0_0_10), .ZN(n_0_521));
   NOR2_X1 i_0_0_109 (.A1(n_0_0_34), .A2(n_0_0_11), .ZN(n_0_522));
   NOR2_X1 i_0_0_110 (.A1(n_0_0_34), .A2(n_0_0_12), .ZN(n_0_523));
   NOR2_X1 i_0_0_111 (.A1(n_0_0_34), .A2(n_0_0_13), .ZN(n_0_524));
   NOR2_X1 i_0_0_112 (.A1(n_0_0_34), .A2(n_0_0_14), .ZN(n_0_525));
   NOR2_X1 i_0_0_113 (.A1(n_0_0_34), .A2(n_0_0_15), .ZN(n_0_526));
   NOR2_X1 i_0_0_114 (.A1(n_0_0_34), .A2(n_0_0_16), .ZN(n_0_527));
   NOR2_X1 i_0_0_115 (.A1(n_0_0_34), .A2(n_0_0_17), .ZN(n_0_528));
   NOR2_X1 i_0_0_116 (.A1(n_0_0_34), .A2(n_0_0_18), .ZN(n_0_529));
   NOR2_X1 i_0_0_117 (.A1(n_0_0_34), .A2(n_0_0_19), .ZN(n_0_530));
   NOR2_X1 i_0_0_118 (.A1(n_0_0_34), .A2(n_0_0_20), .ZN(n_0_531));
   NOR2_X1 i_0_0_119 (.A1(n_0_0_34), .A2(n_0_0_21), .ZN(n_0_532));
   NOR2_X1 i_0_0_120 (.A1(n_0_0_34), .A2(n_0_0_22), .ZN(n_0_533));
   NOR2_X1 i_0_0_121 (.A1(n_0_0_34), .A2(n_0_0_23), .ZN(n_0_534));
   NOR2_X1 i_0_0_122 (.A1(n_0_0_34), .A2(n_0_0_24), .ZN(n_0_535));
   NOR2_X1 i_0_0_123 (.A1(n_0_0_34), .A2(n_0_0_25), .ZN(n_0_536));
   NOR2_X1 i_0_0_124 (.A1(n_0_0_34), .A2(n_0_0_26), .ZN(n_0_537));
   NOR2_X1 i_0_0_125 (.A1(n_0_0_34), .A2(n_0_0_27), .ZN(n_0_538));
   NOR2_X1 i_0_0_126 (.A1(n_0_0_34), .A2(n_0_0_28), .ZN(n_0_539));
   NOR2_X1 i_0_0_127 (.A1(n_0_0_34), .A2(n_0_0_29), .ZN(n_0_540));
   NOR2_X1 i_0_0_128 (.A1(n_0_0_34), .A2(n_0_0_30), .ZN(n_0_541));
   NOR2_X1 i_0_0_129 (.A1(n_0_0_34), .A2(n_0_0_31), .ZN(n_0_542));
   NOR2_X1 i_0_0_130 (.A1(n_0_0_34), .A2(n_0_0_32), .ZN(n_0_543));
   INV_X1 i_0_0_131 (.A(b[3]), .ZN(n_0_0_35));
   NOR2_X1 i_0_0_132 (.A1(n_0_0_35), .A2(n_0_0_1), .ZN(n_0_480));
   NOR2_X1 i_0_0_133 (.A1(n_0_0_35), .A2(n_0_0_2), .ZN(n_0_481));
   NOR2_X1 i_0_0_134 (.A1(n_0_0_35), .A2(n_0_0_3), .ZN(n_0_482));
   NOR2_X1 i_0_0_135 (.A1(n_0_0_35), .A2(n_0_0_4), .ZN(n_0_483));
   NOR2_X1 i_0_0_136 (.A1(n_0_0_35), .A2(n_0_0_5), .ZN(n_0_484));
   NOR2_X1 i_0_0_137 (.A1(n_0_0_35), .A2(n_0_0_6), .ZN(n_0_485));
   NOR2_X1 i_0_0_138 (.A1(n_0_0_35), .A2(n_0_0_7), .ZN(n_0_486));
   NOR2_X1 i_0_0_139 (.A1(n_0_0_35), .A2(n_0_0_8), .ZN(n_0_487));
   NOR2_X1 i_0_0_140 (.A1(n_0_0_35), .A2(n_0_0_9), .ZN(n_0_488));
   NOR2_X1 i_0_0_141 (.A1(n_0_0_35), .A2(n_0_0_10), .ZN(n_0_489));
   NOR2_X1 i_0_0_142 (.A1(n_0_0_35), .A2(n_0_0_11), .ZN(n_0_490));
   NOR2_X1 i_0_0_143 (.A1(n_0_0_35), .A2(n_0_0_12), .ZN(n_0_491));
   NOR2_X1 i_0_0_144 (.A1(n_0_0_35), .A2(n_0_0_13), .ZN(n_0_492));
   NOR2_X1 i_0_0_145 (.A1(n_0_0_35), .A2(n_0_0_14), .ZN(n_0_493));
   NOR2_X1 i_0_0_146 (.A1(n_0_0_35), .A2(n_0_0_15), .ZN(n_0_494));
   NOR2_X1 i_0_0_147 (.A1(n_0_0_35), .A2(n_0_0_16), .ZN(n_0_495));
   NOR2_X1 i_0_0_148 (.A1(n_0_0_35), .A2(n_0_0_17), .ZN(n_0_496));
   NOR2_X1 i_0_0_149 (.A1(n_0_0_35), .A2(n_0_0_18), .ZN(n_0_497));
   NOR2_X1 i_0_0_150 (.A1(n_0_0_35), .A2(n_0_0_19), .ZN(n_0_498));
   NOR2_X1 i_0_0_151 (.A1(n_0_0_35), .A2(n_0_0_20), .ZN(n_0_499));
   NOR2_X1 i_0_0_152 (.A1(n_0_0_35), .A2(n_0_0_21), .ZN(n_0_500));
   NOR2_X1 i_0_0_153 (.A1(n_0_0_35), .A2(n_0_0_22), .ZN(n_0_501));
   NOR2_X1 i_0_0_154 (.A1(n_0_0_35), .A2(n_0_0_23), .ZN(n_0_502));
   NOR2_X1 i_0_0_155 (.A1(n_0_0_35), .A2(n_0_0_24), .ZN(n_0_503));
   NOR2_X1 i_0_0_156 (.A1(n_0_0_35), .A2(n_0_0_25), .ZN(n_0_504));
   NOR2_X1 i_0_0_157 (.A1(n_0_0_35), .A2(n_0_0_26), .ZN(n_0_505));
   NOR2_X1 i_0_0_158 (.A1(n_0_0_35), .A2(n_0_0_27), .ZN(n_0_506));
   NOR2_X1 i_0_0_159 (.A1(n_0_0_35), .A2(n_0_0_28), .ZN(n_0_507));
   NOR2_X1 i_0_0_160 (.A1(n_0_0_35), .A2(n_0_0_29), .ZN(n_0_508));
   NOR2_X1 i_0_0_161 (.A1(n_0_0_35), .A2(n_0_0_30), .ZN(n_0_509));
   NOR2_X1 i_0_0_162 (.A1(n_0_0_35), .A2(n_0_0_31), .ZN(n_0_510));
   NOR2_X1 i_0_0_163 (.A1(n_0_0_35), .A2(n_0_0_32), .ZN(n_0_511));
   INV_X1 i_0_0_164 (.A(b[4]), .ZN(n_0_0_36));
   NOR2_X1 i_0_0_165 (.A1(n_0_0_36), .A2(n_0_0_1), .ZN(n_0_448));
   NOR2_X1 i_0_0_166 (.A1(n_0_0_36), .A2(n_0_0_2), .ZN(n_0_449));
   NOR2_X1 i_0_0_167 (.A1(n_0_0_36), .A2(n_0_0_3), .ZN(n_0_450));
   NOR2_X1 i_0_0_168 (.A1(n_0_0_36), .A2(n_0_0_4), .ZN(n_0_451));
   NOR2_X1 i_0_0_169 (.A1(n_0_0_36), .A2(n_0_0_5), .ZN(n_0_452));
   NOR2_X1 i_0_0_170 (.A1(n_0_0_36), .A2(n_0_0_6), .ZN(n_0_453));
   NOR2_X1 i_0_0_171 (.A1(n_0_0_36), .A2(n_0_0_7), .ZN(n_0_454));
   NOR2_X1 i_0_0_172 (.A1(n_0_0_36), .A2(n_0_0_8), .ZN(n_0_455));
   NOR2_X1 i_0_0_173 (.A1(n_0_0_36), .A2(n_0_0_9), .ZN(n_0_456));
   NOR2_X1 i_0_0_174 (.A1(n_0_0_36), .A2(n_0_0_10), .ZN(n_0_457));
   NOR2_X1 i_0_0_175 (.A1(n_0_0_36), .A2(n_0_0_11), .ZN(n_0_458));
   NOR2_X1 i_0_0_176 (.A1(n_0_0_36), .A2(n_0_0_12), .ZN(n_0_459));
   NOR2_X1 i_0_0_177 (.A1(n_0_0_36), .A2(n_0_0_13), .ZN(n_0_460));
   NOR2_X1 i_0_0_178 (.A1(n_0_0_36), .A2(n_0_0_14), .ZN(n_0_461));
   NOR2_X1 i_0_0_179 (.A1(n_0_0_36), .A2(n_0_0_15), .ZN(n_0_462));
   NOR2_X1 i_0_0_180 (.A1(n_0_0_36), .A2(n_0_0_16), .ZN(n_0_463));
   NOR2_X1 i_0_0_181 (.A1(n_0_0_36), .A2(n_0_0_17), .ZN(n_0_464));
   NOR2_X1 i_0_0_182 (.A1(n_0_0_36), .A2(n_0_0_18), .ZN(n_0_465));
   NOR2_X1 i_0_0_183 (.A1(n_0_0_36), .A2(n_0_0_19), .ZN(n_0_466));
   NOR2_X1 i_0_0_184 (.A1(n_0_0_36), .A2(n_0_0_20), .ZN(n_0_467));
   NOR2_X1 i_0_0_185 (.A1(n_0_0_36), .A2(n_0_0_21), .ZN(n_0_468));
   NOR2_X1 i_0_0_186 (.A1(n_0_0_36), .A2(n_0_0_22), .ZN(n_0_469));
   NOR2_X1 i_0_0_187 (.A1(n_0_0_36), .A2(n_0_0_23), .ZN(n_0_470));
   NOR2_X1 i_0_0_188 (.A1(n_0_0_36), .A2(n_0_0_24), .ZN(n_0_471));
   NOR2_X1 i_0_0_189 (.A1(n_0_0_36), .A2(n_0_0_25), .ZN(n_0_472));
   NOR2_X1 i_0_0_190 (.A1(n_0_0_36), .A2(n_0_0_26), .ZN(n_0_473));
   NOR2_X1 i_0_0_191 (.A1(n_0_0_36), .A2(n_0_0_27), .ZN(n_0_474));
   NOR2_X1 i_0_0_192 (.A1(n_0_0_36), .A2(n_0_0_28), .ZN(n_0_475));
   NOR2_X1 i_0_0_193 (.A1(n_0_0_36), .A2(n_0_0_29), .ZN(n_0_476));
   NOR2_X1 i_0_0_194 (.A1(n_0_0_36), .A2(n_0_0_30), .ZN(n_0_477));
   NOR2_X1 i_0_0_195 (.A1(n_0_0_36), .A2(n_0_0_31), .ZN(n_0_478));
   NOR2_X1 i_0_0_196 (.A1(n_0_0_36), .A2(n_0_0_32), .ZN(n_0_479));
   INV_X1 i_0_0_197 (.A(b[5]), .ZN(n_0_0_37));
   NOR2_X1 i_0_0_198 (.A1(n_0_0_37), .A2(n_0_0_1), .ZN(n_0_416));
   NOR2_X1 i_0_0_199 (.A1(n_0_0_37), .A2(n_0_0_2), .ZN(n_0_417));
   NOR2_X1 i_0_0_200 (.A1(n_0_0_37), .A2(n_0_0_3), .ZN(n_0_418));
   NOR2_X1 i_0_0_201 (.A1(n_0_0_37), .A2(n_0_0_4), .ZN(n_0_419));
   NOR2_X1 i_0_0_202 (.A1(n_0_0_37), .A2(n_0_0_5), .ZN(n_0_420));
   NOR2_X1 i_0_0_203 (.A1(n_0_0_37), .A2(n_0_0_6), .ZN(n_0_421));
   NOR2_X1 i_0_0_204 (.A1(n_0_0_37), .A2(n_0_0_7), .ZN(n_0_422));
   NOR2_X1 i_0_0_205 (.A1(n_0_0_37), .A2(n_0_0_8), .ZN(n_0_423));
   NOR2_X1 i_0_0_206 (.A1(n_0_0_37), .A2(n_0_0_9), .ZN(n_0_424));
   NOR2_X1 i_0_0_207 (.A1(n_0_0_37), .A2(n_0_0_10), .ZN(n_0_425));
   NOR2_X1 i_0_0_208 (.A1(n_0_0_37), .A2(n_0_0_11), .ZN(n_0_426));
   NOR2_X1 i_0_0_209 (.A1(n_0_0_37), .A2(n_0_0_12), .ZN(n_0_427));
   NOR2_X1 i_0_0_210 (.A1(n_0_0_37), .A2(n_0_0_13), .ZN(n_0_428));
   NOR2_X1 i_0_0_211 (.A1(n_0_0_37), .A2(n_0_0_14), .ZN(n_0_429));
   NOR2_X1 i_0_0_212 (.A1(n_0_0_37), .A2(n_0_0_15), .ZN(n_0_430));
   NOR2_X1 i_0_0_213 (.A1(n_0_0_37), .A2(n_0_0_16), .ZN(n_0_431));
   NOR2_X1 i_0_0_214 (.A1(n_0_0_37), .A2(n_0_0_17), .ZN(n_0_432));
   NOR2_X1 i_0_0_215 (.A1(n_0_0_37), .A2(n_0_0_18), .ZN(n_0_433));
   NOR2_X1 i_0_0_216 (.A1(n_0_0_37), .A2(n_0_0_19), .ZN(n_0_434));
   NOR2_X1 i_0_0_217 (.A1(n_0_0_37), .A2(n_0_0_20), .ZN(n_0_435));
   NOR2_X1 i_0_0_218 (.A1(n_0_0_37), .A2(n_0_0_21), .ZN(n_0_436));
   NOR2_X1 i_0_0_219 (.A1(n_0_0_37), .A2(n_0_0_22), .ZN(n_0_437));
   NOR2_X1 i_0_0_220 (.A1(n_0_0_37), .A2(n_0_0_23), .ZN(n_0_438));
   NOR2_X1 i_0_0_221 (.A1(n_0_0_37), .A2(n_0_0_24), .ZN(n_0_439));
   NOR2_X1 i_0_0_222 (.A1(n_0_0_37), .A2(n_0_0_25), .ZN(n_0_440));
   NOR2_X1 i_0_0_223 (.A1(n_0_0_37), .A2(n_0_0_26), .ZN(n_0_441));
   NOR2_X1 i_0_0_224 (.A1(n_0_0_37), .A2(n_0_0_27), .ZN(n_0_442));
   NOR2_X1 i_0_0_225 (.A1(n_0_0_37), .A2(n_0_0_28), .ZN(n_0_443));
   NOR2_X1 i_0_0_226 (.A1(n_0_0_37), .A2(n_0_0_29), .ZN(n_0_444));
   NOR2_X1 i_0_0_227 (.A1(n_0_0_37), .A2(n_0_0_30), .ZN(n_0_445));
   NOR2_X1 i_0_0_228 (.A1(n_0_0_37), .A2(n_0_0_31), .ZN(n_0_446));
   NOR2_X1 i_0_0_229 (.A1(n_0_0_37), .A2(n_0_0_32), .ZN(n_0_447));
   INV_X1 i_0_0_230 (.A(b[6]), .ZN(n_0_0_38));
   NOR2_X1 i_0_0_231 (.A1(n_0_0_38), .A2(n_0_0_1), .ZN(n_0_384));
   NOR2_X1 i_0_0_232 (.A1(n_0_0_38), .A2(n_0_0_2), .ZN(n_0_385));
   NOR2_X1 i_0_0_233 (.A1(n_0_0_38), .A2(n_0_0_3), .ZN(n_0_386));
   NOR2_X1 i_0_0_234 (.A1(n_0_0_38), .A2(n_0_0_4), .ZN(n_0_387));
   NOR2_X1 i_0_0_235 (.A1(n_0_0_38), .A2(n_0_0_5), .ZN(n_0_388));
   NOR2_X1 i_0_0_236 (.A1(n_0_0_38), .A2(n_0_0_6), .ZN(n_0_389));
   NOR2_X1 i_0_0_237 (.A1(n_0_0_38), .A2(n_0_0_7), .ZN(n_0_390));
   NOR2_X1 i_0_0_238 (.A1(n_0_0_38), .A2(n_0_0_8), .ZN(n_0_391));
   NOR2_X1 i_0_0_239 (.A1(n_0_0_38), .A2(n_0_0_9), .ZN(n_0_392));
   NOR2_X1 i_0_0_240 (.A1(n_0_0_38), .A2(n_0_0_10), .ZN(n_0_393));
   NOR2_X1 i_0_0_241 (.A1(n_0_0_38), .A2(n_0_0_11), .ZN(n_0_394));
   NOR2_X1 i_0_0_242 (.A1(n_0_0_38), .A2(n_0_0_12), .ZN(n_0_395));
   NOR2_X1 i_0_0_243 (.A1(n_0_0_38), .A2(n_0_0_13), .ZN(n_0_396));
   NOR2_X1 i_0_0_244 (.A1(n_0_0_38), .A2(n_0_0_14), .ZN(n_0_397));
   NOR2_X1 i_0_0_245 (.A1(n_0_0_38), .A2(n_0_0_15), .ZN(n_0_398));
   NOR2_X1 i_0_0_246 (.A1(n_0_0_38), .A2(n_0_0_16), .ZN(n_0_399));
   NOR2_X1 i_0_0_247 (.A1(n_0_0_38), .A2(n_0_0_17), .ZN(n_0_400));
   NOR2_X1 i_0_0_248 (.A1(n_0_0_38), .A2(n_0_0_18), .ZN(n_0_401));
   NOR2_X1 i_0_0_249 (.A1(n_0_0_38), .A2(n_0_0_19), .ZN(n_0_402));
   NOR2_X1 i_0_0_250 (.A1(n_0_0_38), .A2(n_0_0_20), .ZN(n_0_403));
   NOR2_X1 i_0_0_251 (.A1(n_0_0_38), .A2(n_0_0_21), .ZN(n_0_404));
   NOR2_X1 i_0_0_252 (.A1(n_0_0_38), .A2(n_0_0_22), .ZN(n_0_405));
   NOR2_X1 i_0_0_253 (.A1(n_0_0_38), .A2(n_0_0_23), .ZN(n_0_406));
   NOR2_X1 i_0_0_254 (.A1(n_0_0_38), .A2(n_0_0_24), .ZN(n_0_407));
   NOR2_X1 i_0_0_255 (.A1(n_0_0_38), .A2(n_0_0_25), .ZN(n_0_408));
   NOR2_X1 i_0_0_256 (.A1(n_0_0_38), .A2(n_0_0_26), .ZN(n_0_409));
   NOR2_X1 i_0_0_257 (.A1(n_0_0_38), .A2(n_0_0_27), .ZN(n_0_410));
   NOR2_X1 i_0_0_258 (.A1(n_0_0_38), .A2(n_0_0_28), .ZN(n_0_411));
   NOR2_X1 i_0_0_259 (.A1(n_0_0_38), .A2(n_0_0_29), .ZN(n_0_412));
   NOR2_X1 i_0_0_260 (.A1(n_0_0_38), .A2(n_0_0_30), .ZN(n_0_413));
   NOR2_X1 i_0_0_261 (.A1(n_0_0_38), .A2(n_0_0_31), .ZN(n_0_414));
   NOR2_X1 i_0_0_262 (.A1(n_0_0_38), .A2(n_0_0_32), .ZN(n_0_415));
   INV_X1 i_0_0_263 (.A(b[7]), .ZN(n_0_0_39));
   NOR2_X1 i_0_0_264 (.A1(n_0_0_39), .A2(n_0_0_1), .ZN(n_0_352));
   NOR2_X1 i_0_0_265 (.A1(n_0_0_39), .A2(n_0_0_2), .ZN(n_0_353));
   NOR2_X1 i_0_0_266 (.A1(n_0_0_39), .A2(n_0_0_3), .ZN(n_0_354));
   NOR2_X1 i_0_0_267 (.A1(n_0_0_39), .A2(n_0_0_4), .ZN(n_0_355));
   NOR2_X1 i_0_0_268 (.A1(n_0_0_39), .A2(n_0_0_5), .ZN(n_0_356));
   NOR2_X1 i_0_0_269 (.A1(n_0_0_39), .A2(n_0_0_6), .ZN(n_0_357));
   NOR2_X1 i_0_0_270 (.A1(n_0_0_39), .A2(n_0_0_7), .ZN(n_0_358));
   NOR2_X1 i_0_0_271 (.A1(n_0_0_39), .A2(n_0_0_8), .ZN(n_0_359));
   NOR2_X1 i_0_0_272 (.A1(n_0_0_39), .A2(n_0_0_9), .ZN(n_0_360));
   NOR2_X1 i_0_0_273 (.A1(n_0_0_39), .A2(n_0_0_10), .ZN(n_0_361));
   NOR2_X1 i_0_0_274 (.A1(n_0_0_39), .A2(n_0_0_11), .ZN(n_0_362));
   NOR2_X1 i_0_0_275 (.A1(n_0_0_39), .A2(n_0_0_12), .ZN(n_0_363));
   NOR2_X1 i_0_0_276 (.A1(n_0_0_39), .A2(n_0_0_13), .ZN(n_0_364));
   NOR2_X1 i_0_0_277 (.A1(n_0_0_39), .A2(n_0_0_14), .ZN(n_0_365));
   NOR2_X1 i_0_0_278 (.A1(n_0_0_39), .A2(n_0_0_15), .ZN(n_0_366));
   NOR2_X1 i_0_0_279 (.A1(n_0_0_39), .A2(n_0_0_16), .ZN(n_0_367));
   NOR2_X1 i_0_0_280 (.A1(n_0_0_39), .A2(n_0_0_17), .ZN(n_0_368));
   NOR2_X1 i_0_0_281 (.A1(n_0_0_39), .A2(n_0_0_18), .ZN(n_0_369));
   NOR2_X1 i_0_0_282 (.A1(n_0_0_39), .A2(n_0_0_19), .ZN(n_0_370));
   NOR2_X1 i_0_0_283 (.A1(n_0_0_39), .A2(n_0_0_20), .ZN(n_0_371));
   NOR2_X1 i_0_0_284 (.A1(n_0_0_39), .A2(n_0_0_21), .ZN(n_0_372));
   NOR2_X1 i_0_0_285 (.A1(n_0_0_39), .A2(n_0_0_22), .ZN(n_0_373));
   NOR2_X1 i_0_0_286 (.A1(n_0_0_39), .A2(n_0_0_23), .ZN(n_0_374));
   NOR2_X1 i_0_0_287 (.A1(n_0_0_39), .A2(n_0_0_24), .ZN(n_0_375));
   NOR2_X1 i_0_0_288 (.A1(n_0_0_39), .A2(n_0_0_25), .ZN(n_0_376));
   NOR2_X1 i_0_0_289 (.A1(n_0_0_39), .A2(n_0_0_26), .ZN(n_0_377));
   NOR2_X1 i_0_0_290 (.A1(n_0_0_39), .A2(n_0_0_27), .ZN(n_0_378));
   NOR2_X1 i_0_0_291 (.A1(n_0_0_39), .A2(n_0_0_28), .ZN(n_0_379));
   NOR2_X1 i_0_0_292 (.A1(n_0_0_39), .A2(n_0_0_29), .ZN(n_0_380));
   NOR2_X1 i_0_0_293 (.A1(n_0_0_39), .A2(n_0_0_30), .ZN(n_0_381));
   NOR2_X1 i_0_0_294 (.A1(n_0_0_39), .A2(n_0_0_31), .ZN(n_0_382));
   NOR2_X1 i_0_0_295 (.A1(n_0_0_39), .A2(n_0_0_32), .ZN(n_0_383));
   INV_X1 i_0_0_296 (.A(b[8]), .ZN(n_0_0_40));
   NOR2_X1 i_0_0_297 (.A1(n_0_0_40), .A2(n_0_0_1), .ZN(n_0_320));
   NOR2_X1 i_0_0_298 (.A1(n_0_0_40), .A2(n_0_0_2), .ZN(n_0_321));
   NOR2_X1 i_0_0_299 (.A1(n_0_0_40), .A2(n_0_0_3), .ZN(n_0_322));
   NOR2_X1 i_0_0_300 (.A1(n_0_0_40), .A2(n_0_0_4), .ZN(n_0_323));
   NOR2_X1 i_0_0_301 (.A1(n_0_0_40), .A2(n_0_0_5), .ZN(n_0_324));
   NOR2_X1 i_0_0_302 (.A1(n_0_0_40), .A2(n_0_0_6), .ZN(n_0_325));
   NOR2_X1 i_0_0_303 (.A1(n_0_0_40), .A2(n_0_0_7), .ZN(n_0_326));
   NOR2_X1 i_0_0_304 (.A1(n_0_0_40), .A2(n_0_0_8), .ZN(n_0_327));
   NOR2_X1 i_0_0_305 (.A1(n_0_0_40), .A2(n_0_0_9), .ZN(n_0_328));
   NOR2_X1 i_0_0_306 (.A1(n_0_0_40), .A2(n_0_0_10), .ZN(n_0_329));
   NOR2_X1 i_0_0_307 (.A1(n_0_0_40), .A2(n_0_0_11), .ZN(n_0_330));
   NOR2_X1 i_0_0_308 (.A1(n_0_0_40), .A2(n_0_0_12), .ZN(n_0_331));
   NOR2_X1 i_0_0_309 (.A1(n_0_0_40), .A2(n_0_0_13), .ZN(n_0_332));
   NOR2_X1 i_0_0_310 (.A1(n_0_0_40), .A2(n_0_0_14), .ZN(n_0_333));
   NOR2_X1 i_0_0_311 (.A1(n_0_0_40), .A2(n_0_0_15), .ZN(n_0_334));
   NOR2_X1 i_0_0_312 (.A1(n_0_0_40), .A2(n_0_0_16), .ZN(n_0_335));
   NOR2_X1 i_0_0_313 (.A1(n_0_0_40), .A2(n_0_0_17), .ZN(n_0_336));
   NOR2_X1 i_0_0_314 (.A1(n_0_0_40), .A2(n_0_0_18), .ZN(n_0_337));
   NOR2_X1 i_0_0_315 (.A1(n_0_0_40), .A2(n_0_0_19), .ZN(n_0_338));
   NOR2_X1 i_0_0_316 (.A1(n_0_0_40), .A2(n_0_0_20), .ZN(n_0_339));
   NOR2_X1 i_0_0_317 (.A1(n_0_0_40), .A2(n_0_0_21), .ZN(n_0_340));
   NOR2_X1 i_0_0_318 (.A1(n_0_0_40), .A2(n_0_0_22), .ZN(n_0_341));
   NOR2_X1 i_0_0_319 (.A1(n_0_0_40), .A2(n_0_0_23), .ZN(n_0_342));
   NOR2_X1 i_0_0_320 (.A1(n_0_0_40), .A2(n_0_0_24), .ZN(n_0_343));
   NOR2_X1 i_0_0_321 (.A1(n_0_0_40), .A2(n_0_0_25), .ZN(n_0_344));
   NOR2_X1 i_0_0_322 (.A1(n_0_0_40), .A2(n_0_0_26), .ZN(n_0_345));
   NOR2_X1 i_0_0_323 (.A1(n_0_0_40), .A2(n_0_0_27), .ZN(n_0_346));
   NOR2_X1 i_0_0_324 (.A1(n_0_0_40), .A2(n_0_0_28), .ZN(n_0_347));
   NOR2_X1 i_0_0_325 (.A1(n_0_0_40), .A2(n_0_0_29), .ZN(n_0_348));
   NOR2_X1 i_0_0_326 (.A1(n_0_0_40), .A2(n_0_0_30), .ZN(n_0_349));
   NOR2_X1 i_0_0_327 (.A1(n_0_0_40), .A2(n_0_0_31), .ZN(n_0_350));
   NOR2_X1 i_0_0_328 (.A1(n_0_0_40), .A2(n_0_0_32), .ZN(n_0_351));
   INV_X1 i_0_0_329 (.A(b[9]), .ZN(n_0_0_41));
   NOR2_X1 i_0_0_330 (.A1(n_0_0_41), .A2(n_0_0_1), .ZN(n_0_288));
   NOR2_X1 i_0_0_331 (.A1(n_0_0_41), .A2(n_0_0_2), .ZN(n_0_289));
   NOR2_X1 i_0_0_332 (.A1(n_0_0_41), .A2(n_0_0_3), .ZN(n_0_290));
   NOR2_X1 i_0_0_333 (.A1(n_0_0_41), .A2(n_0_0_4), .ZN(n_0_291));
   NOR2_X1 i_0_0_334 (.A1(n_0_0_41), .A2(n_0_0_5), .ZN(n_0_292));
   NOR2_X1 i_0_0_335 (.A1(n_0_0_41), .A2(n_0_0_6), .ZN(n_0_293));
   NOR2_X1 i_0_0_336 (.A1(n_0_0_41), .A2(n_0_0_7), .ZN(n_0_294));
   NOR2_X1 i_0_0_337 (.A1(n_0_0_41), .A2(n_0_0_8), .ZN(n_0_295));
   NOR2_X1 i_0_0_338 (.A1(n_0_0_41), .A2(n_0_0_9), .ZN(n_0_296));
   NOR2_X1 i_0_0_339 (.A1(n_0_0_41), .A2(n_0_0_10), .ZN(n_0_297));
   NOR2_X1 i_0_0_340 (.A1(n_0_0_41), .A2(n_0_0_11), .ZN(n_0_298));
   NOR2_X1 i_0_0_341 (.A1(n_0_0_41), .A2(n_0_0_12), .ZN(n_0_299));
   NOR2_X1 i_0_0_342 (.A1(n_0_0_41), .A2(n_0_0_13), .ZN(n_0_300));
   NOR2_X1 i_0_0_343 (.A1(n_0_0_41), .A2(n_0_0_14), .ZN(n_0_301));
   NOR2_X1 i_0_0_344 (.A1(n_0_0_41), .A2(n_0_0_15), .ZN(n_0_302));
   NOR2_X1 i_0_0_345 (.A1(n_0_0_41), .A2(n_0_0_16), .ZN(n_0_303));
   NOR2_X1 i_0_0_346 (.A1(n_0_0_41), .A2(n_0_0_17), .ZN(n_0_304));
   NOR2_X1 i_0_0_347 (.A1(n_0_0_41), .A2(n_0_0_18), .ZN(n_0_305));
   NOR2_X1 i_0_0_348 (.A1(n_0_0_41), .A2(n_0_0_19), .ZN(n_0_306));
   NOR2_X1 i_0_0_349 (.A1(n_0_0_41), .A2(n_0_0_20), .ZN(n_0_307));
   NOR2_X1 i_0_0_350 (.A1(n_0_0_41), .A2(n_0_0_21), .ZN(n_0_308));
   NOR2_X1 i_0_0_351 (.A1(n_0_0_41), .A2(n_0_0_22), .ZN(n_0_309));
   NOR2_X1 i_0_0_352 (.A1(n_0_0_41), .A2(n_0_0_23), .ZN(n_0_310));
   NOR2_X1 i_0_0_353 (.A1(n_0_0_41), .A2(n_0_0_24), .ZN(n_0_311));
   NOR2_X1 i_0_0_354 (.A1(n_0_0_41), .A2(n_0_0_25), .ZN(n_0_312));
   NOR2_X1 i_0_0_355 (.A1(n_0_0_41), .A2(n_0_0_26), .ZN(n_0_313));
   NOR2_X1 i_0_0_356 (.A1(n_0_0_41), .A2(n_0_0_27), .ZN(n_0_314));
   NOR2_X1 i_0_0_357 (.A1(n_0_0_41), .A2(n_0_0_28), .ZN(n_0_315));
   NOR2_X1 i_0_0_358 (.A1(n_0_0_41), .A2(n_0_0_29), .ZN(n_0_316));
   NOR2_X1 i_0_0_359 (.A1(n_0_0_41), .A2(n_0_0_30), .ZN(n_0_317));
   NOR2_X1 i_0_0_360 (.A1(n_0_0_41), .A2(n_0_0_31), .ZN(n_0_318));
   NOR2_X1 i_0_0_361 (.A1(n_0_0_41), .A2(n_0_0_32), .ZN(n_0_319));
   INV_X1 i_0_0_362 (.A(b[10]), .ZN(n_0_0_42));
   NOR2_X1 i_0_0_363 (.A1(n_0_0_42), .A2(n_0_0_1), .ZN(n_0_256));
   NOR2_X1 i_0_0_364 (.A1(n_0_0_42), .A2(n_0_0_2), .ZN(n_0_257));
   NOR2_X1 i_0_0_365 (.A1(n_0_0_42), .A2(n_0_0_3), .ZN(n_0_258));
   NOR2_X1 i_0_0_366 (.A1(n_0_0_42), .A2(n_0_0_4), .ZN(n_0_259));
   NOR2_X1 i_0_0_367 (.A1(n_0_0_42), .A2(n_0_0_5), .ZN(n_0_260));
   NOR2_X1 i_0_0_368 (.A1(n_0_0_42), .A2(n_0_0_6), .ZN(n_0_261));
   NOR2_X1 i_0_0_369 (.A1(n_0_0_42), .A2(n_0_0_7), .ZN(n_0_262));
   NOR2_X1 i_0_0_370 (.A1(n_0_0_42), .A2(n_0_0_8), .ZN(n_0_263));
   NOR2_X1 i_0_0_371 (.A1(n_0_0_42), .A2(n_0_0_9), .ZN(n_0_264));
   NOR2_X1 i_0_0_372 (.A1(n_0_0_42), .A2(n_0_0_10), .ZN(n_0_265));
   NOR2_X1 i_0_0_373 (.A1(n_0_0_42), .A2(n_0_0_11), .ZN(n_0_266));
   NOR2_X1 i_0_0_374 (.A1(n_0_0_42), .A2(n_0_0_12), .ZN(n_0_267));
   NOR2_X1 i_0_0_375 (.A1(n_0_0_42), .A2(n_0_0_13), .ZN(n_0_268));
   NOR2_X1 i_0_0_376 (.A1(n_0_0_42), .A2(n_0_0_14), .ZN(n_0_269));
   NOR2_X1 i_0_0_377 (.A1(n_0_0_42), .A2(n_0_0_15), .ZN(n_0_270));
   NOR2_X1 i_0_0_378 (.A1(n_0_0_42), .A2(n_0_0_16), .ZN(n_0_271));
   NOR2_X1 i_0_0_379 (.A1(n_0_0_42), .A2(n_0_0_17), .ZN(n_0_272));
   NOR2_X1 i_0_0_380 (.A1(n_0_0_42), .A2(n_0_0_18), .ZN(n_0_273));
   NOR2_X1 i_0_0_381 (.A1(n_0_0_42), .A2(n_0_0_19), .ZN(n_0_274));
   NOR2_X1 i_0_0_382 (.A1(n_0_0_42), .A2(n_0_0_20), .ZN(n_0_275));
   NOR2_X1 i_0_0_383 (.A1(n_0_0_42), .A2(n_0_0_21), .ZN(n_0_276));
   NOR2_X1 i_0_0_384 (.A1(n_0_0_42), .A2(n_0_0_22), .ZN(n_0_277));
   NOR2_X1 i_0_0_385 (.A1(n_0_0_42), .A2(n_0_0_23), .ZN(n_0_278));
   NOR2_X1 i_0_0_386 (.A1(n_0_0_42), .A2(n_0_0_24), .ZN(n_0_279));
   NOR2_X1 i_0_0_387 (.A1(n_0_0_42), .A2(n_0_0_25), .ZN(n_0_280));
   NOR2_X1 i_0_0_388 (.A1(n_0_0_42), .A2(n_0_0_26), .ZN(n_0_281));
   NOR2_X1 i_0_0_389 (.A1(n_0_0_42), .A2(n_0_0_27), .ZN(n_0_282));
   NOR2_X1 i_0_0_390 (.A1(n_0_0_42), .A2(n_0_0_28), .ZN(n_0_283));
   NOR2_X1 i_0_0_391 (.A1(n_0_0_42), .A2(n_0_0_29), .ZN(n_0_284));
   NOR2_X1 i_0_0_392 (.A1(n_0_0_42), .A2(n_0_0_30), .ZN(n_0_285));
   NOR2_X1 i_0_0_393 (.A1(n_0_0_42), .A2(n_0_0_31), .ZN(n_0_286));
   NOR2_X1 i_0_0_394 (.A1(n_0_0_42), .A2(n_0_0_32), .ZN(n_0_287));
   INV_X1 i_0_0_395 (.A(b[11]), .ZN(n_0_0_43));
   NOR2_X1 i_0_0_396 (.A1(n_0_0_43), .A2(n_0_0_1), .ZN(n_0_224));
   NOR2_X1 i_0_0_397 (.A1(n_0_0_43), .A2(n_0_0_2), .ZN(n_0_225));
   NOR2_X1 i_0_0_398 (.A1(n_0_0_43), .A2(n_0_0_3), .ZN(n_0_226));
   NOR2_X1 i_0_0_399 (.A1(n_0_0_43), .A2(n_0_0_4), .ZN(n_0_227));
   NOR2_X1 i_0_0_400 (.A1(n_0_0_43), .A2(n_0_0_5), .ZN(n_0_228));
   NOR2_X1 i_0_0_401 (.A1(n_0_0_43), .A2(n_0_0_6), .ZN(n_0_229));
   NOR2_X1 i_0_0_402 (.A1(n_0_0_43), .A2(n_0_0_7), .ZN(n_0_230));
   NOR2_X1 i_0_0_403 (.A1(n_0_0_43), .A2(n_0_0_8), .ZN(n_0_231));
   NOR2_X1 i_0_0_404 (.A1(n_0_0_43), .A2(n_0_0_9), .ZN(n_0_232));
   NOR2_X1 i_0_0_405 (.A1(n_0_0_43), .A2(n_0_0_10), .ZN(n_0_233));
   NOR2_X1 i_0_0_406 (.A1(n_0_0_43), .A2(n_0_0_11), .ZN(n_0_234));
   NOR2_X1 i_0_0_407 (.A1(n_0_0_43), .A2(n_0_0_12), .ZN(n_0_235));
   NOR2_X1 i_0_0_408 (.A1(n_0_0_43), .A2(n_0_0_13), .ZN(n_0_236));
   NOR2_X1 i_0_0_409 (.A1(n_0_0_43), .A2(n_0_0_14), .ZN(n_0_237));
   NOR2_X1 i_0_0_410 (.A1(n_0_0_43), .A2(n_0_0_15), .ZN(n_0_238));
   NOR2_X1 i_0_0_411 (.A1(n_0_0_43), .A2(n_0_0_16), .ZN(n_0_239));
   NOR2_X1 i_0_0_412 (.A1(n_0_0_43), .A2(n_0_0_17), .ZN(n_0_240));
   NOR2_X1 i_0_0_413 (.A1(n_0_0_43), .A2(n_0_0_18), .ZN(n_0_241));
   NOR2_X1 i_0_0_414 (.A1(n_0_0_43), .A2(n_0_0_19), .ZN(n_0_242));
   NOR2_X1 i_0_0_415 (.A1(n_0_0_43), .A2(n_0_0_20), .ZN(n_0_243));
   NOR2_X1 i_0_0_416 (.A1(n_0_0_43), .A2(n_0_0_21), .ZN(n_0_244));
   NOR2_X1 i_0_0_417 (.A1(n_0_0_43), .A2(n_0_0_22), .ZN(n_0_245));
   NOR2_X1 i_0_0_418 (.A1(n_0_0_43), .A2(n_0_0_23), .ZN(n_0_246));
   NOR2_X1 i_0_0_419 (.A1(n_0_0_43), .A2(n_0_0_24), .ZN(n_0_247));
   NOR2_X1 i_0_0_420 (.A1(n_0_0_43), .A2(n_0_0_25), .ZN(n_0_248));
   NOR2_X1 i_0_0_421 (.A1(n_0_0_43), .A2(n_0_0_26), .ZN(n_0_249));
   NOR2_X1 i_0_0_422 (.A1(n_0_0_43), .A2(n_0_0_27), .ZN(n_0_250));
   NOR2_X1 i_0_0_423 (.A1(n_0_0_43), .A2(n_0_0_28), .ZN(n_0_251));
   NOR2_X1 i_0_0_424 (.A1(n_0_0_43), .A2(n_0_0_29), .ZN(n_0_252));
   NOR2_X1 i_0_0_425 (.A1(n_0_0_43), .A2(n_0_0_30), .ZN(n_0_253));
   NOR2_X1 i_0_0_426 (.A1(n_0_0_43), .A2(n_0_0_31), .ZN(n_0_254));
   NOR2_X1 i_0_0_427 (.A1(n_0_0_43), .A2(n_0_0_32), .ZN(n_0_255));
   INV_X1 i_0_0_428 (.A(b[12]), .ZN(n_0_0_44));
   NOR2_X1 i_0_0_429 (.A1(n_0_0_44), .A2(n_0_0_1), .ZN(n_0_574));
   NOR2_X1 i_0_0_430 (.A1(n_0_0_44), .A2(n_0_0_2), .ZN(n_0));
   NOR2_X1 i_0_0_431 (.A1(n_0_0_44), .A2(n_0_0_3), .ZN(n_1));
   NOR2_X1 i_0_0_432 (.A1(n_0_0_44), .A2(n_0_0_4), .ZN(n_2));
   NOR2_X1 i_0_0_433 (.A1(n_0_0_44), .A2(n_0_0_5), .ZN(n_3));
   NOR2_X1 i_0_0_434 (.A1(n_0_0_44), .A2(n_0_0_6), .ZN(n_4));
   NOR2_X1 i_0_0_435 (.A1(n_0_0_44), .A2(n_0_0_7), .ZN(n_5));
   NOR2_X1 i_0_0_436 (.A1(n_0_0_44), .A2(n_0_0_8), .ZN(n_6));
   NOR2_X1 i_0_0_437 (.A1(n_0_0_44), .A2(n_0_0_9), .ZN(n_7));
   NOR2_X1 i_0_0_438 (.A1(n_0_0_44), .A2(n_0_0_10), .ZN(n_8));
   NOR2_X1 i_0_0_439 (.A1(n_0_0_44), .A2(n_0_0_11), .ZN(n_9));
   NOR2_X1 i_0_0_440 (.A1(n_0_0_44), .A2(n_0_0_12), .ZN(n_10));
   NOR2_X1 i_0_0_441 (.A1(n_0_0_44), .A2(n_0_0_13), .ZN(n_11));
   NOR2_X1 i_0_0_442 (.A1(n_0_0_44), .A2(n_0_0_14), .ZN(n_12));
   NOR2_X1 i_0_0_443 (.A1(n_0_0_44), .A2(n_0_0_15), .ZN(n_13));
   NOR2_X1 i_0_0_444 (.A1(n_0_0_44), .A2(n_0_0_16), .ZN(n_14));
   NOR2_X1 i_0_0_445 (.A1(n_0_0_44), .A2(n_0_0_17), .ZN(n_15));
   NOR2_X1 i_0_0_446 (.A1(n_0_0_44), .A2(n_0_0_18), .ZN(n_16));
   NOR2_X1 i_0_0_447 (.A1(n_0_0_44), .A2(n_0_0_19), .ZN(n_17));
   NOR2_X1 i_0_0_448 (.A1(n_0_0_44), .A2(n_0_0_20), .ZN(n_18));
   NOR2_X1 i_0_0_449 (.A1(n_0_0_44), .A2(n_0_0_21), .ZN(n_19));
   NOR2_X1 i_0_0_450 (.A1(n_0_0_44), .A2(n_0_0_22), .ZN(n_20));
   NOR2_X1 i_0_0_451 (.A1(n_0_0_44), .A2(n_0_0_23), .ZN(n_21));
   NOR2_X1 i_0_0_452 (.A1(n_0_0_44), .A2(n_0_0_24), .ZN(n_22));
   NOR2_X1 i_0_0_453 (.A1(n_0_0_44), .A2(n_0_0_25), .ZN(n_23));
   NOR2_X1 i_0_0_454 (.A1(n_0_0_44), .A2(n_0_0_26), .ZN(n_24));
   NOR2_X1 i_0_0_455 (.A1(n_0_0_44), .A2(n_0_0_27), .ZN(n_25));
   NOR2_X1 i_0_0_456 (.A1(n_0_0_44), .A2(n_0_0_28), .ZN(n_26));
   NOR2_X1 i_0_0_457 (.A1(n_0_0_44), .A2(n_0_0_29), .ZN(n_27));
   NOR2_X1 i_0_0_458 (.A1(n_0_0_44), .A2(n_0_0_30), .ZN(n_28));
   NOR2_X1 i_0_0_459 (.A1(n_0_0_44), .A2(n_0_0_31), .ZN(n_29));
   NOR2_X1 i_0_0_460 (.A1(n_0_0_44), .A2(n_0_0_32), .ZN(n_30));
   INV_X1 i_0_0_461 (.A(b[13]), .ZN(n_0_0_45));
   NOR2_X1 i_0_0_462 (.A1(n_0_0_45), .A2(n_0_0_1), .ZN(n_31));
   NOR2_X1 i_0_0_463 (.A1(n_0_0_45), .A2(n_0_0_2), .ZN(n_32));
   NOR2_X1 i_0_0_464 (.A1(n_0_0_45), .A2(n_0_0_3), .ZN(n_33));
   NOR2_X1 i_0_0_465 (.A1(n_0_0_45), .A2(n_0_0_4), .ZN(n_34));
   NOR2_X1 i_0_0_466 (.A1(n_0_0_45), .A2(n_0_0_5), .ZN(n_35));
   NOR2_X1 i_0_0_467 (.A1(n_0_0_45), .A2(n_0_0_6), .ZN(n_36));
   NOR2_X1 i_0_0_468 (.A1(n_0_0_45), .A2(n_0_0_7), .ZN(n_37));
   NOR2_X1 i_0_0_469 (.A1(n_0_0_45), .A2(n_0_0_8), .ZN(n_38));
   NOR2_X1 i_0_0_470 (.A1(n_0_0_45), .A2(n_0_0_9), .ZN(n_39));
   NOR2_X1 i_0_0_471 (.A1(n_0_0_45), .A2(n_0_0_10), .ZN(n_40));
   NOR2_X1 i_0_0_472 (.A1(n_0_0_45), .A2(n_0_0_11), .ZN(n_41));
   NOR2_X1 i_0_0_473 (.A1(n_0_0_45), .A2(n_0_0_12), .ZN(n_42));
   NOR2_X1 i_0_0_474 (.A1(n_0_0_45), .A2(n_0_0_13), .ZN(n_43));
   NOR2_X1 i_0_0_475 (.A1(n_0_0_45), .A2(n_0_0_14), .ZN(n_44));
   NOR2_X1 i_0_0_476 (.A1(n_0_0_45), .A2(n_0_0_15), .ZN(n_45));
   NOR2_X1 i_0_0_477 (.A1(n_0_0_45), .A2(n_0_0_16), .ZN(n_46));
   NOR2_X1 i_0_0_478 (.A1(n_0_0_45), .A2(n_0_0_17), .ZN(n_47));
   NOR2_X1 i_0_0_479 (.A1(n_0_0_45), .A2(n_0_0_18), .ZN(n_48));
   NOR2_X1 i_0_0_480 (.A1(n_0_0_45), .A2(n_0_0_19), .ZN(n_49));
   NOR2_X1 i_0_0_481 (.A1(n_0_0_45), .A2(n_0_0_20), .ZN(n_50));
   NOR2_X1 i_0_0_482 (.A1(n_0_0_45), .A2(n_0_0_21), .ZN(n_51));
   NOR2_X1 i_0_0_483 (.A1(n_0_0_45), .A2(n_0_0_22), .ZN(n_52));
   NOR2_X1 i_0_0_484 (.A1(n_0_0_45), .A2(n_0_0_23), .ZN(n_53));
   NOR2_X1 i_0_0_485 (.A1(n_0_0_45), .A2(n_0_0_24), .ZN(n_54));
   NOR2_X1 i_0_0_486 (.A1(n_0_0_45), .A2(n_0_0_25), .ZN(n_55));
   NOR2_X1 i_0_0_487 (.A1(n_0_0_45), .A2(n_0_0_26), .ZN(n_56));
   NOR2_X1 i_0_0_488 (.A1(n_0_0_45), .A2(n_0_0_27), .ZN(n_57));
   NOR2_X1 i_0_0_489 (.A1(n_0_0_45), .A2(n_0_0_28), .ZN(n_58));
   NOR2_X1 i_0_0_490 (.A1(n_0_0_45), .A2(n_0_0_29), .ZN(n_59));
   NOR2_X1 i_0_0_491 (.A1(n_0_0_45), .A2(n_0_0_30), .ZN(n_60));
   NOR2_X1 i_0_0_492 (.A1(n_0_0_45), .A2(n_0_0_31), .ZN(n_61));
   NOR2_X1 i_0_0_493 (.A1(n_0_0_45), .A2(n_0_0_32), .ZN(n_62));
   INV_X1 i_0_0_494 (.A(b[14]), .ZN(n_0_0_46));
   NOR2_X1 i_0_0_495 (.A1(n_0_0_46), .A2(n_0_0_1), .ZN(n_63));
   NOR2_X1 i_0_0_496 (.A1(n_0_0_46), .A2(n_0_0_2), .ZN(n_64));
   NOR2_X1 i_0_0_497 (.A1(n_0_0_46), .A2(n_0_0_3), .ZN(n_65));
   NOR2_X1 i_0_0_498 (.A1(n_0_0_46), .A2(n_0_0_4), .ZN(n_66));
   NOR2_X1 i_0_0_499 (.A1(n_0_0_46), .A2(n_0_0_5), .ZN(n_67));
   NOR2_X1 i_0_0_500 (.A1(n_0_0_46), .A2(n_0_0_6), .ZN(n_68));
   NOR2_X1 i_0_0_501 (.A1(n_0_0_46), .A2(n_0_0_7), .ZN(n_69));
   NOR2_X1 i_0_0_502 (.A1(n_0_0_46), .A2(n_0_0_8), .ZN(n_70));
   NOR2_X1 i_0_0_503 (.A1(n_0_0_46), .A2(n_0_0_9), .ZN(n_71));
   NOR2_X1 i_0_0_504 (.A1(n_0_0_46), .A2(n_0_0_10), .ZN(n_72));
   NOR2_X1 i_0_0_505 (.A1(n_0_0_46), .A2(n_0_0_11), .ZN(n_73));
   NOR2_X1 i_0_0_506 (.A1(n_0_0_46), .A2(n_0_0_12), .ZN(n_74));
   NOR2_X1 i_0_0_507 (.A1(n_0_0_46), .A2(n_0_0_13), .ZN(n_75));
   NOR2_X1 i_0_0_508 (.A1(n_0_0_46), .A2(n_0_0_14), .ZN(n_76));
   NOR2_X1 i_0_0_509 (.A1(n_0_0_46), .A2(n_0_0_15), .ZN(n_77));
   NOR2_X1 i_0_0_510 (.A1(n_0_0_46), .A2(n_0_0_16), .ZN(n_78));
   NOR2_X1 i_0_0_511 (.A1(n_0_0_46), .A2(n_0_0_17), .ZN(n_79));
   NOR2_X1 i_0_0_512 (.A1(n_0_0_46), .A2(n_0_0_18), .ZN(n_80));
   NOR2_X1 i_0_0_513 (.A1(n_0_0_46), .A2(n_0_0_19), .ZN(n_81));
   NOR2_X1 i_0_0_514 (.A1(n_0_0_46), .A2(n_0_0_20), .ZN(n_82));
   NOR2_X1 i_0_0_515 (.A1(n_0_0_46), .A2(n_0_0_21), .ZN(n_83));
   NOR2_X1 i_0_0_516 (.A1(n_0_0_46), .A2(n_0_0_22), .ZN(n_84));
   NOR2_X1 i_0_0_517 (.A1(n_0_0_46), .A2(n_0_0_23), .ZN(n_85));
   NOR2_X1 i_0_0_518 (.A1(n_0_0_46), .A2(n_0_0_24), .ZN(n_86));
   NOR2_X1 i_0_0_519 (.A1(n_0_0_46), .A2(n_0_0_25), .ZN(n_87));
   NOR2_X1 i_0_0_520 (.A1(n_0_0_46), .A2(n_0_0_26), .ZN(n_88));
   NOR2_X1 i_0_0_521 (.A1(n_0_0_46), .A2(n_0_0_27), .ZN(n_89));
   NOR2_X1 i_0_0_522 (.A1(n_0_0_46), .A2(n_0_0_28), .ZN(n_90));
   NOR2_X1 i_0_0_523 (.A1(n_0_0_46), .A2(n_0_0_29), .ZN(n_91));
   NOR2_X1 i_0_0_524 (.A1(n_0_0_46), .A2(n_0_0_30), .ZN(n_92));
   NOR2_X1 i_0_0_525 (.A1(n_0_0_46), .A2(n_0_0_31), .ZN(n_93));
   NOR2_X1 i_0_0_526 (.A1(n_0_0_46), .A2(n_0_0_32), .ZN(n_94));
   INV_X1 i_0_0_527 (.A(b[15]), .ZN(n_0_0_47));
   NOR2_X1 i_0_0_528 (.A1(n_0_0_47), .A2(n_0_0_1), .ZN(n_95));
   NOR2_X1 i_0_0_529 (.A1(n_0_0_47), .A2(n_0_0_2), .ZN(n_96));
   NOR2_X1 i_0_0_530 (.A1(n_0_0_47), .A2(n_0_0_3), .ZN(n_97));
   NOR2_X1 i_0_0_531 (.A1(n_0_0_47), .A2(n_0_0_4), .ZN(n_98));
   NOR2_X1 i_0_0_532 (.A1(n_0_0_47), .A2(n_0_0_5), .ZN(n_99));
   NOR2_X1 i_0_0_533 (.A1(n_0_0_47), .A2(n_0_0_6), .ZN(n_100));
   NOR2_X1 i_0_0_534 (.A1(n_0_0_47), .A2(n_0_0_7), .ZN(n_101));
   NOR2_X1 i_0_0_535 (.A1(n_0_0_47), .A2(n_0_0_8), .ZN(n_102));
   NOR2_X1 i_0_0_536 (.A1(n_0_0_47), .A2(n_0_0_9), .ZN(n_103));
   NOR2_X1 i_0_0_537 (.A1(n_0_0_47), .A2(n_0_0_10), .ZN(n_104));
   NOR2_X1 i_0_0_538 (.A1(n_0_0_47), .A2(n_0_0_11), .ZN(n_105));
   NOR2_X1 i_0_0_539 (.A1(n_0_0_47), .A2(n_0_0_12), .ZN(n_106));
   NOR2_X1 i_0_0_540 (.A1(n_0_0_47), .A2(n_0_0_13), .ZN(n_107));
   NOR2_X1 i_0_0_541 (.A1(n_0_0_47), .A2(n_0_0_14), .ZN(n_108));
   NOR2_X1 i_0_0_542 (.A1(n_0_0_47), .A2(n_0_0_15), .ZN(n_109));
   NOR2_X1 i_0_0_543 (.A1(n_0_0_47), .A2(n_0_0_16), .ZN(n_110));
   NOR2_X1 i_0_0_544 (.A1(n_0_0_47), .A2(n_0_0_17), .ZN(n_111));
   NOR2_X1 i_0_0_545 (.A1(n_0_0_47), .A2(n_0_0_18), .ZN(n_112));
   NOR2_X1 i_0_0_546 (.A1(n_0_0_47), .A2(n_0_0_19), .ZN(n_113));
   NOR2_X1 i_0_0_547 (.A1(n_0_0_47), .A2(n_0_0_20), .ZN(n_114));
   NOR2_X1 i_0_0_548 (.A1(n_0_0_47), .A2(n_0_0_21), .ZN(n_115));
   NOR2_X1 i_0_0_549 (.A1(n_0_0_47), .A2(n_0_0_22), .ZN(n_116));
   NOR2_X1 i_0_0_550 (.A1(n_0_0_47), .A2(n_0_0_23), .ZN(n_117));
   NOR2_X1 i_0_0_551 (.A1(n_0_0_47), .A2(n_0_0_24), .ZN(n_118));
   NOR2_X1 i_0_0_552 (.A1(n_0_0_47), .A2(n_0_0_25), .ZN(n_119));
   NOR2_X1 i_0_0_553 (.A1(n_0_0_47), .A2(n_0_0_26), .ZN(n_120));
   NOR2_X1 i_0_0_554 (.A1(n_0_0_47), .A2(n_0_0_27), .ZN(n_121));
   NOR2_X1 i_0_0_555 (.A1(n_0_0_47), .A2(n_0_0_28), .ZN(n_122));
   NOR2_X1 i_0_0_556 (.A1(n_0_0_47), .A2(n_0_0_29), .ZN(n_123));
   NOR2_X1 i_0_0_557 (.A1(n_0_0_47), .A2(n_0_0_30), .ZN(n_124));
   NOR2_X1 i_0_0_558 (.A1(n_0_0_47), .A2(n_0_0_31), .ZN(n_125));
   NOR2_X1 i_0_0_559 (.A1(n_0_0_47), .A2(n_0_0_32), .ZN(n_126));
   INV_X1 i_0_0_560 (.A(b[16]), .ZN(n_0_0_48));
   NOR2_X1 i_0_0_561 (.A1(n_0_0_48), .A2(n_0_0_1), .ZN(n_127));
   NOR2_X1 i_0_0_562 (.A1(n_0_0_48), .A2(n_0_0_2), .ZN(n_128));
   NOR2_X1 i_0_0_563 (.A1(n_0_0_48), .A2(n_0_0_3), .ZN(n_129));
   NOR2_X1 i_0_0_564 (.A1(n_0_0_48), .A2(n_0_0_4), .ZN(n_130));
   NOR2_X1 i_0_0_565 (.A1(n_0_0_48), .A2(n_0_0_5), .ZN(n_131));
   NOR2_X1 i_0_0_566 (.A1(n_0_0_48), .A2(n_0_0_6), .ZN(n_132));
   NOR2_X1 i_0_0_567 (.A1(n_0_0_48), .A2(n_0_0_7), .ZN(n_133));
   NOR2_X1 i_0_0_568 (.A1(n_0_0_48), .A2(n_0_0_8), .ZN(n_134));
   NOR2_X1 i_0_0_569 (.A1(n_0_0_48), .A2(n_0_0_9), .ZN(n_135));
   NOR2_X1 i_0_0_570 (.A1(n_0_0_48), .A2(n_0_0_10), .ZN(n_136));
   NOR2_X1 i_0_0_571 (.A1(n_0_0_48), .A2(n_0_0_11), .ZN(n_137));
   NOR2_X1 i_0_0_572 (.A1(n_0_0_48), .A2(n_0_0_12), .ZN(n_138));
   NOR2_X1 i_0_0_573 (.A1(n_0_0_48), .A2(n_0_0_13), .ZN(n_139));
   NOR2_X1 i_0_0_574 (.A1(n_0_0_48), .A2(n_0_0_14), .ZN(n_140));
   NOR2_X1 i_0_0_575 (.A1(n_0_0_48), .A2(n_0_0_15), .ZN(n_141));
   NOR2_X1 i_0_0_576 (.A1(n_0_0_48), .A2(n_0_0_16), .ZN(n_142));
   NOR2_X1 i_0_0_577 (.A1(n_0_0_48), .A2(n_0_0_17), .ZN(n_143));
   NOR2_X1 i_0_0_578 (.A1(n_0_0_48), .A2(n_0_0_18), .ZN(n_144));
   NOR2_X1 i_0_0_579 (.A1(n_0_0_48), .A2(n_0_0_19), .ZN(n_145));
   NOR2_X1 i_0_0_580 (.A1(n_0_0_48), .A2(n_0_0_20), .ZN(n_146));
   NOR2_X1 i_0_0_581 (.A1(n_0_0_48), .A2(n_0_0_21), .ZN(n_147));
   NOR2_X1 i_0_0_582 (.A1(n_0_0_48), .A2(n_0_0_22), .ZN(n_148));
   NOR2_X1 i_0_0_583 (.A1(n_0_0_48), .A2(n_0_0_23), .ZN(n_149));
   NOR2_X1 i_0_0_584 (.A1(n_0_0_48), .A2(n_0_0_24), .ZN(n_150));
   NOR2_X1 i_0_0_585 (.A1(n_0_0_48), .A2(n_0_0_25), .ZN(n_151));
   NOR2_X1 i_0_0_586 (.A1(n_0_0_48), .A2(n_0_0_26), .ZN(n_152));
   NOR2_X1 i_0_0_587 (.A1(n_0_0_48), .A2(n_0_0_27), .ZN(n_153));
   NOR2_X1 i_0_0_588 (.A1(n_0_0_48), .A2(n_0_0_28), .ZN(n_154));
   NOR2_X1 i_0_0_589 (.A1(n_0_0_48), .A2(n_0_0_29), .ZN(n_155));
   NOR2_X1 i_0_0_590 (.A1(n_0_0_48), .A2(n_0_0_30), .ZN(n_156));
   NOR2_X1 i_0_0_591 (.A1(n_0_0_48), .A2(n_0_0_31), .ZN(n_157));
   NOR2_X1 i_0_0_592 (.A1(n_0_0_48), .A2(n_0_0_32), .ZN(n_158));
   INV_X1 i_0_0_593 (.A(b[17]), .ZN(n_0_0_49));
   NOR2_X1 i_0_0_594 (.A1(n_0_0_49), .A2(n_0_0_1), .ZN(n_159));
   NOR2_X1 i_0_0_595 (.A1(n_0_0_49), .A2(n_0_0_2), .ZN(n_160));
   NOR2_X1 i_0_0_596 (.A1(n_0_0_49), .A2(n_0_0_3), .ZN(n_161));
   NOR2_X1 i_0_0_597 (.A1(n_0_0_49), .A2(n_0_0_4), .ZN(n_162));
   NOR2_X1 i_0_0_598 (.A1(n_0_0_49), .A2(n_0_0_5), .ZN(n_163));
   NOR2_X1 i_0_0_599 (.A1(n_0_0_49), .A2(n_0_0_6), .ZN(n_164));
   NOR2_X1 i_0_0_600 (.A1(n_0_0_49), .A2(n_0_0_7), .ZN(n_165));
   NOR2_X1 i_0_0_601 (.A1(n_0_0_49), .A2(n_0_0_8), .ZN(n_166));
   NOR2_X1 i_0_0_602 (.A1(n_0_0_49), .A2(n_0_0_9), .ZN(n_167));
   NOR2_X1 i_0_0_603 (.A1(n_0_0_49), .A2(n_0_0_10), .ZN(n_168));
   NOR2_X1 i_0_0_604 (.A1(n_0_0_49), .A2(n_0_0_11), .ZN(n_169));
   NOR2_X1 i_0_0_605 (.A1(n_0_0_49), .A2(n_0_0_12), .ZN(n_170));
   NOR2_X1 i_0_0_606 (.A1(n_0_0_49), .A2(n_0_0_13), .ZN(n_171));
   NOR2_X1 i_0_0_607 (.A1(n_0_0_49), .A2(n_0_0_14), .ZN(n_172));
   NOR2_X1 i_0_0_608 (.A1(n_0_0_49), .A2(n_0_0_15), .ZN(n_173));
   NOR2_X1 i_0_0_609 (.A1(n_0_0_49), .A2(n_0_0_16), .ZN(n_174));
   NOR2_X1 i_0_0_610 (.A1(n_0_0_49), .A2(n_0_0_17), .ZN(n_175));
   NOR2_X1 i_0_0_611 (.A1(n_0_0_49), .A2(n_0_0_18), .ZN(n_176));
   NOR2_X1 i_0_0_612 (.A1(n_0_0_49), .A2(n_0_0_19), .ZN(n_177));
   NOR2_X1 i_0_0_613 (.A1(n_0_0_49), .A2(n_0_0_20), .ZN(n_178));
   NOR2_X1 i_0_0_614 (.A1(n_0_0_49), .A2(n_0_0_21), .ZN(n_179));
   NOR2_X1 i_0_0_615 (.A1(n_0_0_49), .A2(n_0_0_22), .ZN(n_180));
   NOR2_X1 i_0_0_616 (.A1(n_0_0_49), .A2(n_0_0_23), .ZN(n_181));
   NOR2_X1 i_0_0_617 (.A1(n_0_0_49), .A2(n_0_0_24), .ZN(n_182));
   NOR2_X1 i_0_0_618 (.A1(n_0_0_49), .A2(n_0_0_25), .ZN(n_183));
   NOR2_X1 i_0_0_619 (.A1(n_0_0_49), .A2(n_0_0_26), .ZN(n_184));
   NOR2_X1 i_0_0_620 (.A1(n_0_0_49), .A2(n_0_0_27), .ZN(n_185));
   NOR2_X1 i_0_0_621 (.A1(n_0_0_49), .A2(n_0_0_28), .ZN(n_186));
   NOR2_X1 i_0_0_622 (.A1(n_0_0_49), .A2(n_0_0_29), .ZN(n_187));
   NOR2_X1 i_0_0_623 (.A1(n_0_0_49), .A2(n_0_0_30), .ZN(n_188));
   NOR2_X1 i_0_0_624 (.A1(n_0_0_49), .A2(n_0_0_31), .ZN(n_189));
   NOR2_X1 i_0_0_625 (.A1(n_0_0_49), .A2(n_0_0_32), .ZN(n_190));
   INV_X1 i_0_0_626 (.A(b[18]), .ZN(n_0_0_50));
   NOR2_X1 i_0_0_627 (.A1(n_0_0_50), .A2(n_0_0_1), .ZN(n_191));
   NOR2_X1 i_0_0_628 (.A1(n_0_0_50), .A2(n_0_0_2), .ZN(n_192));
   NOR2_X1 i_0_0_629 (.A1(n_0_0_50), .A2(n_0_0_3), .ZN(n_193));
   NOR2_X1 i_0_0_630 (.A1(n_0_0_50), .A2(n_0_0_4), .ZN(n_194));
   NOR2_X1 i_0_0_631 (.A1(n_0_0_50), .A2(n_0_0_5), .ZN(n_195));
   NOR2_X1 i_0_0_632 (.A1(n_0_0_50), .A2(n_0_0_6), .ZN(n_196));
   NOR2_X1 i_0_0_633 (.A1(n_0_0_50), .A2(n_0_0_7), .ZN(n_197));
   NOR2_X1 i_0_0_634 (.A1(n_0_0_50), .A2(n_0_0_8), .ZN(n_198));
   NOR2_X1 i_0_0_635 (.A1(n_0_0_50), .A2(n_0_0_9), .ZN(n_199));
   NOR2_X1 i_0_0_636 (.A1(n_0_0_50), .A2(n_0_0_10), .ZN(n_200));
   NOR2_X1 i_0_0_637 (.A1(n_0_0_50), .A2(n_0_0_11), .ZN(n_201));
   NOR2_X1 i_0_0_638 (.A1(n_0_0_50), .A2(n_0_0_12), .ZN(n_202));
   NOR2_X1 i_0_0_639 (.A1(n_0_0_50), .A2(n_0_0_13), .ZN(n_203));
   NOR2_X1 i_0_0_640 (.A1(n_0_0_50), .A2(n_0_0_14), .ZN(n_204));
   NOR2_X1 i_0_0_641 (.A1(n_0_0_50), .A2(n_0_0_15), .ZN(n_205));
   NOR2_X1 i_0_0_642 (.A1(n_0_0_50), .A2(n_0_0_16), .ZN(n_206));
   NOR2_X1 i_0_0_643 (.A1(n_0_0_50), .A2(n_0_0_17), .ZN(n_207));
   NOR2_X1 i_0_0_644 (.A1(n_0_0_50), .A2(n_0_0_18), .ZN(n_208));
   NOR2_X1 i_0_0_645 (.A1(n_0_0_50), .A2(n_0_0_19), .ZN(n_209));
   NOR2_X1 i_0_0_646 (.A1(n_0_0_50), .A2(n_0_0_20), .ZN(n_210));
   NOR2_X1 i_0_0_647 (.A1(n_0_0_50), .A2(n_0_0_21), .ZN(n_211));
   NOR2_X1 i_0_0_648 (.A1(n_0_0_50), .A2(n_0_0_22), .ZN(n_212));
   NOR2_X1 i_0_0_649 (.A1(n_0_0_50), .A2(n_0_0_23), .ZN(n_213));
   NOR2_X1 i_0_0_650 (.A1(n_0_0_50), .A2(n_0_0_24), .ZN(n_214));
   NOR2_X1 i_0_0_651 (.A1(n_0_0_50), .A2(n_0_0_25), .ZN(n_215));
   NOR2_X1 i_0_0_652 (.A1(n_0_0_50), .A2(n_0_0_26), .ZN(n_216));
   NOR2_X1 i_0_0_653 (.A1(n_0_0_50), .A2(n_0_0_27), .ZN(n_217));
   NOR2_X1 i_0_0_654 (.A1(n_0_0_50), .A2(n_0_0_28), .ZN(n_218));
   NOR2_X1 i_0_0_655 (.A1(n_0_0_50), .A2(n_0_0_29), .ZN(n_219));
   NOR2_X1 i_0_0_656 (.A1(n_0_0_50), .A2(n_0_0_30), .ZN(n_220));
   NOR2_X1 i_0_0_657 (.A1(n_0_0_50), .A2(n_0_0_31), .ZN(n_221));
   NOR2_X1 i_0_0_658 (.A1(n_0_0_50), .A2(n_0_0_32), .ZN(n_222));
   INV_X1 i_0_0_659 (.A(b[19]), .ZN(n_0_0_51));
   NOR2_X1 i_0_0_660 (.A1(n_0_0_51), .A2(n_0_0_1), .ZN(n_223));
   NOR2_X1 i_0_0_661 (.A1(n_0_0_51), .A2(n_0_0_2), .ZN(n_224));
   NOR2_X1 i_0_0_662 (.A1(n_0_0_51), .A2(n_0_0_3), .ZN(n_225));
   NOR2_X1 i_0_0_663 (.A1(n_0_0_51), .A2(n_0_0_4), .ZN(n_226));
   NOR2_X1 i_0_0_664 (.A1(n_0_0_51), .A2(n_0_0_5), .ZN(n_227));
   NOR2_X1 i_0_0_665 (.A1(n_0_0_51), .A2(n_0_0_6), .ZN(n_228));
   NOR2_X1 i_0_0_666 (.A1(n_0_0_51), .A2(n_0_0_7), .ZN(n_229));
   NOR2_X1 i_0_0_667 (.A1(n_0_0_51), .A2(n_0_0_8), .ZN(n_230));
   NOR2_X1 i_0_0_668 (.A1(n_0_0_51), .A2(n_0_0_9), .ZN(n_231));
   NOR2_X1 i_0_0_669 (.A1(n_0_0_51), .A2(n_0_0_10), .ZN(n_232));
   NOR2_X1 i_0_0_670 (.A1(n_0_0_51), .A2(n_0_0_11), .ZN(n_233));
   NOR2_X1 i_0_0_671 (.A1(n_0_0_51), .A2(n_0_0_12), .ZN(n_234));
   NOR2_X1 i_0_0_672 (.A1(n_0_0_51), .A2(n_0_0_13), .ZN(n_235));
   NOR2_X1 i_0_0_673 (.A1(n_0_0_51), .A2(n_0_0_14), .ZN(n_236));
   NOR2_X1 i_0_0_674 (.A1(n_0_0_51), .A2(n_0_0_15), .ZN(n_237));
   NOR2_X1 i_0_0_675 (.A1(n_0_0_51), .A2(n_0_0_16), .ZN(n_238));
   NOR2_X1 i_0_0_676 (.A1(n_0_0_51), .A2(n_0_0_17), .ZN(n_239));
   NOR2_X1 i_0_0_677 (.A1(n_0_0_51), .A2(n_0_0_18), .ZN(n_240));
   NOR2_X1 i_0_0_678 (.A1(n_0_0_51), .A2(n_0_0_19), .ZN(n_241));
   NOR2_X1 i_0_0_679 (.A1(n_0_0_51), .A2(n_0_0_20), .ZN(n_242));
   NOR2_X1 i_0_0_680 (.A1(n_0_0_51), .A2(n_0_0_21), .ZN(n_243));
   NOR2_X1 i_0_0_681 (.A1(n_0_0_51), .A2(n_0_0_22), .ZN(n_244));
   NOR2_X1 i_0_0_682 (.A1(n_0_0_51), .A2(n_0_0_23), .ZN(n_245));
   NOR2_X1 i_0_0_683 (.A1(n_0_0_51), .A2(n_0_0_24), .ZN(n_246));
   NOR2_X1 i_0_0_684 (.A1(n_0_0_51), .A2(n_0_0_25), .ZN(n_247));
   NOR2_X1 i_0_0_685 (.A1(n_0_0_51), .A2(n_0_0_26), .ZN(n_248));
   NOR2_X1 i_0_0_686 (.A1(n_0_0_51), .A2(n_0_0_27), .ZN(n_249));
   NOR2_X1 i_0_0_687 (.A1(n_0_0_51), .A2(n_0_0_28), .ZN(n_250));
   NOR2_X1 i_0_0_688 (.A1(n_0_0_51), .A2(n_0_0_29), .ZN(n_251));
   NOR2_X1 i_0_0_689 (.A1(n_0_0_51), .A2(n_0_0_30), .ZN(n_252));
   NOR2_X1 i_0_0_690 (.A1(n_0_0_51), .A2(n_0_0_31), .ZN(n_253));
   NOR2_X1 i_0_0_691 (.A1(n_0_0_51), .A2(n_0_0_32), .ZN(n_254));
   INV_X1 i_0_0_692 (.A(b[20]), .ZN(n_0_0_52));
   NOR2_X1 i_0_0_693 (.A1(n_0_0_52), .A2(n_0_0_1), .ZN(n_255));
   NOR2_X1 i_0_0_694 (.A1(n_0_0_52), .A2(n_0_0_2), .ZN(n_256));
   NOR2_X1 i_0_0_695 (.A1(n_0_0_52), .A2(n_0_0_3), .ZN(n_257));
   NOR2_X1 i_0_0_696 (.A1(n_0_0_52), .A2(n_0_0_4), .ZN(n_258));
   NOR2_X1 i_0_0_697 (.A1(n_0_0_52), .A2(n_0_0_5), .ZN(n_259));
   NOR2_X1 i_0_0_698 (.A1(n_0_0_52), .A2(n_0_0_6), .ZN(n_260));
   NOR2_X1 i_0_0_699 (.A1(n_0_0_52), .A2(n_0_0_7), .ZN(n_261));
   NOR2_X1 i_0_0_700 (.A1(n_0_0_52), .A2(n_0_0_8), .ZN(n_262));
   NOR2_X1 i_0_0_701 (.A1(n_0_0_52), .A2(n_0_0_9), .ZN(n_263));
   NOR2_X1 i_0_0_702 (.A1(n_0_0_52), .A2(n_0_0_10), .ZN(n_264));
   NOR2_X1 i_0_0_703 (.A1(n_0_0_52), .A2(n_0_0_11), .ZN(n_265));
   NOR2_X1 i_0_0_704 (.A1(n_0_0_52), .A2(n_0_0_12), .ZN(n_266));
   NOR2_X1 i_0_0_705 (.A1(n_0_0_52), .A2(n_0_0_13), .ZN(n_267));
   NOR2_X1 i_0_0_706 (.A1(n_0_0_52), .A2(n_0_0_14), .ZN(n_268));
   NOR2_X1 i_0_0_707 (.A1(n_0_0_52), .A2(n_0_0_15), .ZN(n_269));
   NOR2_X1 i_0_0_708 (.A1(n_0_0_52), .A2(n_0_0_16), .ZN(n_270));
   NOR2_X1 i_0_0_709 (.A1(n_0_0_52), .A2(n_0_0_17), .ZN(n_271));
   NOR2_X1 i_0_0_710 (.A1(n_0_0_52), .A2(n_0_0_18), .ZN(n_272));
   NOR2_X1 i_0_0_711 (.A1(n_0_0_52), .A2(n_0_0_19), .ZN(n_273));
   NOR2_X1 i_0_0_712 (.A1(n_0_0_52), .A2(n_0_0_20), .ZN(n_274));
   NOR2_X1 i_0_0_713 (.A1(n_0_0_52), .A2(n_0_0_21), .ZN(n_275));
   NOR2_X1 i_0_0_714 (.A1(n_0_0_52), .A2(n_0_0_22), .ZN(n_276));
   NOR2_X1 i_0_0_715 (.A1(n_0_0_52), .A2(n_0_0_23), .ZN(n_277));
   NOR2_X1 i_0_0_716 (.A1(n_0_0_52), .A2(n_0_0_24), .ZN(n_278));
   NOR2_X1 i_0_0_717 (.A1(n_0_0_52), .A2(n_0_0_25), .ZN(n_279));
   NOR2_X1 i_0_0_718 (.A1(n_0_0_52), .A2(n_0_0_26), .ZN(n_280));
   NOR2_X1 i_0_0_719 (.A1(n_0_0_52), .A2(n_0_0_27), .ZN(n_281));
   NOR2_X1 i_0_0_720 (.A1(n_0_0_52), .A2(n_0_0_28), .ZN(n_282));
   NOR2_X1 i_0_0_721 (.A1(n_0_0_52), .A2(n_0_0_29), .ZN(n_283));
   NOR2_X1 i_0_0_722 (.A1(n_0_0_52), .A2(n_0_0_30), .ZN(n_284));
   NOR2_X1 i_0_0_723 (.A1(n_0_0_52), .A2(n_0_0_31), .ZN(n_285));
   NOR2_X1 i_0_0_724 (.A1(n_0_0_52), .A2(n_0_0_32), .ZN(n_286));
   INV_X1 i_0_0_725 (.A(b[21]), .ZN(n_0_0_53));
   NOR2_X1 i_0_0_726 (.A1(n_0_0_53), .A2(n_0_0_1), .ZN(\s1[7] [21]));
   NOR2_X1 i_0_0_727 (.A1(n_0_0_53), .A2(n_0_0_2), .ZN(n_0_193));
   NOR2_X1 i_0_0_728 (.A1(n_0_0_53), .A2(n_0_0_3), .ZN(n_0_194));
   NOR2_X1 i_0_0_729 (.A1(n_0_0_53), .A2(n_0_0_4), .ZN(n_0_195));
   NOR2_X1 i_0_0_730 (.A1(n_0_0_53), .A2(n_0_0_5), .ZN(n_0_196));
   NOR2_X1 i_0_0_731 (.A1(n_0_0_53), .A2(n_0_0_6), .ZN(n_0_197));
   NOR2_X1 i_0_0_732 (.A1(n_0_0_53), .A2(n_0_0_7), .ZN(n_0_198));
   NOR2_X1 i_0_0_733 (.A1(n_0_0_53), .A2(n_0_0_8), .ZN(n_0_199));
   NOR2_X1 i_0_0_734 (.A1(n_0_0_53), .A2(n_0_0_9), .ZN(n_0_200));
   NOR2_X1 i_0_0_735 (.A1(n_0_0_53), .A2(n_0_0_10), .ZN(n_0_201));
   NOR2_X1 i_0_0_736 (.A1(n_0_0_53), .A2(n_0_0_11), .ZN(n_0_202));
   NOR2_X1 i_0_0_737 (.A1(n_0_0_53), .A2(n_0_0_12), .ZN(n_0_203));
   NOR2_X1 i_0_0_738 (.A1(n_0_0_53), .A2(n_0_0_13), .ZN(n_0_204));
   NOR2_X1 i_0_0_739 (.A1(n_0_0_53), .A2(n_0_0_14), .ZN(n_0_205));
   NOR2_X1 i_0_0_740 (.A1(n_0_0_53), .A2(n_0_0_15), .ZN(n_0_206));
   NOR2_X1 i_0_0_741 (.A1(n_0_0_53), .A2(n_0_0_16), .ZN(n_0_207));
   NOR2_X1 i_0_0_742 (.A1(n_0_0_53), .A2(n_0_0_17), .ZN(n_0_208));
   NOR2_X1 i_0_0_743 (.A1(n_0_0_53), .A2(n_0_0_18), .ZN(n_0_209));
   NOR2_X1 i_0_0_744 (.A1(n_0_0_53), .A2(n_0_0_19), .ZN(n_0_210));
   NOR2_X1 i_0_0_745 (.A1(n_0_0_53), .A2(n_0_0_20), .ZN(n_0_211));
   NOR2_X1 i_0_0_746 (.A1(n_0_0_53), .A2(n_0_0_21), .ZN(n_0_212));
   NOR2_X1 i_0_0_747 (.A1(n_0_0_53), .A2(n_0_0_22), .ZN(n_0_213));
   NOR2_X1 i_0_0_748 (.A1(n_0_0_53), .A2(n_0_0_23), .ZN(n_0_214));
   NOR2_X1 i_0_0_749 (.A1(n_0_0_53), .A2(n_0_0_24), .ZN(n_0_215));
   NOR2_X1 i_0_0_750 (.A1(n_0_0_53), .A2(n_0_0_25), .ZN(n_0_216));
   NOR2_X1 i_0_0_751 (.A1(n_0_0_53), .A2(n_0_0_26), .ZN(n_0_217));
   NOR2_X1 i_0_0_752 (.A1(n_0_0_53), .A2(n_0_0_27), .ZN(n_0_218));
   NOR2_X1 i_0_0_753 (.A1(n_0_0_53), .A2(n_0_0_28), .ZN(n_0_219));
   NOR2_X1 i_0_0_754 (.A1(n_0_0_53), .A2(n_0_0_29), .ZN(n_0_220));
   NOR2_X1 i_0_0_755 (.A1(n_0_0_53), .A2(n_0_0_30), .ZN(n_0_221));
   NOR2_X1 i_0_0_756 (.A1(n_0_0_53), .A2(n_0_0_31), .ZN(n_0_222));
   NOR2_X1 i_0_0_757 (.A1(n_0_0_53), .A2(n_0_0_32), .ZN(n_0_223));
   INV_X1 i_0_0_758 (.A(b[22]), .ZN(n_0_0_54));
   NOR2_X1 i_0_0_759 (.A1(n_0_0_54), .A2(n_0_0_1), .ZN(n_0_160));
   NOR2_X1 i_0_0_760 (.A1(n_0_0_54), .A2(n_0_0_2), .ZN(n_0_161));
   NOR2_X1 i_0_0_761 (.A1(n_0_0_54), .A2(n_0_0_3), .ZN(n_0_162));
   NOR2_X1 i_0_0_762 (.A1(n_0_0_54), .A2(n_0_0_4), .ZN(n_0_163));
   NOR2_X1 i_0_0_763 (.A1(n_0_0_54), .A2(n_0_0_5), .ZN(n_0_164));
   NOR2_X1 i_0_0_764 (.A1(n_0_0_54), .A2(n_0_0_6), .ZN(n_0_165));
   NOR2_X1 i_0_0_765 (.A1(n_0_0_54), .A2(n_0_0_7), .ZN(n_0_166));
   NOR2_X1 i_0_0_766 (.A1(n_0_0_54), .A2(n_0_0_8), .ZN(n_0_167));
   NOR2_X1 i_0_0_767 (.A1(n_0_0_54), .A2(n_0_0_9), .ZN(n_0_168));
   NOR2_X1 i_0_0_768 (.A1(n_0_0_54), .A2(n_0_0_10), .ZN(n_0_169));
   NOR2_X1 i_0_0_769 (.A1(n_0_0_54), .A2(n_0_0_11), .ZN(n_0_170));
   NOR2_X1 i_0_0_770 (.A1(n_0_0_54), .A2(n_0_0_12), .ZN(n_0_171));
   NOR2_X1 i_0_0_771 (.A1(n_0_0_54), .A2(n_0_0_13), .ZN(n_0_172));
   NOR2_X1 i_0_0_772 (.A1(n_0_0_54), .A2(n_0_0_14), .ZN(n_0_173));
   NOR2_X1 i_0_0_773 (.A1(n_0_0_54), .A2(n_0_0_15), .ZN(n_0_174));
   NOR2_X1 i_0_0_774 (.A1(n_0_0_54), .A2(n_0_0_16), .ZN(n_0_175));
   NOR2_X1 i_0_0_775 (.A1(n_0_0_54), .A2(n_0_0_17), .ZN(n_0_176));
   NOR2_X1 i_0_0_776 (.A1(n_0_0_54), .A2(n_0_0_18), .ZN(n_0_177));
   NOR2_X1 i_0_0_777 (.A1(n_0_0_54), .A2(n_0_0_19), .ZN(n_0_178));
   NOR2_X1 i_0_0_778 (.A1(n_0_0_54), .A2(n_0_0_20), .ZN(n_0_179));
   NOR2_X1 i_0_0_779 (.A1(n_0_0_54), .A2(n_0_0_21), .ZN(n_0_180));
   NOR2_X1 i_0_0_780 (.A1(n_0_0_54), .A2(n_0_0_22), .ZN(n_0_181));
   NOR2_X1 i_0_0_781 (.A1(n_0_0_54), .A2(n_0_0_23), .ZN(n_0_182));
   NOR2_X1 i_0_0_782 (.A1(n_0_0_54), .A2(n_0_0_24), .ZN(n_0_183));
   NOR2_X1 i_0_0_783 (.A1(n_0_0_54), .A2(n_0_0_25), .ZN(n_0_184));
   NOR2_X1 i_0_0_784 (.A1(n_0_0_54), .A2(n_0_0_26), .ZN(n_0_185));
   NOR2_X1 i_0_0_785 (.A1(n_0_0_54), .A2(n_0_0_27), .ZN(n_0_186));
   NOR2_X1 i_0_0_786 (.A1(n_0_0_54), .A2(n_0_0_28), .ZN(n_0_187));
   NOR2_X1 i_0_0_787 (.A1(n_0_0_54), .A2(n_0_0_29), .ZN(n_0_188));
   NOR2_X1 i_0_0_788 (.A1(n_0_0_54), .A2(n_0_0_30), .ZN(n_0_189));
   NOR2_X1 i_0_0_789 (.A1(n_0_0_54), .A2(n_0_0_31), .ZN(n_0_190));
   NOR2_X1 i_0_0_790 (.A1(n_0_0_54), .A2(n_0_0_32), .ZN(n_0_191));
   INV_X1 i_0_0_791 (.A(b[23]), .ZN(n_0_0_55));
   NOR2_X1 i_0_0_792 (.A1(n_0_0_55), .A2(n_0_0_1), .ZN(n_0_128));
   NOR2_X1 i_0_0_793 (.A1(n_0_0_55), .A2(n_0_0_2), .ZN(n_0_129));
   NOR2_X1 i_0_0_794 (.A1(n_0_0_55), .A2(n_0_0_3), .ZN(n_0_130));
   NOR2_X1 i_0_0_795 (.A1(n_0_0_55), .A2(n_0_0_4), .ZN(n_0_131));
   NOR2_X1 i_0_0_796 (.A1(n_0_0_55), .A2(n_0_0_5), .ZN(n_0_132));
   NOR2_X1 i_0_0_797 (.A1(n_0_0_55), .A2(n_0_0_6), .ZN(n_0_133));
   NOR2_X1 i_0_0_798 (.A1(n_0_0_55), .A2(n_0_0_7), .ZN(n_0_134));
   NOR2_X1 i_0_0_799 (.A1(n_0_0_55), .A2(n_0_0_8), .ZN(n_0_135));
   NOR2_X1 i_0_0_800 (.A1(n_0_0_55), .A2(n_0_0_9), .ZN(n_0_136));
   NOR2_X1 i_0_0_801 (.A1(n_0_0_55), .A2(n_0_0_10), .ZN(n_0_137));
   NOR2_X1 i_0_0_802 (.A1(n_0_0_55), .A2(n_0_0_11), .ZN(n_0_138));
   NOR2_X1 i_0_0_803 (.A1(n_0_0_55), .A2(n_0_0_12), .ZN(n_0_139));
   NOR2_X1 i_0_0_804 (.A1(n_0_0_55), .A2(n_0_0_13), .ZN(n_0_140));
   NOR2_X1 i_0_0_805 (.A1(n_0_0_55), .A2(n_0_0_14), .ZN(n_0_141));
   NOR2_X1 i_0_0_806 (.A1(n_0_0_55), .A2(n_0_0_15), .ZN(n_0_142));
   NOR2_X1 i_0_0_807 (.A1(n_0_0_55), .A2(n_0_0_16), .ZN(n_0_143));
   NOR2_X1 i_0_0_808 (.A1(n_0_0_55), .A2(n_0_0_17), .ZN(n_0_144));
   NOR2_X1 i_0_0_809 (.A1(n_0_0_55), .A2(n_0_0_18), .ZN(n_0_145));
   NOR2_X1 i_0_0_810 (.A1(n_0_0_55), .A2(n_0_0_19), .ZN(n_0_146));
   NOR2_X1 i_0_0_811 (.A1(n_0_0_55), .A2(n_0_0_20), .ZN(n_0_147));
   NOR2_X1 i_0_0_812 (.A1(n_0_0_55), .A2(n_0_0_21), .ZN(n_0_148));
   NOR2_X1 i_0_0_813 (.A1(n_0_0_55), .A2(n_0_0_22), .ZN(n_0_149));
   NOR2_X1 i_0_0_814 (.A1(n_0_0_55), .A2(n_0_0_23), .ZN(n_0_150));
   NOR2_X1 i_0_0_815 (.A1(n_0_0_55), .A2(n_0_0_24), .ZN(n_0_151));
   NOR2_X1 i_0_0_816 (.A1(n_0_0_55), .A2(n_0_0_25), .ZN(n_0_152));
   NOR2_X1 i_0_0_817 (.A1(n_0_0_55), .A2(n_0_0_26), .ZN(n_0_153));
   NOR2_X1 i_0_0_818 (.A1(n_0_0_55), .A2(n_0_0_27), .ZN(n_0_154));
   NOR2_X1 i_0_0_819 (.A1(n_0_0_55), .A2(n_0_0_28), .ZN(n_0_155));
   NOR2_X1 i_0_0_820 (.A1(n_0_0_55), .A2(n_0_0_29), .ZN(n_0_156));
   NOR2_X1 i_0_0_821 (.A1(n_0_0_55), .A2(n_0_0_30), .ZN(n_0_157));
   NOR2_X1 i_0_0_822 (.A1(n_0_0_55), .A2(n_0_0_31), .ZN(n_0_158));
   NOR2_X1 i_0_0_823 (.A1(n_0_0_55), .A2(n_0_0_32), .ZN(n_0_159));
   INV_X1 i_0_0_824 (.A(b[24]), .ZN(n_0_0_56));
   NOR2_X1 i_0_0_825 (.A1(n_0_0_56), .A2(n_0_0_1), .ZN(n_0_96));
   NOR2_X1 i_0_0_826 (.A1(n_0_0_56), .A2(n_0_0_2), .ZN(n_0_97));
   NOR2_X1 i_0_0_827 (.A1(n_0_0_56), .A2(n_0_0_3), .ZN(n_0_98));
   NOR2_X1 i_0_0_828 (.A1(n_0_0_56), .A2(n_0_0_4), .ZN(n_0_99));
   NOR2_X1 i_0_0_829 (.A1(n_0_0_56), .A2(n_0_0_5), .ZN(n_0_100));
   NOR2_X1 i_0_0_830 (.A1(n_0_0_56), .A2(n_0_0_6), .ZN(n_0_101));
   NOR2_X1 i_0_0_831 (.A1(n_0_0_56), .A2(n_0_0_7), .ZN(n_0_102));
   NOR2_X1 i_0_0_832 (.A1(n_0_0_56), .A2(n_0_0_8), .ZN(n_0_103));
   NOR2_X1 i_0_0_833 (.A1(n_0_0_56), .A2(n_0_0_9), .ZN(n_0_104));
   NOR2_X1 i_0_0_834 (.A1(n_0_0_56), .A2(n_0_0_10), .ZN(n_0_105));
   NOR2_X1 i_0_0_835 (.A1(n_0_0_56), .A2(n_0_0_11), .ZN(n_0_106));
   NOR2_X1 i_0_0_836 (.A1(n_0_0_56), .A2(n_0_0_12), .ZN(n_0_107));
   NOR2_X1 i_0_0_837 (.A1(n_0_0_56), .A2(n_0_0_13), .ZN(n_0_108));
   NOR2_X1 i_0_0_838 (.A1(n_0_0_56), .A2(n_0_0_14), .ZN(n_0_109));
   NOR2_X1 i_0_0_839 (.A1(n_0_0_56), .A2(n_0_0_15), .ZN(n_0_110));
   NOR2_X1 i_0_0_840 (.A1(n_0_0_56), .A2(n_0_0_16), .ZN(n_0_111));
   NOR2_X1 i_0_0_841 (.A1(n_0_0_56), .A2(n_0_0_17), .ZN(n_0_112));
   NOR2_X1 i_0_0_842 (.A1(n_0_0_56), .A2(n_0_0_18), .ZN(n_0_113));
   NOR2_X1 i_0_0_843 (.A1(n_0_0_56), .A2(n_0_0_19), .ZN(n_0_114));
   NOR2_X1 i_0_0_844 (.A1(n_0_0_56), .A2(n_0_0_20), .ZN(n_0_115));
   NOR2_X1 i_0_0_845 (.A1(n_0_0_56), .A2(n_0_0_21), .ZN(n_0_116));
   NOR2_X1 i_0_0_846 (.A1(n_0_0_56), .A2(n_0_0_22), .ZN(n_0_117));
   NOR2_X1 i_0_0_847 (.A1(n_0_0_56), .A2(n_0_0_23), .ZN(n_0_118));
   NOR2_X1 i_0_0_848 (.A1(n_0_0_56), .A2(n_0_0_24), .ZN(n_0_119));
   NOR2_X1 i_0_0_849 (.A1(n_0_0_56), .A2(n_0_0_25), .ZN(n_0_120));
   NOR2_X1 i_0_0_850 (.A1(n_0_0_56), .A2(n_0_0_26), .ZN(n_0_121));
   NOR2_X1 i_0_0_851 (.A1(n_0_0_56), .A2(n_0_0_27), .ZN(n_0_122));
   NOR2_X1 i_0_0_852 (.A1(n_0_0_56), .A2(n_0_0_28), .ZN(n_0_123));
   NOR2_X1 i_0_0_853 (.A1(n_0_0_56), .A2(n_0_0_29), .ZN(n_0_124));
   NOR2_X1 i_0_0_854 (.A1(n_0_0_56), .A2(n_0_0_30), .ZN(n_0_125));
   NOR2_X1 i_0_0_855 (.A1(n_0_0_56), .A2(n_0_0_31), .ZN(n_0_126));
   NOR2_X1 i_0_0_856 (.A1(n_0_0_56), .A2(n_0_0_32), .ZN(n_0_127));
   INV_X1 i_0_0_857 (.A(b[25]), .ZN(n_0_0_57));
   NOR2_X1 i_0_0_858 (.A1(n_0_0_57), .A2(n_0_0_1), .ZN(n_0_64));
   NOR2_X1 i_0_0_859 (.A1(n_0_0_57), .A2(n_0_0_2), .ZN(n_0_65));
   NOR2_X1 i_0_0_860 (.A1(n_0_0_57), .A2(n_0_0_3), .ZN(n_0_66));
   NOR2_X1 i_0_0_861 (.A1(n_0_0_57), .A2(n_0_0_4), .ZN(n_0_67));
   NOR2_X1 i_0_0_862 (.A1(n_0_0_57), .A2(n_0_0_5), .ZN(n_0_68));
   NOR2_X1 i_0_0_863 (.A1(n_0_0_57), .A2(n_0_0_6), .ZN(n_0_69));
   NOR2_X1 i_0_0_864 (.A1(n_0_0_57), .A2(n_0_0_7), .ZN(n_0_70));
   NOR2_X1 i_0_0_865 (.A1(n_0_0_57), .A2(n_0_0_8), .ZN(n_0_71));
   NOR2_X1 i_0_0_866 (.A1(n_0_0_57), .A2(n_0_0_9), .ZN(n_0_72));
   NOR2_X1 i_0_0_867 (.A1(n_0_0_57), .A2(n_0_0_10), .ZN(n_0_73));
   NOR2_X1 i_0_0_868 (.A1(n_0_0_57), .A2(n_0_0_11), .ZN(n_0_74));
   NOR2_X1 i_0_0_869 (.A1(n_0_0_57), .A2(n_0_0_12), .ZN(n_0_75));
   NOR2_X1 i_0_0_870 (.A1(n_0_0_57), .A2(n_0_0_13), .ZN(n_0_76));
   NOR2_X1 i_0_0_871 (.A1(n_0_0_57), .A2(n_0_0_14), .ZN(n_0_77));
   NOR2_X1 i_0_0_872 (.A1(n_0_0_57), .A2(n_0_0_15), .ZN(n_0_78));
   NOR2_X1 i_0_0_873 (.A1(n_0_0_57), .A2(n_0_0_16), .ZN(n_0_79));
   NOR2_X1 i_0_0_874 (.A1(n_0_0_57), .A2(n_0_0_17), .ZN(n_0_80));
   NOR2_X1 i_0_0_875 (.A1(n_0_0_57), .A2(n_0_0_18), .ZN(n_0_81));
   NOR2_X1 i_0_0_876 (.A1(n_0_0_57), .A2(n_0_0_19), .ZN(n_0_82));
   NOR2_X1 i_0_0_877 (.A1(n_0_0_57), .A2(n_0_0_20), .ZN(n_0_83));
   NOR2_X1 i_0_0_878 (.A1(n_0_0_57), .A2(n_0_0_21), .ZN(n_0_84));
   NOR2_X1 i_0_0_879 (.A1(n_0_0_57), .A2(n_0_0_22), .ZN(n_0_85));
   NOR2_X1 i_0_0_880 (.A1(n_0_0_57), .A2(n_0_0_23), .ZN(n_0_86));
   NOR2_X1 i_0_0_881 (.A1(n_0_0_57), .A2(n_0_0_24), .ZN(n_0_87));
   NOR2_X1 i_0_0_882 (.A1(n_0_0_57), .A2(n_0_0_25), .ZN(n_0_88));
   NOR2_X1 i_0_0_883 (.A1(n_0_0_57), .A2(n_0_0_26), .ZN(n_0_89));
   NOR2_X1 i_0_0_884 (.A1(n_0_0_57), .A2(n_0_0_27), .ZN(n_0_90));
   NOR2_X1 i_0_0_885 (.A1(n_0_0_57), .A2(n_0_0_28), .ZN(n_0_91));
   NOR2_X1 i_0_0_886 (.A1(n_0_0_57), .A2(n_0_0_29), .ZN(n_0_92));
   NOR2_X1 i_0_0_887 (.A1(n_0_0_57), .A2(n_0_0_30), .ZN(n_0_93));
   NOR2_X1 i_0_0_888 (.A1(n_0_0_57), .A2(n_0_0_31), .ZN(n_0_94));
   NOR2_X1 i_0_0_889 (.A1(n_0_0_57), .A2(n_0_0_32), .ZN(n_0_95));
   INV_X1 i_0_0_890 (.A(b[26]), .ZN(n_0_0_58));
   NOR2_X1 i_0_0_891 (.A1(n_0_0_58), .A2(n_0_0_1), .ZN(n_0_33));
   NOR2_X1 i_0_0_892 (.A1(n_0_0_58), .A2(n_0_0_2), .ZN(n_0_34));
   NOR2_X1 i_0_0_893 (.A1(n_0_0_58), .A2(n_0_0_3), .ZN(n_0_35));
   NOR2_X1 i_0_0_894 (.A1(n_0_0_58), .A2(n_0_0_4), .ZN(n_0_36));
   NOR2_X1 i_0_0_895 (.A1(n_0_0_58), .A2(n_0_0_5), .ZN(n_0_37));
   NOR2_X1 i_0_0_896 (.A1(n_0_0_58), .A2(n_0_0_6), .ZN(n_0_38));
   NOR2_X1 i_0_0_897 (.A1(n_0_0_58), .A2(n_0_0_7), .ZN(n_0_39));
   NOR2_X1 i_0_0_898 (.A1(n_0_0_58), .A2(n_0_0_8), .ZN(n_0_40));
   NOR2_X1 i_0_0_899 (.A1(n_0_0_58), .A2(n_0_0_9), .ZN(n_0_41));
   NOR2_X1 i_0_0_900 (.A1(n_0_0_58), .A2(n_0_0_10), .ZN(n_0_42));
   NOR2_X1 i_0_0_901 (.A1(n_0_0_58), .A2(n_0_0_11), .ZN(n_0_43));
   NOR2_X1 i_0_0_902 (.A1(n_0_0_58), .A2(n_0_0_12), .ZN(n_0_44));
   NOR2_X1 i_0_0_903 (.A1(n_0_0_58), .A2(n_0_0_13), .ZN(n_0_45));
   NOR2_X1 i_0_0_904 (.A1(n_0_0_58), .A2(n_0_0_14), .ZN(n_0_46));
   NOR2_X1 i_0_0_905 (.A1(n_0_0_58), .A2(n_0_0_15), .ZN(n_0_47));
   NOR2_X1 i_0_0_906 (.A1(n_0_0_58), .A2(n_0_0_16), .ZN(n_0_48));
   NOR2_X1 i_0_0_907 (.A1(n_0_0_58), .A2(n_0_0_17), .ZN(n_0_49));
   NOR2_X1 i_0_0_908 (.A1(n_0_0_58), .A2(n_0_0_18), .ZN(n_0_50));
   NOR2_X1 i_0_0_909 (.A1(n_0_0_58), .A2(n_0_0_19), .ZN(n_0_51));
   NOR2_X1 i_0_0_910 (.A1(n_0_0_58), .A2(n_0_0_20), .ZN(n_0_52));
   NOR2_X1 i_0_0_911 (.A1(n_0_0_58), .A2(n_0_0_21), .ZN(n_0_53));
   NOR2_X1 i_0_0_912 (.A1(n_0_0_58), .A2(n_0_0_22), .ZN(n_0_54));
   NOR2_X1 i_0_0_913 (.A1(n_0_0_58), .A2(n_0_0_23), .ZN(n_0_55));
   NOR2_X1 i_0_0_914 (.A1(n_0_0_58), .A2(n_0_0_24), .ZN(n_0_56));
   NOR2_X1 i_0_0_915 (.A1(n_0_0_58), .A2(n_0_0_25), .ZN(n_0_57));
   NOR2_X1 i_0_0_916 (.A1(n_0_0_58), .A2(n_0_0_26), .ZN(n_0_58));
   NOR2_X1 i_0_0_917 (.A1(n_0_0_58), .A2(n_0_0_27), .ZN(n_0_59));
   NOR2_X1 i_0_0_918 (.A1(n_0_0_58), .A2(n_0_0_28), .ZN(n_0_60));
   NOR2_X1 i_0_0_919 (.A1(n_0_0_58), .A2(n_0_0_29), .ZN(n_0_61));
   NOR2_X1 i_0_0_920 (.A1(n_0_0_58), .A2(n_0_0_30), .ZN(n_0_62));
   NOR2_X1 i_0_0_921 (.A1(n_0_0_58), .A2(n_0_0_31), .ZN(n_0_63));
   NOR2_X1 i_0_0_922 (.A1(n_0_0_58), .A2(n_0_0_32), .ZN(n_0_192));
   INV_X1 i_0_0_923 (.A(b[27]), .ZN(n_0_0_59));
   NOR2_X1 i_0_0_924 (.A1(n_0_0_59), .A2(n_0_0_1), .ZN(n_287));
   NOR2_X1 i_0_0_925 (.A1(n_0_0_59), .A2(n_0_0_2), .ZN(n_288));
   NOR2_X1 i_0_0_926 (.A1(n_0_0_59), .A2(n_0_0_3), .ZN(n_289));
   NOR2_X1 i_0_0_927 (.A1(n_0_0_59), .A2(n_0_0_4), .ZN(n_290));
   NOR2_X1 i_0_0_928 (.A1(n_0_0_59), .A2(n_0_0_5), .ZN(n_291));
   NOR2_X1 i_0_0_929 (.A1(n_0_0_59), .A2(n_0_0_6), .ZN(n_292));
   NOR2_X1 i_0_0_930 (.A1(n_0_0_59), .A2(n_0_0_7), .ZN(n_293));
   NOR2_X1 i_0_0_931 (.A1(n_0_0_59), .A2(n_0_0_8), .ZN(n_294));
   NOR2_X1 i_0_0_932 (.A1(n_0_0_59), .A2(n_0_0_9), .ZN(n_295));
   NOR2_X1 i_0_0_933 (.A1(n_0_0_59), .A2(n_0_0_10), .ZN(n_296));
   NOR2_X1 i_0_0_934 (.A1(n_0_0_59), .A2(n_0_0_11), .ZN(n_297));
   NOR2_X1 i_0_0_935 (.A1(n_0_0_59), .A2(n_0_0_12), .ZN(n_298));
   NOR2_X1 i_0_0_936 (.A1(n_0_0_59), .A2(n_0_0_13), .ZN(n_299));
   NOR2_X1 i_0_0_937 (.A1(n_0_0_59), .A2(n_0_0_14), .ZN(n_300));
   NOR2_X1 i_0_0_938 (.A1(n_0_0_59), .A2(n_0_0_15), .ZN(n_301));
   NOR2_X1 i_0_0_939 (.A1(n_0_0_59), .A2(n_0_0_16), .ZN(n_302));
   NOR2_X1 i_0_0_940 (.A1(n_0_0_59), .A2(n_0_0_17), .ZN(n_303));
   NOR2_X1 i_0_0_941 (.A1(n_0_0_59), .A2(n_0_0_18), .ZN(n_304));
   NOR2_X1 i_0_0_942 (.A1(n_0_0_59), .A2(n_0_0_19), .ZN(n_305));
   NOR2_X1 i_0_0_943 (.A1(n_0_0_59), .A2(n_0_0_20), .ZN(n_306));
   NOR2_X1 i_0_0_944 (.A1(n_0_0_59), .A2(n_0_0_21), .ZN(n_307));
   NOR2_X1 i_0_0_945 (.A1(n_0_0_59), .A2(n_0_0_22), .ZN(n_308));
   NOR2_X1 i_0_0_946 (.A1(n_0_0_59), .A2(n_0_0_23), .ZN(n_309));
   NOR2_X1 i_0_0_947 (.A1(n_0_0_59), .A2(n_0_0_24), .ZN(n_310));
   NOR2_X1 i_0_0_948 (.A1(n_0_0_59), .A2(n_0_0_25), .ZN(n_311));
   NOR2_X1 i_0_0_949 (.A1(n_0_0_59), .A2(n_0_0_26), .ZN(n_312));
   NOR2_X1 i_0_0_950 (.A1(n_0_0_59), .A2(n_0_0_27), .ZN(n_313));
   NOR2_X1 i_0_0_951 (.A1(n_0_0_59), .A2(n_0_0_28), .ZN(n_314));
   NOR2_X1 i_0_0_952 (.A1(n_0_0_59), .A2(n_0_0_29), .ZN(n_315));
   NOR2_X1 i_0_0_953 (.A1(n_0_0_59), .A2(n_0_0_30), .ZN(n_316));
   NOR2_X1 i_0_0_954 (.A1(n_0_0_59), .A2(n_0_0_31), .ZN(n_317));
   NOR2_X1 i_0_0_955 (.A1(n_0_0_59), .A2(n_0_0_32), .ZN(n_318));
   INV_X1 i_0_0_956 (.A(b[28]), .ZN(n_0_0_60));
   NOR2_X1 i_0_0_957 (.A1(n_0_0_60), .A2(n_0_0_1), .ZN(n_319));
   NOR2_X1 i_0_0_958 (.A1(n_0_0_60), .A2(n_0_0_2), .ZN(n_320));
   NOR2_X1 i_0_0_959 (.A1(n_0_0_60), .A2(n_0_0_3), .ZN(n_321));
   NOR2_X1 i_0_0_960 (.A1(n_0_0_60), .A2(n_0_0_4), .ZN(n_322));
   NOR2_X1 i_0_0_961 (.A1(n_0_0_60), .A2(n_0_0_5), .ZN(n_323));
   NOR2_X1 i_0_0_962 (.A1(n_0_0_60), .A2(n_0_0_6), .ZN(n_324));
   NOR2_X1 i_0_0_963 (.A1(n_0_0_60), .A2(n_0_0_7), .ZN(n_325));
   NOR2_X1 i_0_0_964 (.A1(n_0_0_60), .A2(n_0_0_8), .ZN(n_326));
   NOR2_X1 i_0_0_965 (.A1(n_0_0_60), .A2(n_0_0_9), .ZN(n_327));
   NOR2_X1 i_0_0_966 (.A1(n_0_0_60), .A2(n_0_0_10), .ZN(n_328));
   NOR2_X1 i_0_0_967 (.A1(n_0_0_60), .A2(n_0_0_11), .ZN(n_329));
   NOR2_X1 i_0_0_968 (.A1(n_0_0_60), .A2(n_0_0_12), .ZN(n_330));
   NOR2_X1 i_0_0_969 (.A1(n_0_0_60), .A2(n_0_0_13), .ZN(n_331));
   NOR2_X1 i_0_0_970 (.A1(n_0_0_60), .A2(n_0_0_14), .ZN(n_332));
   NOR2_X1 i_0_0_971 (.A1(n_0_0_60), .A2(n_0_0_15), .ZN(n_333));
   NOR2_X1 i_0_0_972 (.A1(n_0_0_60), .A2(n_0_0_16), .ZN(n_334));
   NOR2_X1 i_0_0_973 (.A1(n_0_0_60), .A2(n_0_0_17), .ZN(n_335));
   NOR2_X1 i_0_0_974 (.A1(n_0_0_60), .A2(n_0_0_18), .ZN(n_336));
   NOR2_X1 i_0_0_975 (.A1(n_0_0_60), .A2(n_0_0_19), .ZN(n_337));
   NOR2_X1 i_0_0_976 (.A1(n_0_0_60), .A2(n_0_0_20), .ZN(n_338));
   NOR2_X1 i_0_0_977 (.A1(n_0_0_60), .A2(n_0_0_21), .ZN(n_339));
   NOR2_X1 i_0_0_978 (.A1(n_0_0_60), .A2(n_0_0_22), .ZN(n_340));
   NOR2_X1 i_0_0_979 (.A1(n_0_0_60), .A2(n_0_0_23), .ZN(n_341));
   NOR2_X1 i_0_0_980 (.A1(n_0_0_60), .A2(n_0_0_24), .ZN(n_342));
   NOR2_X1 i_0_0_981 (.A1(n_0_0_60), .A2(n_0_0_25), .ZN(n_343));
   NOR2_X1 i_0_0_982 (.A1(n_0_0_60), .A2(n_0_0_26), .ZN(n_344));
   NOR2_X1 i_0_0_983 (.A1(n_0_0_60), .A2(n_0_0_27), .ZN(n_345));
   NOR2_X1 i_0_0_984 (.A1(n_0_0_60), .A2(n_0_0_28), .ZN(n_346));
   NOR2_X1 i_0_0_985 (.A1(n_0_0_60), .A2(n_0_0_29), .ZN(n_347));
   NOR2_X1 i_0_0_986 (.A1(n_0_0_60), .A2(n_0_0_30), .ZN(n_348));
   NOR2_X1 i_0_0_987 (.A1(n_0_0_60), .A2(n_0_0_31), .ZN(n_349));
   NOR2_X1 i_0_0_988 (.A1(n_0_0_60), .A2(n_0_0_32), .ZN(n_350));
   INV_X1 i_0_0_989 (.A(b[29]), .ZN(n_0_0_61));
   NOR2_X1 i_0_0_990 (.A1(n_0_0_61), .A2(n_0_0_1), .ZN(n_351));
   NOR2_X1 i_0_0_991 (.A1(n_0_0_61), .A2(n_0_0_2), .ZN(n_352));
   NOR2_X1 i_0_0_992 (.A1(n_0_0_61), .A2(n_0_0_3), .ZN(n_353));
   NOR2_X1 i_0_0_993 (.A1(n_0_0_61), .A2(n_0_0_4), .ZN(n_354));
   NOR2_X1 i_0_0_994 (.A1(n_0_0_61), .A2(n_0_0_5), .ZN(n_355));
   NOR2_X1 i_0_0_995 (.A1(n_0_0_61), .A2(n_0_0_6), .ZN(n_356));
   NOR2_X1 i_0_0_996 (.A1(n_0_0_61), .A2(n_0_0_7), .ZN(n_357));
   NOR2_X1 i_0_0_997 (.A1(n_0_0_61), .A2(n_0_0_8), .ZN(n_358));
   NOR2_X1 i_0_0_998 (.A1(n_0_0_61), .A2(n_0_0_9), .ZN(n_359));
   NOR2_X1 i_0_0_999 (.A1(n_0_0_61), .A2(n_0_0_10), .ZN(n_360));
   NOR2_X1 i_0_0_1000 (.A1(n_0_0_61), .A2(n_0_0_11), .ZN(n_361));
   NOR2_X1 i_0_0_1001 (.A1(n_0_0_61), .A2(n_0_0_12), .ZN(n_362));
   NOR2_X1 i_0_0_1002 (.A1(n_0_0_61), .A2(n_0_0_13), .ZN(n_363));
   NOR2_X1 i_0_0_1003 (.A1(n_0_0_61), .A2(n_0_0_14), .ZN(n_364));
   NOR2_X1 i_0_0_1004 (.A1(n_0_0_61), .A2(n_0_0_15), .ZN(n_365));
   NOR2_X1 i_0_0_1005 (.A1(n_0_0_61), .A2(n_0_0_16), .ZN(n_366));
   NOR2_X1 i_0_0_1006 (.A1(n_0_0_61), .A2(n_0_0_17), .ZN(n_367));
   NOR2_X1 i_0_0_1007 (.A1(n_0_0_61), .A2(n_0_0_18), .ZN(n_368));
   NOR2_X1 i_0_0_1008 (.A1(n_0_0_61), .A2(n_0_0_19), .ZN(n_369));
   NOR2_X1 i_0_0_1009 (.A1(n_0_0_61), .A2(n_0_0_20), .ZN(n_370));
   NOR2_X1 i_0_0_1010 (.A1(n_0_0_61), .A2(n_0_0_21), .ZN(n_371));
   NOR2_X1 i_0_0_1011 (.A1(n_0_0_61), .A2(n_0_0_22), .ZN(n_372));
   NOR2_X1 i_0_0_1012 (.A1(n_0_0_61), .A2(n_0_0_23), .ZN(n_373));
   NOR2_X1 i_0_0_1013 (.A1(n_0_0_61), .A2(n_0_0_24), .ZN(n_374));
   NOR2_X1 i_0_0_1014 (.A1(n_0_0_61), .A2(n_0_0_25), .ZN(n_375));
   NOR2_X1 i_0_0_1015 (.A1(n_0_0_61), .A2(n_0_0_26), .ZN(n_376));
   NOR2_X1 i_0_0_1016 (.A1(n_0_0_61), .A2(n_0_0_27), .ZN(n_377));
   NOR2_X1 i_0_0_1017 (.A1(n_0_0_61), .A2(n_0_0_28), .ZN(n_378));
   NOR2_X1 i_0_0_1018 (.A1(n_0_0_61), .A2(n_0_0_29), .ZN(n_379));
   NOR2_X1 i_0_0_1019 (.A1(n_0_0_61), .A2(n_0_0_30), .ZN(n_380));
   NOR2_X1 i_0_0_1020 (.A1(n_0_0_61), .A2(n_0_0_31), .ZN(n_381));
   NOR2_X1 i_0_0_1021 (.A1(n_0_0_61), .A2(n_0_0_32), .ZN(n_382));
   INV_X1 i_0_0_1022 (.A(b[30]), .ZN(n_0_0_62));
   NOR2_X1 i_0_0_1023 (.A1(n_0_0_62), .A2(n_0_0_1), .ZN(n_383));
   NOR2_X1 i_0_0_1024 (.A1(n_0_0_62), .A2(n_0_0_2), .ZN(n_384));
   NOR2_X1 i_0_0_1025 (.A1(n_0_0_62), .A2(n_0_0_3), .ZN(n_385));
   NOR2_X1 i_0_0_1026 (.A1(n_0_0_62), .A2(n_0_0_4), .ZN(n_386));
   NOR2_X1 i_0_0_1027 (.A1(n_0_0_62), .A2(n_0_0_5), .ZN(n_387));
   NOR2_X1 i_0_0_1028 (.A1(n_0_0_62), .A2(n_0_0_6), .ZN(n_388));
   NOR2_X1 i_0_0_1029 (.A1(n_0_0_62), .A2(n_0_0_7), .ZN(n_389));
   NOR2_X1 i_0_0_1030 (.A1(n_0_0_62), .A2(n_0_0_8), .ZN(n_390));
   NOR2_X1 i_0_0_1031 (.A1(n_0_0_62), .A2(n_0_0_9), .ZN(n_391));
   NOR2_X1 i_0_0_1032 (.A1(n_0_0_62), .A2(n_0_0_10), .ZN(n_392));
   NOR2_X1 i_0_0_1033 (.A1(n_0_0_62), .A2(n_0_0_11), .ZN(n_393));
   NOR2_X1 i_0_0_1034 (.A1(n_0_0_62), .A2(n_0_0_12), .ZN(n_394));
   NOR2_X1 i_0_0_1035 (.A1(n_0_0_62), .A2(n_0_0_13), .ZN(n_395));
   NOR2_X1 i_0_0_1036 (.A1(n_0_0_62), .A2(n_0_0_14), .ZN(n_396));
   NOR2_X1 i_0_0_1037 (.A1(n_0_0_62), .A2(n_0_0_15), .ZN(n_397));
   NOR2_X1 i_0_0_1038 (.A1(n_0_0_62), .A2(n_0_0_16), .ZN(n_398));
   NOR2_X1 i_0_0_1039 (.A1(n_0_0_62), .A2(n_0_0_17), .ZN(n_399));
   NOR2_X1 i_0_0_1040 (.A1(n_0_0_62), .A2(n_0_0_18), .ZN(n_400));
   NOR2_X1 i_0_0_1041 (.A1(n_0_0_62), .A2(n_0_0_19), .ZN(n_401));
   NOR2_X1 i_0_0_1042 (.A1(n_0_0_62), .A2(n_0_0_20), .ZN(n_402));
   NOR2_X1 i_0_0_1043 (.A1(n_0_0_62), .A2(n_0_0_21), .ZN(n_403));
   NOR2_X1 i_0_0_1044 (.A1(n_0_0_62), .A2(n_0_0_22), .ZN(n_404));
   NOR2_X1 i_0_0_1045 (.A1(n_0_0_62), .A2(n_0_0_23), .ZN(n_405));
   NOR2_X1 i_0_0_1046 (.A1(n_0_0_62), .A2(n_0_0_24), .ZN(n_406));
   NOR2_X1 i_0_0_1047 (.A1(n_0_0_62), .A2(n_0_0_25), .ZN(n_407));
   NOR2_X1 i_0_0_1048 (.A1(n_0_0_62), .A2(n_0_0_26), .ZN(n_408));
   NOR2_X1 i_0_0_1049 (.A1(n_0_0_62), .A2(n_0_0_27), .ZN(n_409));
   NOR2_X1 i_0_0_1050 (.A1(n_0_0_62), .A2(n_0_0_28), .ZN(n_410));
   NOR2_X1 i_0_0_1051 (.A1(n_0_0_62), .A2(n_0_0_29), .ZN(n_411));
   NOR2_X1 i_0_0_1052 (.A1(n_0_0_62), .A2(n_0_0_30), .ZN(n_412));
   NOR2_X1 i_0_0_1053 (.A1(n_0_0_62), .A2(n_0_0_31), .ZN(n_413));
   NOR2_X1 i_0_0_1054 (.A1(n_0_0_62), .A2(n_0_0_32), .ZN(n_414));
   INV_X1 i_0_0_1055 (.A(b[31]), .ZN(n_0_0_63));
   NOR2_X1 i_0_0_1056 (.A1(n_0_0_63), .A2(a[0]), .ZN(n_415));
   NOR2_X1 i_0_0_1057 (.A1(n_0_0_63), .A2(a[1]), .ZN(n_416));
   NOR2_X1 i_0_0_1058 (.A1(n_0_0_63), .A2(a[2]), .ZN(n_417));
   NOR2_X1 i_0_0_1059 (.A1(n_0_0_63), .A2(a[3]), .ZN(n_418));
   NOR2_X1 i_0_0_1060 (.A1(n_0_0_63), .A2(a[4]), .ZN(n_419));
   NOR2_X1 i_0_0_1061 (.A1(n_0_0_63), .A2(a[5]), .ZN(n_420));
   NOR2_X1 i_0_0_1062 (.A1(n_0_0_63), .A2(a[6]), .ZN(n_421));
   NOR2_X1 i_0_0_1063 (.A1(n_0_0_63), .A2(a[7]), .ZN(n_422));
   NOR2_X1 i_0_0_1064 (.A1(n_0_0_63), .A2(a[8]), .ZN(n_423));
   NOR2_X1 i_0_0_1065 (.A1(n_0_0_63), .A2(a[9]), .ZN(n_424));
   NOR2_X1 i_0_0_1066 (.A1(n_0_0_63), .A2(a[10]), .ZN(n_425));
   NOR2_X1 i_0_0_1067 (.A1(n_0_0_63), .A2(a[11]), .ZN(n_426));
   NOR2_X1 i_0_0_1068 (.A1(n_0_0_63), .A2(a[12]), .ZN(n_427));
   NOR2_X1 i_0_0_1069 (.A1(n_0_0_63), .A2(a[13]), .ZN(n_428));
   NOR2_X1 i_0_0_1070 (.A1(n_0_0_63), .A2(a[14]), .ZN(n_429));
   NOR2_X1 i_0_0_1071 (.A1(n_0_0_63), .A2(a[15]), .ZN(n_430));
   NOR2_X1 i_0_0_1072 (.A1(n_0_0_63), .A2(a[16]), .ZN(n_431));
   NOR2_X1 i_0_0_1073 (.A1(n_0_0_63), .A2(a[17]), .ZN(n_432));
   NOR2_X1 i_0_0_1074 (.A1(n_0_0_63), .A2(a[18]), .ZN(n_433));
   NOR2_X1 i_0_0_1075 (.A1(n_0_0_63), .A2(a[19]), .ZN(n_434));
   NOR2_X1 i_0_0_1076 (.A1(n_0_0_63), .A2(a[20]), .ZN(n_435));
   NOR2_X1 i_0_0_1077 (.A1(n_0_0_63), .A2(a[21]), .ZN(n_436));
   NOR2_X1 i_0_0_1078 (.A1(n_0_0_63), .A2(a[22]), .ZN(n_437));
   NOR2_X1 i_0_0_1079 (.A1(n_0_0_63), .A2(a[23]), .ZN(n_438));
   NOR2_X1 i_0_0_1080 (.A1(n_0_0_63), .A2(a[24]), .ZN(n_439));
   NOR2_X1 i_0_0_1081 (.A1(n_0_0_63), .A2(a[25]), .ZN(n_440));
   NOR2_X1 i_0_0_1082 (.A1(n_0_0_63), .A2(a[26]), .ZN(n_441));
   NOR2_X1 i_0_0_1083 (.A1(n_0_0_63), .A2(a[27]), .ZN(n_442));
   NOR2_X1 i_0_0_1084 (.A1(n_0_0_63), .A2(a[28]), .ZN(n_443));
   NOR2_X1 i_0_0_1085 (.A1(n_0_0_63), .A2(a[29]), .ZN(n_444));
   NOR2_X1 i_0_0_1086 (.A1(n_0_0_63), .A2(a[30]), .ZN(n_445));
   NOR2_X1 i_0_0_1087 (.A1(n_0_0_63), .A2(a[31]), .ZN(n_446));
   INV_X1 i_0_0_0 (.A(b[1]), .ZN(n_0_0_33));
   INV_X1 i_0_0_63 (.A(a[31]), .ZN(n_0_0_32));
   INV_X1 i_0_0_64 (.A(b[0]), .ZN(n_0_0_0));
   INV_X1 i_0_0_65 (.A(n_0_0_64), .ZN(n_0_30));
   NAND2_X1 i_0_0_97 (.A1(a[31]), .A2(b[0]), .ZN(n_0_0_64));
   INV_X1 i_0_0_1088 (.A(n_0_0_65), .ZN(n_0_32));
   NAND2_X1 i_0_0_1089 (.A1(a[31]), .A2(b[1]), .ZN(n_0_0_65));
   CSA__2_2 A2_4 (.in1({\c1[4] [46], uc_2097, uc_2098, uc_2099, uc_2100, uc_2101, 
      uc_2102, uc_2103, uc_2104, uc_2105, uc_2106, uc_2107, uc_2108, uc_2109, 
      uc_2110, uc_2111, uc_2112, uc_2113, \c1[4] [45], \c1[4] [44], \c1[4] [43], 
      \c1[4] [42], \c1[4] [41], \c1[4] [40], \c1[4] [39], \c1[4] [38], 
      \c1[4] [37], \c1[4] [36], \c1[4] [35], \c1[4] [34], \c1[4] [33], 
      \c1[4] [32], \c1[4] [31], \c1[4] [30], \c1[4] [29], \c1[4] [28], 
      \c1[4] [27], \c1[4] [26], \c1[4] [25], \c1[4] [24], \c1[4] [23], 
      \c1[4] [22], \c1[4] [21], \c1[4] [20], \c1[4] [19], \c1[4] [18], 
      \c1[4] [17], \c1[4] [16], \c1[4] [15], uc_2114, uc_2115, uc_2116, uc_2117, 
      uc_2118, uc_2119, uc_2120, uc_2121, uc_2122, uc_2123, uc_2124, uc_2125, 
      uc_2126, uc_2127, uc_2128}), .in2({\s1[5] [48], uc_2129, uc_2130, uc_2131, 
      uc_2132, uc_2133, uc_2134, uc_2135, uc_2136, uc_2137, uc_2138, uc_2139, 
      uc_2140, uc_2141, uc_2142, uc_2143, \s1[5] [47], \s1[5] [46], \s1[5] [45], 
      \s1[5] [44], \s1[5] [43], \s1[5] [42], \s1[5] [41], \s1[5] [40], 
      \s1[5] [39], \s1[5] [38], \s1[5] [37], \s1[5] [36], \s1[5] [35], 
      \s1[5] [34], \s1[5] [33], \s1[5] [32], \s1[5] [31], \s1[5] [30], 
      \s1[5] [29], \s1[5] [28], \s1[5] [27], \s1[5] [26], \s1[5] [25], 
      \s1[5] [24], \s1[5] [23], \s1[5] [22], \s1[5] [21], \s1[5] [20], 
      \s1[5] [19], \s1[5] [18], \s1[5] [17], \s1[5] [16], n_95, uc_2144, uc_2145, 
      uc_2146, uc_2147, uc_2148, uc_2149, uc_2150, uc_2151, uc_2152, uc_2153, 
      uc_2154, uc_2155, uc_2156, uc_2157, uc_2158}), .in3({\c1[5] [49], uc_2159, 
      uc_2160, uc_2161, uc_2162, uc_2163, uc_2164, uc_2165, uc_2166, uc_2167, 
      uc_2168, uc_2169, uc_2170, uc_2171, uc_2172, \c1[5] [48], \c1[5] [47], 
      \c1[5] [46], \c1[5] [45], \c1[5] [44], \c1[5] [43], \c1[5] [42], 
      \c1[5] [41], \c1[5] [40], \c1[5] [39], \c1[5] [38], \c1[5] [37], 
      \c1[5] [36], \c1[5] [35], \c1[5] [34], \c1[5] [33], \c1[5] [32], 
      \c1[5] [31], \c1[5] [30], \c1[5] [29], \c1[5] [28], \c1[5] [27], 
      \c1[5] [26], \c1[5] [25], \c1[5] [24], \c1[5] [23], \c1[5] [22], 
      \c1[5] [21], \c1[5] [20], \c1[5] [19], \c1[5] [18], \c1[5] [17], uc_2173, 
      uc_2174, uc_2175, uc_2176, uc_2177, uc_2178, uc_2179, uc_2180, uc_2181, 
      uc_2182, uc_2183, uc_2184, uc_2185, uc_2186, uc_2187, uc_2188, uc_2189}), 
      .sum({\s2[3] [49], uc_2190, uc_2191, uc_2192, uc_2193, uc_2194, uc_2195, 
      uc_2196, uc_2197, uc_2198, uc_2199, uc_2200, uc_2201, uc_2202, uc_2203, 
      \s2[3] [48], \s2[3] [47], \s2[3] [46], \s2[3] [45], \s2[3] [44], 
      \s2[3] [43], \s2[3] [42], \s2[3] [41], \s2[3] [40], \s2[3] [39], 
      \s2[3] [38], \s2[3] [37], \s2[3] [36], \s2[3] [35], \s2[3] [34], 
      \s2[3] [33], \s2[3] [32], \s2[3] [31], \s2[3] [30], \s2[3] [29], 
      \s2[3] [28], \s2[3] [27], \s2[3] [26], \s2[3] [25], \s2[3] [24], 
      \s2[3] [23], \s2[3] [22], \s2[3] [21], \s2[3] [20], \s2[3] [19], 
      \s2[3] [18], \s2[3] [17], \s2[3] [16], \s2[3] [15], uc_2204, uc_2205, 
      uc_2206, uc_2207, uc_2208, uc_2209, uc_2210, uc_2211, uc_2212, uc_2213, 
      uc_2214, uc_2215, uc_2216, uc_2217, uc_2218}), .c({\c2[3] [50], uc_2219, 
      uc_2220, uc_2221, uc_2222, uc_2223, uc_2224, uc_2225, uc_2226, uc_2227, 
      uc_2228, uc_2229, uc_2230, uc_2231, \c2[3] [49], \c2[3] [48], \c2[3] [47], 
      \c2[3] [46], \c2[3] [45], \c2[3] [44], \c2[3] [43], \c2[3] [42], 
      \c2[3] [41], \c2[3] [40], \c2[3] [39], \c2[3] [38], \c2[3] [37], 
      \c2[3] [36], \c2[3] [35], \c2[3] [34], \c2[3] [33], \c2[3] [32], 
      \c2[3] [31], \c2[3] [30], \c2[3] [29], \c2[3] [28], \c2[3] [27], 
      \c2[3] [26], \c2[3] [25], \c2[3] [24], \c2[3] [23], \c2[3] [22], 
      \c2[3] [21], \c2[3] [20], \c2[3] [19], \c2[3] [18], \c2[3] [17], 
      \c2[3] [16], uc_2232, uc_2233, uc_2234, uc_2235, uc_2236, uc_2237, uc_2238, 
      uc_2239, uc_2240, uc_2241, uc_2242, uc_2243, uc_2244, uc_2245, uc_2246, 
      uc_2247}));
   CSA__2_5 A1_6 (.in1({n_126, uc_2248, uc_2249, uc_2250, uc_2251, uc_2252, 
      uc_2253, uc_2254, uc_2255, uc_2256, uc_2257, uc_2258, uc_2259, uc_2260, 
      uc_2261, uc_2262, uc_2263, uc_2264, n_125, n_124, n_123, n_122, n_121, 
      n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, 
      n_110, n_109, n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, 
      n_100, n_99, n_98, n_97, n_96, uc_2265, uc_2266, uc_2267, uc_2268, uc_2269, 
      uc_2270, uc_2271, uc_2272, uc_2273, uc_2274, uc_2275, uc_2276, uc_2277, 
      uc_2278, uc_2279, uc_2280}), .in2({n_158, uc_2281, uc_2282, uc_2283, 
      uc_2284, uc_2285, uc_2286, uc_2287, uc_2288, uc_2289, uc_2290, uc_2291, 
      uc_2292, uc_2293, uc_2294, uc_2295, uc_2296, n_157, n_156, n_155, n_154, 
      n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, 
      n_143, n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, 
      n_133, n_132, n_131, n_130, n_129, n_128, n_127, uc_2297, uc_2298, uc_2299, 
      uc_2300, uc_2301, uc_2302, uc_2303, uc_2304, uc_2305, uc_2306, uc_2307, 
      uc_2308, uc_2309, uc_2310, uc_2311, uc_2312}), .in3({n_190, uc_2313, 
      uc_2314, uc_2315, uc_2316, uc_2317, uc_2318, uc_2319, uc_2320, uc_2321, 
      uc_2322, uc_2323, uc_2324, uc_2325, uc_2326, uc_2327, n_189, n_188, n_187, 
      n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_178, n_177, 
      n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, 
      n_166, n_165, n_164, n_163, n_162, n_161, n_160, n_159, uc_2328, uc_2329, 
      uc_2330, uc_2331, uc_2332, uc_2333, uc_2334, uc_2335, uc_2336, uc_2337, 
      uc_2338, uc_2339, uc_2340, uc_2341, uc_2342, uc_2343, uc_2344}), .sum({
      \s1[5] [48], uc_2345, uc_2346, uc_2347, uc_2348, uc_2349, uc_2350, uc_2351, 
      uc_2352, uc_2353, uc_2354, uc_2355, uc_2356, uc_2357, uc_2358, uc_2359, 
      \s1[5] [47], \s1[5] [46], \s1[5] [45], \s1[5] [44], \s1[5] [43], 
      \s1[5] [42], \s1[5] [41], \s1[5] [40], \s1[5] [39], \s1[5] [38], 
      \s1[5] [37], \s1[5] [36], \s1[5] [35], \s1[5] [34], \s1[5] [33], 
      \s1[5] [32], \s1[5] [31], \s1[5] [30], \s1[5] [29], \s1[5] [28], 
      \s1[5] [27], \s1[5] [26], \s1[5] [25], \s1[5] [24], \s1[5] [23], 
      \s1[5] [22], \s1[5] [21], \s1[5] [20], \s1[5] [19], \s1[5] [18], 
      \s1[5] [17], \s1[5] [16], uc_2360, uc_2361, uc_2362, uc_2363, uc_2364, 
      uc_2365, uc_2366, uc_2367, uc_2368, uc_2369, uc_2370, uc_2371, uc_2372, 
      uc_2373, uc_2374, uc_2375}), .c({\c1[5] [49], uc_2376, uc_2377, uc_2378, 
      uc_2379, uc_2380, uc_2381, uc_2382, uc_2383, uc_2384, uc_2385, uc_2386, 
      uc_2387, uc_2388, uc_2389, \c1[5] [48], \c1[5] [47], \c1[5] [46], 
      \c1[5] [45], \c1[5] [44], \c1[5] [43], \c1[5] [42], \c1[5] [41], 
      \c1[5] [40], \c1[5] [39], \c1[5] [38], \c1[5] [37], \c1[5] [36], 
      \c1[5] [35], \c1[5] [34], \c1[5] [33], \c1[5] [32], \c1[5] [31], 
      \c1[5] [30], \c1[5] [29], \c1[5] [28], \c1[5] [27], \c1[5] [26], 
      \c1[5] [25], \c1[5] [24], \c1[5] [23], \c1[5] [22], \c1[5] [21], 
      \c1[5] [20], \c1[5] [19], \c1[5] [18], \c1[5] [17], uc_2390, uc_2391, 
      uc_2392, uc_2393, uc_2394, uc_2395, uc_2396, uc_2397, uc_2398, uc_2399, 
      uc_2400, uc_2401, uc_2402, uc_2403, uc_2404, uc_2405, uc_2406}));
   CSA__0_71 A1_5 (.in1({n_30, uc_2407, uc_2408, uc_2409, uc_2410, uc_2411, 
      uc_2412, uc_2413, uc_2414, uc_2415, uc_2416, uc_2417, uc_2418, uc_2419, 
      uc_2420, uc_2421, uc_2422, uc_2423, uc_2424, uc_2425, uc_2426, n_29, n_28, 
      n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, 
      n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, 
      n_1, n_0, uc_2427, uc_2428, uc_2429, uc_2430, uc_2431, uc_2432, uc_2433, 
      uc_2434, uc_2435, uc_2436, uc_2437, uc_2438, uc_2439}), .in2({n_62, 
      uc_2440, uc_2441, uc_2442, uc_2443, uc_2444, uc_2445, uc_2446, uc_2447, 
      uc_2448, uc_2449, uc_2450, uc_2451, uc_2452, uc_2453, uc_2454, uc_2455, 
      uc_2456, uc_2457, uc_2458, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
      n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
      n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, uc_2459, 
      uc_2460, uc_2461, uc_2462, uc_2463, uc_2464, uc_2465, uc_2466, uc_2467, 
      uc_2468, uc_2469, uc_2470, uc_2471}), .in3({n_94, uc_2472, uc_2473, 
      uc_2474, uc_2475, uc_2476, uc_2477, uc_2478, uc_2479, uc_2480, uc_2481, 
      uc_2482, uc_2483, uc_2484, uc_2485, uc_2486, uc_2487, uc_2488, uc_2489, 
      n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, 
      n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, 
      n_69, n_68, n_67, n_66, n_65, n_64, n_63, uc_2490, uc_2491, uc_2492, 
      uc_2493, uc_2494, uc_2495, uc_2496, uc_2497, uc_2498, uc_2499, uc_2500, 
      uc_2501, uc_2502, uc_2503}), .sum({\s1[4] [45], uc_2504, uc_2505, uc_2506, 
      uc_2507, uc_2508, uc_2509, uc_2510, uc_2511, uc_2512, uc_2513, uc_2514, 
      uc_2515, uc_2516, uc_2517, uc_2518, uc_2519, uc_2520, uc_2521, \s1[4] [44], 
      \s1[4] [43], \s1[4] [42], \s1[4] [41], \s1[4] [40], \s1[4] [39], 
      \s1[4] [38], \s1[4] [37], \s1[4] [36], \s1[4] [35], \s1[4] [34], 
      \s1[4] [33], \s1[4] [32], \s1[4] [31], \s1[4] [30], \s1[4] [29], 
      \s1[4] [28], \s1[4] [27], \s1[4] [26], \s1[4] [25], \s1[4] [24], 
      \s1[4] [23], \s1[4] [22], \s1[4] [21], \s1[4] [20], \s1[4] [19], 
      \s1[4] [18], \s1[4] [17], \s1[4] [16], \s1[4] [15], \s1[4] [14], 
      \s1[4] [13], uc_2522, uc_2523, uc_2524, uc_2525, uc_2526, uc_2527, uc_2528, 
      uc_2529, uc_2530, uc_2531, uc_2532, uc_2533, uc_2534}), .c({\c1[4] [46], 
      uc_2535, uc_2536, uc_2537, uc_2538, uc_2539, uc_2540, uc_2541, uc_2542, 
      uc_2543, uc_2544, uc_2545, uc_2546, uc_2547, uc_2548, uc_2549, uc_2550, 
      uc_2551, \c1[4] [45], \c1[4] [44], \c1[4] [43], \c1[4] [42], \c1[4] [41], 
      \c1[4] [40], \c1[4] [39], \c1[4] [38], \c1[4] [37], \c1[4] [36], 
      \c1[4] [35], \c1[4] [34], \c1[4] [33], \c1[4] [32], \c1[4] [31], 
      \c1[4] [30], \c1[4] [29], \c1[4] [28], \c1[4] [27], \c1[4] [26], 
      \c1[4] [25], \c1[4] [24], \c1[4] [23], \c1[4] [22], \c1[4] [21], 
      \c1[4] [20], \c1[4] [19], \c1[4] [18], \c1[4] [17], \c1[4] [16], 
      \c1[4] [15], \s2[3] [14], uc_2552, uc_2553, uc_2554, uc_2555, uc_2556, 
      uc_2557, uc_2558, uc_2559, uc_2560, uc_2561, uc_2562, uc_2563, uc_2564, 
      uc_2565}));
   CSA__3_2 A5_1 (.in1({\s4[0] [46], uc_2566, uc_2567, uc_2568, uc_2569, uc_2570, 
      uc_2571, uc_2572, uc_2573, uc_2574, uc_2575, uc_2576, uc_2577, uc_2578, 
      uc_2579, uc_2580, uc_2581, uc_2582, \s4[0] [45], \s4[0] [44], \s4[0] [43], 
      \s4[0] [42], \s4[0] [41], \s4[0] [40], \s4[0] [39], \s4[0] [38], 
      \s4[0] [37], \s4[0] [36], \s4[0] [35], \s4[0] [34], \s4[0] [33], 
      \s4[0] [32], \s4[0] [31], \s4[0] [30], \s4[0] [29], \s4[0] [28], 
      \s4[0] [27], \s4[0] [26], \s4[0] [25], \s4[0] [24], \s4[0] [23], 
      \s4[0] [22], \s4[0] [21], \s4[0] [20], \s4[0] [19], \s4[0] [18], 
      \s4[0] [17], \s4[0] [16], \s4[0] [15], \s4[0] [14], \s4[0] [13], 
      \s4[0] [12], \s4[0] [11], \s4[0] [10], \s4[0] [9], \s4[0] [8], \s4[0] [7], 
      \s4[0] [6], \s4[0] [5], uc_2583, uc_2584, uc_2585, uc_2586, uc_2587}), 
      .in2({\c4[0] [47], uc_2588, uc_2589, uc_2590, uc_2591, uc_2592, uc_2593, 
      uc_2594, uc_2595, uc_2596, uc_2597, uc_2598, uc_2599, uc_2600, uc_2601, 
      uc_2602, uc_2603, \c4[0] [46], \c4[0] [45], \c4[0] [44], \c4[0] [43], 
      \c4[0] [42], \c4[0] [41], \c4[0] [40], \c4[0] [39], \c4[0] [38], 
      \c4[0] [37], \c4[0] [36], \c4[0] [35], \c4[0] [34], \c4[0] [33], 
      \c4[0] [32], \c4[0] [31], \c4[0] [30], \c4[0] [29], \c4[0] [28], 
      \c4[0] [27], \c4[0] [26], \c4[0] [25], \c4[0] [24], \c4[0] [23], 
      \c4[0] [22], \c4[0] [21], \c4[0] [20], \c4[0] [19], \c4[0] [18], 
      \c4[0] [17], \c4[0] [16], \c4[0] [15], \c4[0] [14], \c4[0] [13], 
      \c4[0] [12], \c4[0] [11], \c4[0] [10], \c4[0] [9], \c4[0] [8], \c4[0] [7], 
      \c4[0] [6], \c4[0] [5], uc_2604, uc_2605, uc_2606, uc_2607, uc_2608}), 
      .in3({\s4[1] [55], uc_2609, uc_2610, uc_2611, uc_2612, uc_2613, uc_2614, 
      uc_2615, uc_2616, \s4[1] [54], \s4[1] [53], \s4[1] [52], \s4[1] [51], 
      \s4[1] [50], \s4[1] [49], \s4[1] [48], \s4[1] [47], \s4[1] [46], 
      \s4[1] [45], \s4[1] [44], \s4[1] [43], \s4[1] [42], \s4[1] [41], 
      \s4[1] [40], \s4[1] [39], \s4[1] [38], \s4[1] [37], \s4[1] [36], 
      \s4[1] [35], \s4[1] [34], \s4[1] [33], \s4[1] [32], \s4[1] [31], 
      \s4[1] [30], \s4[1] [29], \s4[1] [28], \s4[1] [27], \s4[1] [26], 
      \s4[1] [25], \s4[1] [24], \s4[1] [23], \s4[1] [22], \s4[1] [21], 
      \s4[1] [20], \s4[1] [19], \s4[1] [18], \s4[1] [17], \s4[1] [16], 
      \s4[1] [15], \s4[1] [14], \c3[1] [13], \c3[1] [12], \c3[1] [11], 
      \c3[1] [10], uc_2617, uc_2618, uc_2619, uc_2620, uc_2621, uc_2622, uc_2623, 
      uc_2624, uc_2625, uc_2626}), .sum({\s5[0] [55], uc_2627, uc_2628, uc_2629, 
      uc_2630, uc_2631, uc_2632, uc_2633, uc_2634, \s5[0] [54], \s5[0] [53], 
      \s5[0] [52], \s5[0] [51], \s5[0] [50], \s5[0] [49], \s5[0] [48], 
      \s5[0] [47], \s5[0] [46], \s5[0] [45], \s5[0] [44], \s5[0] [43], 
      \s5[0] [42], \s5[0] [41], \s5[0] [40], \s5[0] [39], \s5[0] [38], 
      \s5[0] [37], \s5[0] [36], \s5[0] [35], \s5[0] [34], \s5[0] [33], 
      \s5[0] [32], \s5[0] [31], \s5[0] [30], \s5[0] [29], \s5[0] [28], 
      \s5[0] [27], \s5[0] [26], \s5[0] [25], \s5[0] [24], \s5[0] [23], 
      \s5[0] [22], \s5[0] [21], \s5[0] [20], \s5[0] [19], \s5[0] [18], 
      \s5[0] [17], \s5[0] [16], \s5[0] [15], \s5[0] [14], \s5[0] [13], 
      \s5[0] [12], \s5[0] [11], \s5[0] [10], \s5[0] [9], \s5[0] [8], \s5[0] [7], 
      \s5[0] [6], c[5], uc_2635, uc_2636, uc_2637, uc_2638, uc_2639}), .c({
      \c5[0] [56], uc_2640, uc_2641, uc_2642, uc_2643, uc_2644, uc_2645, uc_2646, 
      \c5[0] [55], \c5[0] [54], \c5[0] [53], \c5[0] [52], \c5[0] [51], 
      \c5[0] [50], \c5[0] [49], \c5[0] [48], \c5[0] [47], \c5[0] [46], 
      \c5[0] [45], \c5[0] [44], \c5[0] [43], \c5[0] [42], \c5[0] [41], 
      \c5[0] [40], \c5[0] [39], \c5[0] [38], \c5[0] [37], \c5[0] [36], 
      \c5[0] [35], \c5[0] [34], \c5[0] [33], \c5[0] [32], \c5[0] [31], 
      \c5[0] [30], \c5[0] [29], \c5[0] [28], \c5[0] [27], \c5[0] [26], 
      \c5[0] [25], \c5[0] [24], \c5[0] [23], \c5[0] [22], \c5[0] [21], 
      \c5[0] [20], \c5[0] [19], \c5[0] [18], \c5[0] [17], \c5[0] [16], 
      \c5[0] [15], \c5[0] [14], \c5[0] [13], \c5[0] [12], \c5[0] [11], 
      \c5[0] [10], \c5[0] [9], \c5[0] [8], \c5[0] [7], \c5[0] [6], uc_2647, 
      uc_2648, uc_2649, uc_2650, uc_2651, uc_2652}));
   CSA__3_5 A4_2 (.in1({\c3[1] [47], uc_2653, uc_2654, uc_2655, uc_2656, uc_2657, 
      uc_2658, uc_2659, uc_2660, uc_2661, uc_2662, uc_2663, uc_2664, uc_2665, 
      uc_2666, uc_2667, uc_2668, \c3[1] [46], \c3[1] [45], \c3[1] [44], 
      \c3[1] [43], \c3[1] [42], \c3[1] [41], \c3[1] [40], \c3[1] [39], 
      \c3[1] [38], \c3[1] [37], \c3[1] [36], \c3[1] [35], \c3[1] [34], 
      \c3[1] [33], \c3[1] [32], \c3[1] [31], \c3[1] [30], \c3[1] [29], 
      \c3[1] [28], \c3[1] [27], \c3[1] [26], \c3[1] [25], \c3[1] [24], 
      \c3[1] [23], \c3[1] [22], \c3[1] [21], \c3[1] [20], \c3[1] [19], 
      \c3[1] [18], \c3[1] [17], \c3[1] [16], \c3[1] [15], \c3[1] [14], uc_2669, 
      uc_2670, uc_2671, uc_2672, uc_2673, uc_2674, uc_2675, uc_2676, uc_2677, 
      uc_2678, uc_2679, uc_2680, uc_2681, uc_2682}), .in2({\s3[2] [54], uc_2683, 
      uc_2684, uc_2685, uc_2686, uc_2687, uc_2688, uc_2689, uc_2690, uc_2691, 
      \s3[2] [53], \s3[2] [52], \s3[2] [51], \s3[2] [50], \s3[2] [49], 
      \s3[2] [48], \s3[2] [47], \s3[2] [46], \s3[2] [45], \s3[2] [44], 
      \s3[2] [43], \s3[2] [42], \s3[2] [41], \s3[2] [40], \s3[2] [39], 
      \s3[2] [38], \s3[2] [37], \s3[2] [36], \s3[2] [35], \s3[2] [34], 
      \s3[2] [33], \s3[2] [32], \s3[2] [31], \s3[2] [30], \s3[2] [29], 
      \s3[2] [28], \s3[2] [27], \s3[2] [26], \s3[2] [25], \s3[2] [24], 
      \s3[2] [23], \s3[2] [22], \s3[2] [21], \s3[2] [20], \s3[2] [19], 
      \s3[2] [18], \s3[2] [17], \s3[2] [16], \s2[3] [15], \s2[3] [14], uc_2692, 
      uc_2693, uc_2694, uc_2695, uc_2696, uc_2697, uc_2698, uc_2699, uc_2700, 
      uc_2701, uc_2702, uc_2703, uc_2704, uc_2705}), .in3({\c3[2] [55], uc_2706, 
      uc_2707, uc_2708, uc_2709, uc_2710, uc_2711, uc_2712, uc_2713, \c3[2] [54], 
      \c3[2] [53], \c3[2] [52], \c3[2] [51], \c3[2] [50], \c3[2] [49], 
      \c3[2] [48], \c3[2] [47], \c3[2] [46], \c3[2] [45], \c3[2] [44], 
      \c3[2] [43], \c3[2] [42], \c3[2] [41], \c3[2] [40], \c3[2] [39], 
      \c3[2] [38], \c3[2] [37], \c3[2] [36], \c3[2] [35], \c3[2] [34], 
      \c3[2] [33], \c3[2] [32], \c3[2] [31], \c3[2] [30], \c3[2] [29], 
      \c3[2] [28], \c3[2] [27], \c3[2] [26], \c3[2] [25], \c3[2] [24], 
      \c3[2] [23], \c3[2] [22], \c3[2] [21], \c3[2] [20], \c3[2] [19], 
      \c3[2] [18], \c3[2] [17], uc_2714, uc_2715, uc_2716, uc_2717, uc_2718, 
      uc_2719, uc_2720, uc_2721, uc_2722, uc_2723, uc_2724, uc_2725, uc_2726, 
      uc_2727, uc_2728, uc_2729, uc_2730}), .sum({\s4[1] [55], uc_2731, uc_2732, 
      uc_2733, uc_2734, uc_2735, uc_2736, uc_2737, uc_2738, \s4[1] [54], 
      \s4[1] [53], \s4[1] [52], \s4[1] [51], \s4[1] [50], \s4[1] [49], 
      \s4[1] [48], \s4[1] [47], \s4[1] [46], \s4[1] [45], \s4[1] [44], 
      \s4[1] [43], \s4[1] [42], \s4[1] [41], \s4[1] [40], \s4[1] [39], 
      \s4[1] [38], \s4[1] [37], \s4[1] [36], \s4[1] [35], \s4[1] [34], 
      \s4[1] [33], \s4[1] [32], \s4[1] [31], \s4[1] [30], \s4[1] [29], 
      \s4[1] [28], \s4[1] [27], \s4[1] [26], \s4[1] [25], \s4[1] [24], 
      \s4[1] [23], \s4[1] [22], \s4[1] [21], \s4[1] [20], \s4[1] [19], 
      \s4[1] [18], \s4[1] [17], \s4[1] [16], \s4[1] [15], \s4[1] [14], uc_2739, 
      uc_2740, uc_2741, uc_2742, uc_2743, uc_2744, uc_2745, uc_2746, uc_2747, 
      uc_2748, uc_2749, uc_2750, uc_2751, uc_2752}), .c({\c4[1] [56], uc_2753, 
      uc_2754, uc_2755, uc_2756, uc_2757, uc_2758, uc_2759, \c4[1] [55], 
      \c4[1] [54], \c4[1] [53], \c4[1] [52], \c4[1] [51], \c4[1] [50], 
      \c4[1] [49], \c4[1] [48], \c4[1] [47], \c4[1] [46], \c4[1] [45], 
      \c4[1] [44], \c4[1] [43], \c4[1] [42], \c4[1] [41], \c4[1] [40], 
      \c4[1] [39], \c4[1] [38], \c4[1] [37], \c4[1] [36], \c4[1] [35], 
      \c4[1] [34], \c4[1] [33], \c4[1] [32], \c4[1] [31], \c4[1] [30], 
      \c4[1] [29], \c4[1] [28], \c4[1] [27], \c4[1] [26], \c4[1] [25], 
      \c4[1] [24], \c4[1] [23], \c4[1] [22], \c4[1] [21], \c4[1] [20], 
      \c4[1] [19], \c4[1] [18], \c4[1] [17], \c4[1] [16], \c4[1] [15], uc_2760, 
      uc_2761, uc_2762, uc_2763, uc_2764, uc_2765, uc_2766, uc_2767, uc_2768, 
      uc_2769, uc_2770, uc_2771, uc_2772, uc_2773, uc_2774}));
   CSA__3_8 A3_3 (.in1({\s2[3] [49], uc_2775, uc_2776, uc_2777, uc_2778, uc_2779, 
      uc_2780, uc_2781, uc_2782, uc_2783, uc_2784, uc_2785, uc_2786, uc_2787, 
      uc_2788, \s2[3] [48], \s2[3] [47], \s2[3] [46], \s2[3] [45], \s2[3] [44], 
      \s2[3] [43], \s2[3] [42], \s2[3] [41], \s2[3] [40], \s2[3] [39], 
      \s2[3] [38], \s2[3] [37], \s2[3] [36], \s2[3] [35], \s2[3] [34], 
      \s2[3] [33], \s2[3] [32], \s2[3] [31], \s2[3] [30], \s2[3] [29], 
      \s2[3] [28], \s2[3] [27], \s2[3] [26], \s2[3] [25], \s2[3] [24], 
      \s2[3] [23], \s2[3] [22], \s2[3] [21], \s2[3] [20], \s2[3] [19], 
      \s2[3] [18], \s2[3] [17], \s2[3] [16], uc_2789, uc_2790, uc_2791, uc_2792, 
      uc_2793, uc_2794, uc_2795, uc_2796, uc_2797, uc_2798, uc_2799, uc_2800, 
      uc_2801, uc_2802, uc_2803, uc_2804}), .in2({\c2[3] [50], uc_2805, uc_2806, 
      uc_2807, uc_2808, uc_2809, uc_2810, uc_2811, uc_2812, uc_2813, uc_2814, 
      uc_2815, uc_2816, uc_2817, \c2[3] [49], \c2[3] [48], \c2[3] [47], 
      \c2[3] [46], \c2[3] [45], \c2[3] [44], \c2[3] [43], \c2[3] [42], 
      \c2[3] [41], \c2[3] [40], \c2[3] [39], \c2[3] [38], \c2[3] [37], 
      \c2[3] [36], \c2[3] [35], \c2[3] [34], \c2[3] [33], \c2[3] [32], 
      \c2[3] [31], \c2[3] [30], \c2[3] [29], \c2[3] [28], \c2[3] [27], 
      \c2[3] [26], \c2[3] [25], \c2[3] [24], \c2[3] [23], \c2[3] [22], 
      \c2[3] [21], \c2[3] [20], \c2[3] [19], \c2[3] [18], \c2[3] [17], 
      \c2[3] [16], uc_2818, uc_2819, uc_2820, uc_2821, uc_2822, uc_2823, uc_2824, 
      uc_2825, uc_2826, uc_2827, uc_2828, uc_2829, uc_2830, uc_2831, uc_2832, 
      uc_2833}), .in3({\s2[4] [54], uc_2834, uc_2835, uc_2836, uc_2837, uc_2838, 
      uc_2839, uc_2840, uc_2841, uc_2842, \s2[4] [53], \s2[4] [52], \s2[4] [51], 
      \s2[4] [50], \s2[4] [49], \s2[4] [48], \s2[4] [47], \s2[4] [46], 
      \s2[4] [45], \s2[4] [44], \s2[4] [43], \s2[4] [42], \s2[4] [41], 
      \s2[4] [40], \s2[4] [39], \s2[4] [38], \s2[4] [37], \s2[4] [36], 
      \s2[4] [35], \s2[4] [34], \s2[4] [33], \s2[4] [32], \s2[4] [31], 
      \s2[4] [30], \s2[4] [29], \s2[4] [28], \s2[4] [27], \s2[4] [26], 
      \s2[4] [25], \s2[4] [24], \s2[4] [23], \s2[4] [22], \s2[4] [21], 
      \s2[4] [20], \s1[6] [19], n_191, uc_2843, uc_2844, uc_2845, uc_2846, 
      uc_2847, uc_2848, uc_2849, uc_2850, uc_2851, uc_2852, uc_2853, uc_2854, 
      uc_2855, uc_2856, uc_2857, uc_2858, uc_2859, uc_2860}), .sum({\s3[2] [54], 
      uc_2861, uc_2862, uc_2863, uc_2864, uc_2865, uc_2866, uc_2867, uc_2868, 
      uc_2869, \s3[2] [53], \s3[2] [52], \s3[2] [51], \s3[2] [50], \s3[2] [49], 
      \s3[2] [48], \s3[2] [47], \s3[2] [46], \s3[2] [45], \s3[2] [44], 
      \s3[2] [43], \s3[2] [42], \s3[2] [41], \s3[2] [40], \s3[2] [39], 
      \s3[2] [38], \s3[2] [37], \s3[2] [36], \s3[2] [35], \s3[2] [34], 
      \s3[2] [33], \s3[2] [32], \s3[2] [31], \s3[2] [30], \s3[2] [29], 
      \s3[2] [28], \s3[2] [27], \s3[2] [26], \s3[2] [25], \s3[2] [24], 
      \s3[2] [23], \s3[2] [22], \s3[2] [21], \s3[2] [20], \s3[2] [19], 
      \s3[2] [18], \s3[2] [17], \s3[2] [16], uc_2870, uc_2871, uc_2872, uc_2873, 
      uc_2874, uc_2875, uc_2876, uc_2877, uc_2878, uc_2879, uc_2880, uc_2881, 
      uc_2882, uc_2883, uc_2884, uc_2885}), .c({\c3[2] [55], uc_2886, uc_2887, 
      uc_2888, uc_2889, uc_2890, uc_2891, uc_2892, uc_2893, \c3[2] [54], 
      \c3[2] [53], \c3[2] [52], \c3[2] [51], \c3[2] [50], \c3[2] [49], 
      \c3[2] [48], \c3[2] [47], \c3[2] [46], \c3[2] [45], \c3[2] [44], 
      \c3[2] [43], \c3[2] [42], \c3[2] [41], \c3[2] [40], \c3[2] [39], 
      \c3[2] [38], \c3[2] [37], \c3[2] [36], \c3[2] [35], \c3[2] [34], 
      \c3[2] [33], \c3[2] [32], \c3[2] [31], \c3[2] [30], \c3[2] [29], 
      \c3[2] [28], \c3[2] [27], \c3[2] [26], \c3[2] [25], \c3[2] [24], 
      \c3[2] [23], \c3[2] [22], \c3[2] [21], \c3[2] [20], \c3[2] [19], 
      \c3[2] [18], \c3[2] [17], uc_2894, uc_2895, uc_2896, uc_2897, uc_2898, 
      uc_2899, uc_2900, uc_2901, uc_2902, uc_2903, uc_2904, uc_2905, uc_2906, 
      uc_2907, uc_2908, uc_2909, uc_2910}));
   CSA__3_11 A2_5 (.in1({\s1[6] [51], uc_2911, uc_2912, uc_2913, uc_2914, 
      uc_2915, uc_2916, uc_2917, uc_2918, uc_2919, uc_2920, uc_2921, uc_2922, 
      \s1[6] [50], \s1[6] [49], \s1[6] [48], \s1[6] [47], \s1[6] [46], 
      \s1[6] [45], \s1[6] [44], \s1[6] [43], \s1[6] [42], \s1[6] [41], 
      \s1[6] [40], \s1[6] [39], \s1[6] [38], \s1[6] [37], \s1[6] [36], 
      \s1[6] [35], \s1[6] [34], \s1[6] [33], \s1[6] [32], \s1[6] [31], 
      \s1[6] [30], \s1[6] [29], \s1[6] [28], \s1[6] [27], \s1[6] [26], 
      \s1[6] [25], \s1[6] [24], \s1[6] [23], \s1[6] [22], \s1[6] [21], 
      \s1[6] [20], uc_2923, uc_2924, uc_2925, uc_2926, uc_2927, uc_2928, uc_2929, 
      uc_2930, uc_2931, uc_2932, uc_2933, uc_2934, uc_2935, uc_2936, uc_2937, 
      uc_2938, uc_2939, uc_2940, uc_2941, uc_2942}), .in2({\c1[6] [52], uc_2943, 
      uc_2944, uc_2945, uc_2946, uc_2947, uc_2948, uc_2949, uc_2950, uc_2951, 
      uc_2952, uc_2953, \c1[6] [51], \c1[6] [50], \c1[6] [49], \c1[6] [48], 
      \c1[6] [47], \c1[6] [46], \c1[6] [45], \c1[6] [44], \c1[6] [43], 
      \c1[6] [42], \c1[6] [41], \c1[6] [40], \c1[6] [39], \c1[6] [38], 
      \c1[6] [37], \c1[6] [36], \c1[6] [35], \c1[6] [34], \c1[6] [33], 
      \c1[6] [32], \c1[6] [31], \c1[6] [30], \c1[6] [29], \c1[6] [28], 
      \c1[6] [27], \c1[6] [26], \c1[6] [25], \c1[6] [24], \c1[6] [23], 
      \c1[6] [22], \c1[6] [21], \c1[6] [20], uc_2954, uc_2955, uc_2956, uc_2957, 
      uc_2958, uc_2959, uc_2960, uc_2961, uc_2962, uc_2963, uc_2964, uc_2965, 
      uc_2966, uc_2967, uc_2968, uc_2969, uc_2970, uc_2971, uc_2972, uc_2973}), 
      .in3({\s1[7] [54], uc_2974, uc_2975, uc_2976, uc_2977, uc_2978, uc_2979, 
      uc_2980, uc_2981, uc_2982, \s1[7] [53], \s1[7] [52], \s1[7] [51], 
      \s1[7] [50], \s1[7] [49], \s1[7] [48], \s1[7] [47], \s1[7] [46], 
      \s1[7] [45], \s1[7] [44], \s1[7] [43], \s1[7] [42], \s1[7] [41], 
      \s1[7] [40], \s1[7] [39], \s1[7] [38], \s1[7] [37], \s1[7] [36], 
      \s1[7] [35], \s1[7] [34], \s1[7] [33], \s1[7] [32], \s1[7] [31], 
      \s1[7] [30], \s1[7] [29], \s1[7] [28], \s1[7] [27], \s1[7] [26], 
      \s1[7] [25], \s1[7] [24], \s1[7] [23], \s1[7] [22], \s1[7] [21], uc_2983, 
      uc_2984, uc_2985, uc_2986, uc_2987, uc_2988, uc_2989, uc_2990, uc_2991, 
      uc_2992, uc_2993, uc_2994, uc_2995, uc_2996, uc_2997, uc_2998, uc_2999, 
      uc_3000, uc_3001, uc_3002, uc_3003}), .sum({\s2[4] [54], uc_3004, uc_3005, 
      uc_3006, uc_3007, uc_3008, uc_3009, uc_3010, uc_3011, uc_3012, \s2[4] [53], 
      \s2[4] [52], \s2[4] [51], \s2[4] [50], \s2[4] [49], \s2[4] [48], 
      \s2[4] [47], \s2[4] [46], \s2[4] [45], \s2[4] [44], \s2[4] [43], 
      \s2[4] [42], \s2[4] [41], \s2[4] [40], \s2[4] [39], \s2[4] [38], 
      \s2[4] [37], \s2[4] [36], \s2[4] [35], \s2[4] [34], \s2[4] [33], 
      \s2[4] [32], \s2[4] [31], \s2[4] [30], \s2[4] [29], \s2[4] [28], 
      \s2[4] [27], \s2[4] [26], \s2[4] [25], \s2[4] [24], \s2[4] [23], 
      \s2[4] [22], \s2[4] [21], \s2[4] [20], uc_3013, uc_3014, uc_3015, uc_3016, 
      uc_3017, uc_3018, uc_3019, uc_3020, uc_3021, uc_3022, uc_3023, uc_3024, 
      uc_3025, uc_3026, uc_3027, uc_3028, uc_3029, uc_3030, uc_3031, uc_3032}), 
      .c({\c2[4] [55], uc_3033, uc_3034, uc_3035, uc_3036, uc_3037, uc_3038, 
      uc_3039, uc_3040, \c2[4] [54], \c2[4] [53], \c2[4] [52], \c2[4] [51], 
      \c2[4] [50], \c2[4] [49], \c2[4] [48], \c2[4] [47], \c2[4] [46], 
      \c2[4] [45], \c2[4] [44], \c2[4] [43], \c2[4] [42], \c2[4] [41], 
      \c2[4] [40], \c2[4] [39], \c2[4] [38], \c2[4] [37], \c2[4] [36], 
      \c2[4] [35], \c2[4] [34], \c2[4] [33], \c2[4] [32], \c2[4] [31], 
      \c2[4] [30], \c2[4] [29], \c2[4] [28], \c2[4] [27], \c2[4] [26], 
      \c2[4] [25], \c2[4] [24], \c2[4] [23], \c2[4] [22], \c2[4] [21], uc_3041, 
      uc_3042, uc_3043, uc_3044, uc_3045, uc_3046, uc_3047, uc_3048, uc_3049, 
      uc_3050, uc_3051, uc_3052, uc_3053, uc_3054, uc_3055, uc_3056, uc_3057, 
      uc_3058, uc_3059, uc_3060, uc_3061}));
   CSA__0_74 A1_7 (.in1({n_222, uc_3062, uc_3063, uc_3064, uc_3065, uc_3066, 
      uc_3067, uc_3068, uc_3069, uc_3070, uc_3071, uc_3072, uc_3073, uc_3074, 
      uc_3075, n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, 
      n_212, n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, 
      n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, n_193, 
      n_192, uc_3076, uc_3077, uc_3078, uc_3079, uc_3080, uc_3081, uc_3082, 
      uc_3083, uc_3084, uc_3085, uc_3086, uc_3087, uc_3088, uc_3089, uc_3090, 
      uc_3091, uc_3092, uc_3093, uc_3094}), .in2({n_254, uc_3095, uc_3096, 
      uc_3097, uc_3098, uc_3099, uc_3100, uc_3101, uc_3102, uc_3103, uc_3104, 
      uc_3105, uc_3106, uc_3107, n_253, n_252, n_251, n_250, n_249, n_248, n_247, 
      n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, n_238, n_237, 
      n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, n_228, n_227, 
      n_226, n_225, n_224, n_223, uc_3108, uc_3109, uc_3110, uc_3111, uc_3112, 
      uc_3113, uc_3114, uc_3115, uc_3116, uc_3117, uc_3118, uc_3119, uc_3120, 
      uc_3121, uc_3122, uc_3123, uc_3124, uc_3125, uc_3126}), .in3({n_286, 
      uc_3127, uc_3128, uc_3129, uc_3130, uc_3131, uc_3132, uc_3133, uc_3134, 
      uc_3135, uc_3136, uc_3137, uc_3138, n_285, n_284, n_283, n_282, n_281, 
      n_280, n_279, n_278, n_277, n_276, n_275, n_274, n_273, n_272, n_271, 
      n_270, n_269, n_268, n_267, n_266, n_265, n_264, n_263, n_262, n_261, 
      n_260, n_259, n_258, n_257, n_256, n_255, uc_3139, uc_3140, uc_3141, 
      uc_3142, uc_3143, uc_3144, uc_3145, uc_3146, uc_3147, uc_3148, uc_3149, 
      uc_3150, uc_3151, uc_3152, uc_3153, uc_3154, uc_3155, uc_3156, uc_3157, 
      uc_3158}), .sum({\s1[6] [51], uc_3159, uc_3160, uc_3161, uc_3162, uc_3163, 
      uc_3164, uc_3165, uc_3166, uc_3167, uc_3168, uc_3169, uc_3170, \s1[6] [50], 
      \s1[6] [49], \s1[6] [48], \s1[6] [47], \s1[6] [46], \s1[6] [45], 
      \s1[6] [44], \s1[6] [43], \s1[6] [42], \s1[6] [41], \s1[6] [40], 
      \s1[6] [39], \s1[6] [38], \s1[6] [37], \s1[6] [36], \s1[6] [35], 
      \s1[6] [34], \s1[6] [33], \s1[6] [32], \s1[6] [31], \s1[6] [30], 
      \s1[6] [29], \s1[6] [28], \s1[6] [27], \s1[6] [26], \s1[6] [25], 
      \s1[6] [24], \s1[6] [23], \s1[6] [22], \s1[6] [21], \s1[6] [20], 
      \s1[6] [19], uc_3171, uc_3172, uc_3173, uc_3174, uc_3175, uc_3176, uc_3177, 
      uc_3178, uc_3179, uc_3180, uc_3181, uc_3182, uc_3183, uc_3184, uc_3185, 
      uc_3186, uc_3187, uc_3188, uc_3189}), .c({\c1[6] [52], uc_3190, uc_3191, 
      uc_3192, uc_3193, uc_3194, uc_3195, uc_3196, uc_3197, uc_3198, uc_3199, 
      uc_3200, \c1[6] [51], \c1[6] [50], \c1[6] [49], \c1[6] [48], \c1[6] [47], 
      \c1[6] [46], \c1[6] [45], \c1[6] [44], \c1[6] [43], \c1[6] [42], 
      \c1[6] [41], \c1[6] [40], \c1[6] [39], \c1[6] [38], \c1[6] [37], 
      \c1[6] [36], \c1[6] [35], \c1[6] [34], \c1[6] [33], \c1[6] [32], 
      \c1[6] [31], \c1[6] [30], \c1[6] [29], \c1[6] [28], \c1[6] [27], 
      \c1[6] [26], \c1[6] [25], \c1[6] [24], \c1[6] [23], \c1[6] [22], 
      \c1[6] [21], \c1[6] [20], uc_3201, uc_3202, uc_3203, uc_3204, uc_3205, 
      uc_3206, uc_3207, uc_3208, uc_3209, uc_3210, uc_3211, uc_3212, uc_3213, 
      uc_3214, uc_3215, uc_3216, uc_3217, uc_3218, uc_3219, uc_3220}));
   CSA__4_2 A2_7 (.in1({\s1[9] [60], uc_3221, uc_3222, uc_3223, \s1[9] [59], 
      \s1[9] [58], \s1[9] [57], \s1[9] [56], \s1[9] [55], \s1[9] [54], 
      \s1[9] [53], \s1[9] [52], \s1[9] [51], \s1[9] [50], \s1[9] [49], 
      \s1[9] [48], \s1[9] [47], \s1[9] [46], \s1[9] [45], \s1[9] [44], 
      \s1[9] [43], \s1[9] [42], \s1[9] [41], \s1[9] [40], \s1[9] [39], 
      \s1[9] [38], \s1[9] [37], \s1[9] [36], \s1[9] [35], \s1[9] [34], 
      \s1[9] [33], \s1[9] [32], \s1[9] [31], \s1[9] [30], \s1[9] [29], uc_3224, 
      uc_3225, uc_3226, uc_3227, uc_3228, uc_3229, uc_3230, uc_3231, uc_3232, 
      uc_3233, uc_3234, uc_3235, uc_3236, uc_3237, uc_3238, uc_3239, uc_3240, 
      uc_3241, uc_3242, uc_3243, uc_3244, uc_3245, uc_3246, uc_3247, uc_3248, 
      uc_3249, uc_3250, uc_3251, uc_3252}), .in2({\c1[9] [61], uc_3253, uc_3254, 
      \c1[9] [60], \c1[9] [59], \c1[9] [58], \c1[9] [57], \c1[9] [56], 
      \c1[9] [55], \c1[9] [54], \c1[9] [53], \c1[9] [52], \c1[9] [51], 
      \c1[9] [50], \c1[9] [49], \c1[9] [48], \c1[9] [47], \c1[9] [46], 
      \c1[9] [45], \c1[9] [44], \c1[9] [43], \c1[9] [42], \c1[9] [41], 
      \c1[9] [40], \c1[9] [39], \c1[9] [38], \c1[9] [37], \c1[9] [36], 
      \c1[9] [35], \c1[9] [34], \c1[9] [33], \c1[9] [32], \c1[9] [31], 
      \c1[9] [30], \c1[9] [29], uc_3255, uc_3256, uc_3257, uc_3258, uc_3259, 
      uc_3260, uc_3261, uc_3262, uc_3263, uc_3264, uc_3265, uc_3266, uc_3267, 
      uc_3268, uc_3269, uc_3270, uc_3271, uc_3272, uc_3273, uc_3274, uc_3275, 
      uc_3276, uc_3277, uc_3278, uc_3279, uc_3280, uc_3281, uc_3282, uc_3283}), 
      .in3({n_414, uc_3284, uc_3285, n_413, n_412, n_411, n_410, n_409, n_408, 
      n_407, n_406, n_405, n_404, n_403, n_402, n_401, n_400, n_399, n_398, 
      n_397, n_396, n_395, n_394, n_393, n_392, n_391, n_390, n_389, n_388, 
      n_387, n_386, n_385, n_384, n_383, uc_3286, uc_3287, uc_3288, uc_3289, 
      uc_3290, uc_3291, uc_3292, uc_3293, uc_3294, uc_3295, uc_3296, uc_3297, 
      uc_3298, uc_3299, uc_3300, uc_3301, uc_3302, uc_3303, uc_3304, uc_3305, 
      uc_3306, uc_3307, uc_3308, uc_3309, uc_3310, uc_3311, uc_3312, uc_3313, 
      uc_3314, uc_3315}), .sum({\s2[6] [61], uc_3316, uc_3317, \s2[6] [60], 
      \s2[6] [59], \s2[6] [58], \s2[6] [57], \s2[6] [56], \s2[6] [55], 
      \s2[6] [54], \s2[6] [53], \s2[6] [52], \s2[6] [51], \s2[6] [50], 
      \s2[6] [49], \s2[6] [48], \s2[6] [47], \s2[6] [46], \s2[6] [45], 
      \s2[6] [44], \s2[6] [43], \s2[6] [42], \s2[6] [41], \s2[6] [40], 
      \s2[6] [39], \s2[6] [38], \s2[6] [37], \s2[6] [36], \s2[6] [35], 
      \s2[6] [34], \s2[6] [33], \s2[6] [32], \s2[6] [31], \s2[6] [30], 
      \s2[6] [29], uc_3318, uc_3319, uc_3320, uc_3321, uc_3322, uc_3323, uc_3324, 
      uc_3325, uc_3326, uc_3327, uc_3328, uc_3329, uc_3330, uc_3331, uc_3332, 
      uc_3333, uc_3334, uc_3335, uc_3336, uc_3337, uc_3338, uc_3339, uc_3340, 
      uc_3341, uc_3342, uc_3343, uc_3344, uc_3345, uc_3346}), .c({\c2[6] [62], 
      uc_3347, \c2[6] [61], \c2[6] [60], \c2[6] [59], \c2[6] [58], \c2[6] [57], 
      \c2[6] [56], \c2[6] [55], \c2[6] [54], \c2[6] [53], \c2[6] [52], 
      \c2[6] [51], \c2[6] [50], \c2[6] [49], \c2[6] [48], \c2[6] [47], 
      \c2[6] [46], \c2[6] [45], \c2[6] [44], \c2[6] [43], \c2[6] [42], 
      \c2[6] [41], \c2[6] [40], \c2[6] [39], \c2[6] [38], \c2[6] [37], 
      \c2[6] [36], \c2[6] [35], \c2[6] [34], \c2[6] [33], \c2[6] [32], 
      \c2[6] [31], \c2[6] [30], uc_3348, uc_3349, uc_3350, uc_3351, uc_3352, 
      uc_3353, uc_3354, uc_3355, uc_3356, uc_3357, uc_3358, uc_3359, uc_3360, 
      uc_3361, uc_3362, uc_3363, uc_3364, uc_3365, uc_3366, uc_3367, uc_3368, 
      uc_3369, uc_3370, uc_3371, uc_3372, uc_3373, uc_3374, uc_3375, uc_3376, 
      uc_3377}));
   CSA__4_5 A3_5 (.in1({\s2[6] [61], uc_3378, uc_3379, \s2[6] [60], \s2[6] [59], 
      \s2[6] [58], \s2[6] [57], \s2[6] [56], \s2[6] [55], \s2[6] [54], 
      \s2[6] [53], \s2[6] [52], \s2[6] [51], \s2[6] [50], \s2[6] [49], 
      \s2[6] [48], \s2[6] [47], \s2[6] [46], \s2[6] [45], \s2[6] [44], 
      \s2[6] [43], \s2[6] [42], \s2[6] [41], \s2[6] [40], \s2[6] [39], 
      \s2[6] [38], \s2[6] [37], \s2[6] [36], \s2[6] [35], \s2[6] [34], 
      \s2[6] [33], \s2[6] [32], \s2[6] [31], \s2[6] [30], uc_3380, uc_3381, 
      uc_3382, uc_3383, uc_3384, uc_3385, uc_3386, uc_3387, uc_3388, uc_3389, 
      uc_3390, uc_3391, uc_3392, uc_3393, uc_3394, uc_3395, uc_3396, uc_3397, 
      uc_3398, uc_3399, uc_3400, uc_3401, uc_3402, uc_3403, uc_3404, uc_3405, 
      uc_3406, uc_3407, uc_3408, uc_3409}), .in2({\c2[6] [62], uc_3410, 
      \c2[6] [61], \c2[6] [60], \c2[6] [59], \c2[6] [58], \c2[6] [57], 
      \c2[6] [56], \c2[6] [55], \c2[6] [54], \c2[6] [53], \c2[6] [52], 
      \c2[6] [51], \c2[6] [50], \c2[6] [49], \c2[6] [48], \c2[6] [47], 
      \c2[6] [46], \c2[6] [45], \c2[6] [44], \c2[6] [43], \c2[6] [42], 
      \c2[6] [41], \c2[6] [40], \c2[6] [39], \c2[6] [38], \c2[6] [37], 
      \c2[6] [36], \c2[6] [35], \c2[6] [34], \c2[6] [33], \c2[6] [32], 
      \c2[6] [31], \c2[6] [30], uc_3411, uc_3412, uc_3413, uc_3414, uc_3415, 
      uc_3416, uc_3417, uc_3418, uc_3419, uc_3420, uc_3421, uc_3422, uc_3423, 
      uc_3424, uc_3425, uc_3426, uc_3427, uc_3428, uc_3429, uc_3430, uc_3431, 
      uc_3432, uc_3433, uc_3434, uc_3435, uc_3436, uc_3437, uc_3438, uc_3439, 
      uc_3440}), .in3({n_446, uc_3441, n_445, n_444, n_443, n_442, n_441, n_440, 
      n_439, n_438, n_437, n_436, n_435, n_434, n_433, n_432, n_431, n_430, 
      n_429, n_428, n_427, n_426, n_425, n_424, n_423, n_422, n_421, n_420, 
      n_419, n_418, n_417, n_416, n_415, uc_3442, uc_3443, uc_3444, uc_3445, 
      uc_3446, uc_3447, uc_3448, uc_3449, uc_3450, uc_3451, uc_3452, uc_3453, 
      uc_3454, uc_3455, uc_3456, uc_3457, uc_3458, uc_3459, uc_3460, uc_3461, 
      uc_3462, uc_3463, uc_3464, uc_3465, uc_3466, uc_3467, uc_3468, uc_3469, 
      uc_3470, uc_3471, uc_3472}), .sum({\s3[4] [62], uc_3473, \s3[4] [61], 
      \s3[4] [60], \s3[4] [59], \s3[4] [58], \s3[4] [57], \s3[4] [56], 
      \s3[4] [55], \s3[4] [54], \s3[4] [53], \s3[4] [52], \s3[4] [51], 
      \s3[4] [50], \s3[4] [49], \s3[4] [48], \s3[4] [47], \s3[4] [46], 
      \s3[4] [45], \s3[4] [44], \s3[4] [43], \s3[4] [42], \s3[4] [41], 
      \s3[4] [40], \s3[4] [39], \s3[4] [38], \s3[4] [37], \s3[4] [36], 
      \s3[4] [35], \s3[4] [34], \s3[4] [33], \s3[4] [32], \s3[4] [31], 
      \s3[4] [30], uc_3474, uc_3475, uc_3476, uc_3477, uc_3478, uc_3479, uc_3480, 
      uc_3481, uc_3482, uc_3483, uc_3484, uc_3485, uc_3486, uc_3487, uc_3488, 
      uc_3489, uc_3490, uc_3491, uc_3492, uc_3493, uc_3494, uc_3495, uc_3496, 
      uc_3497, uc_3498, uc_3499, uc_3500, uc_3501, uc_3502, uc_3503}), .c({
      \c3[4] [63], \c3[4] [62], \c3[4] [61], \c3[4] [60], \c3[4] [59], 
      \c3[4] [58], \c3[4] [57], \c3[4] [56], \c3[4] [55], \c3[4] [54], 
      \c3[4] [53], \c3[4] [52], \c3[4] [51], \c3[4] [50], \c3[4] [49], 
      \c3[4] [48], \c3[4] [47], \c3[4] [46], \c3[4] [45], \c3[4] [44], 
      \c3[4] [43], \c3[4] [42], \c3[4] [41], \c3[4] [40], \c3[4] [39], 
      \c3[4] [38], \c3[4] [37], \c3[4] [36], \c3[4] [35], \c3[4] [34], 
      \c3[4] [33], \c3[4] [32], \c3[4] [31], uc_3504, uc_3505, uc_3506, uc_3507, 
      uc_3508, uc_3509, uc_3510, uc_3511, uc_3512, uc_3513, uc_3514, uc_3515, 
      uc_3516, uc_3517, uc_3518, uc_3519, uc_3520, uc_3521, uc_3522, uc_3523, 
      uc_3524, uc_3525, uc_3526, uc_3527, uc_3528, uc_3529, uc_3530, uc_3531, 
      uc_3532, uc_3533, uc_3534}));
   CSA__4_8 A4_3 (.in1({\s3[3] [59], uc_3535, uc_3536, uc_3537, uc_3538, 
      \s3[3] [58], \s3[3] [57], \s3[3] [56], \s3[3] [55], \s3[3] [54], 
      \s3[3] [53], \s3[3] [52], \s3[3] [51], \s3[3] [50], \s3[3] [49], 
      \s3[3] [48], \s3[3] [47], \s3[3] [46], \s3[3] [45], \s3[3] [44], 
      \s3[3] [43], \s3[3] [42], \s3[3] [41], \s3[3] [40], \s3[3] [39], 
      \s3[3] [38], \s3[3] [37], \s3[3] [36], \s3[3] [35], \s3[3] [34], 
      \s3[3] [33], \s3[3] [32], \s3[3] [31], \s3[3] [30], \s3[3] [29], 
      \s3[3] [28], \s3[3] [27], \s3[3] [26], \s3[3] [25], \s3[3] [24], uc_3539, 
      uc_3540, uc_3541, uc_3542, uc_3543, uc_3544, uc_3545, uc_3546, uc_3547, 
      uc_3548, uc_3549, uc_3550, uc_3551, uc_3552, uc_3553, uc_3554, uc_3555, 
      uc_3556, uc_3557, uc_3558, uc_3559, uc_3560, uc_3561, uc_3562}), .in2({
      \c3[3] [60], uc_3563, uc_3564, uc_3565, \c3[3] [59], \c3[3] [58], 
      \c3[3] [57], \c3[3] [56], \c3[3] [55], \c3[3] [54], \c3[3] [53], 
      \c3[3] [52], \c3[3] [51], \c3[3] [50], \c3[3] [49], \c3[3] [48], 
      \c3[3] [47], \c3[3] [46], \c3[3] [45], \c3[3] [44], \c3[3] [43], 
      \c3[3] [42], \c3[3] [41], \c3[3] [40], \c3[3] [39], \c3[3] [38], 
      \c3[3] [37], \c3[3] [36], \c3[3] [35], \c3[3] [34], \c3[3] [33], 
      \c3[3] [32], \c3[3] [31], \c3[3] [30], \c3[3] [29], \c3[3] [28], 
      \c3[3] [27], \c3[3] [26], \c3[3] [25], \c3[3] [24], uc_3566, uc_3567, 
      uc_3568, uc_3569, uc_3570, uc_3571, uc_3572, uc_3573, uc_3574, uc_3575, 
      uc_3576, uc_3577, uc_3578, uc_3579, uc_3580, uc_3581, uc_3582, uc_3583, 
      uc_3584, uc_3585, uc_3586, uc_3587, uc_3588, uc_3589}), .in3({\s3[4] [62], 
      uc_3590, \s3[4] [61], \s3[4] [60], \s3[4] [59], \s3[4] [58], \s3[4] [57], 
      \s3[4] [56], \s3[4] [55], \s3[4] [54], \s3[4] [53], \s3[4] [52], 
      \s3[4] [51], \s3[4] [50], \s3[4] [49], \s3[4] [48], \s3[4] [47], 
      \s3[4] [46], \s3[4] [45], \s3[4] [44], \s3[4] [43], \s3[4] [42], 
      \s3[4] [41], \s3[4] [40], \s3[4] [39], \s3[4] [38], \s3[4] [37], 
      \s3[4] [36], \s3[4] [35], \s3[4] [34], \s3[4] [33], \s3[4] [32], 
      \s3[4] [31], \s3[4] [30], \s2[6] [29], \s1[9] [28], n_287, uc_3591, 
      uc_3592, uc_3593, uc_3594, uc_3595, uc_3596, uc_3597, uc_3598, uc_3599, 
      uc_3600, uc_3601, uc_3602, uc_3603, uc_3604, uc_3605, uc_3606, uc_3607, 
      uc_3608, uc_3609, uc_3610, uc_3611, uc_3612, uc_3613, uc_3614, uc_3615, 
      uc_3616, uc_3617}), .sum({\s4[2] [62], uc_3618, \s4[2] [61], \s4[2] [60], 
      \s4[2] [59], \s4[2] [58], \s4[2] [57], \s4[2] [56], \s4[2] [55], 
      \s4[2] [54], \s4[2] [53], \s4[2] [52], \s4[2] [51], \s4[2] [50], 
      \s4[2] [49], \s4[2] [48], \s4[2] [47], \s4[2] [46], \s4[2] [45], 
      \s4[2] [44], \s4[2] [43], \s4[2] [42], \s4[2] [41], \s4[2] [40], 
      \s4[2] [39], \s4[2] [38], \s4[2] [37], \s4[2] [36], \s4[2] [35], 
      \s4[2] [34], \s4[2] [33], \s4[2] [32], \s4[2] [31], \s4[2] [30], 
      \s4[2] [29], \s4[2] [28], \s4[2] [27], \s4[2] [26], \s4[2] [25], 
      \s4[2] [24], uc_3619, uc_3620, uc_3621, uc_3622, uc_3623, uc_3624, uc_3625, 
      uc_3626, uc_3627, uc_3628, uc_3629, uc_3630, uc_3631, uc_3632, uc_3633, 
      uc_3634, uc_3635, uc_3636, uc_3637, uc_3638, uc_3639, uc_3640, uc_3641, 
      uc_3642}), .c({\c4[2] [63], \c4[2] [62], \c4[2] [61], \c4[2] [60], 
      \c4[2] [59], \c4[2] [58], \c4[2] [57], \c4[2] [56], \c4[2] [55], 
      \c4[2] [54], \c4[2] [53], \c4[2] [52], \c4[2] [51], \c4[2] [50], 
      \c4[2] [49], \c4[2] [48], \c4[2] [47], \c4[2] [46], \c4[2] [45], 
      \c4[2] [44], \c4[2] [43], \c4[2] [42], \c4[2] [41], \c4[2] [40], 
      \c4[2] [39], \c4[2] [38], \c4[2] [37], \c4[2] [36], \c4[2] [35], 
      \c4[2] [34], \c4[2] [33], \c4[2] [32], \c4[2] [31], \c4[2] [30], 
      \c4[2] [29], \c4[2] [28], \c4[2] [27], \c4[2] [26], \c4[2] [25], uc_3643, 
      uc_3644, uc_3645, uc_3646, uc_3647, uc_3648, uc_3649, uc_3650, uc_3651, 
      uc_3652, uc_3653, uc_3654, uc_3655, uc_3656, uc_3657, uc_3658, uc_3659, 
      uc_3660, uc_3661, uc_3662, uc_3663, uc_3664, uc_3665, uc_3666, uc_3667}));
   CSA__4_11 A5_2 (.in1({\c4[1] [56], uc_3668, uc_3669, uc_3670, uc_3671, 
      uc_3672, uc_3673, uc_3674, \c4[1] [55], \c4[1] [54], \c4[1] [53], 
      \c4[1] [52], \c4[1] [51], \c4[1] [50], \c4[1] [49], \c4[1] [48], 
      \c4[1] [47], \c4[1] [46], \c4[1] [45], \c4[1] [44], \c4[1] [43], 
      \c4[1] [42], \c4[1] [41], \c4[1] [40], \c4[1] [39], \c4[1] [38], 
      \c4[1] [37], \c4[1] [36], \c4[1] [35], \c4[1] [34], \c4[1] [33], 
      \c4[1] [32], \c4[1] [31], \c4[1] [30], \c4[1] [29], \c4[1] [28], 
      \c4[1] [27], \c4[1] [26], \c4[1] [25], \c4[1] [24], \c4[1] [23], 
      \c4[1] [22], \c4[1] [21], uc_3675, uc_3676, uc_3677, uc_3678, uc_3679, 
      uc_3680, uc_3681, uc_3682, uc_3683, uc_3684, uc_3685, uc_3686, uc_3687, 
      uc_3688, uc_3689, uc_3690, uc_3691, uc_3692, uc_3693, uc_3694, uc_3695}), 
      .in2({\s4[2] [62], uc_3696, \s4[2] [61], \s4[2] [60], \s4[2] [59], 
      \s4[2] [58], \s4[2] [57], \s4[2] [56], \s4[2] [55], \s4[2] [54], 
      \s4[2] [53], \s4[2] [52], \s4[2] [51], \s4[2] [50], \s4[2] [49], 
      \s4[2] [48], \s4[2] [47], \s4[2] [46], \s4[2] [45], \s4[2] [44], 
      \s4[2] [43], \s4[2] [42], \s4[2] [41], \s4[2] [40], \s4[2] [39], 
      \s4[2] [38], \s4[2] [37], \s4[2] [36], \s4[2] [35], \s4[2] [34], 
      \s4[2] [33], \s4[2] [32], \s4[2] [31], \s4[2] [30], \s4[2] [29], 
      \s4[2] [28], \s4[2] [27], \s4[2] [26], \s4[2] [25], \s4[2] [24], 
      \s3[3] [23], \c2[4] [22], \c2[4] [21], uc_3697, uc_3698, uc_3699, uc_3700, 
      uc_3701, uc_3702, uc_3703, uc_3704, uc_3705, uc_3706, uc_3707, uc_3708, 
      uc_3709, uc_3710, uc_3711, uc_3712, uc_3713, uc_3714, uc_3715, uc_3716, 
      uc_3717}), .in3({\c4[2] [63], \c4[2] [62], \c4[2] [61], \c4[2] [60], 
      \c4[2] [59], \c4[2] [58], \c4[2] [57], \c4[2] [56], \c4[2] [55], 
      \c4[2] [54], \c4[2] [53], \c4[2] [52], \c4[2] [51], \c4[2] [50], 
      \c4[2] [49], \c4[2] [48], \c4[2] [47], \c4[2] [46], \c4[2] [45], 
      \c4[2] [44], \c4[2] [43], \c4[2] [42], \c4[2] [41], \c4[2] [40], 
      \c4[2] [39], \c4[2] [38], \c4[2] [37], \c4[2] [36], \c4[2] [35], 
      \c4[2] [34], \c4[2] [33], \c4[2] [32], \c4[2] [31], \c4[2] [30], 
      \c4[2] [29], \c4[2] [28], \c4[2] [27], \c4[2] [26], \c4[2] [25], uc_3718, 
      uc_3719, uc_3720, uc_3721, uc_3722, uc_3723, uc_3724, uc_3725, uc_3726, 
      uc_3727, uc_3728, uc_3729, uc_3730, uc_3731, uc_3732, uc_3733, uc_3734, 
      uc_3735, uc_3736, uc_3737, uc_3738, uc_3739, uc_3740, uc_3741, uc_3742}), 
      .sum({\s5[1] [63], \s5[1] [62], \s5[1] [61], \s5[1] [60], \s5[1] [59], 
      \s5[1] [58], \s5[1] [57], \s5[1] [56], \s5[1] [55], \s5[1] [54], 
      \s5[1] [53], \s5[1] [52], \s5[1] [51], \s5[1] [50], \s5[1] [49], 
      \s5[1] [48], \s5[1] [47], \s5[1] [46], \s5[1] [45], \s5[1] [44], 
      \s5[1] [43], \s5[1] [42], \s5[1] [41], \s5[1] [40], \s5[1] [39], 
      \s5[1] [38], \s5[1] [37], \s5[1] [36], \s5[1] [35], \s5[1] [34], 
      \s5[1] [33], \s5[1] [32], \s5[1] [31], \s5[1] [30], \s5[1] [29], 
      \s5[1] [28], \s5[1] [27], \s5[1] [26], \s5[1] [25], \s5[1] [24], 
      \s5[1] [23], \s5[1] [22], \s5[1] [21], uc_3743, uc_3744, uc_3745, uc_3746, 
      uc_3747, uc_3748, uc_3749, uc_3750, uc_3751, uc_3752, uc_3753, uc_3754, 
      uc_3755, uc_3756, uc_3757, uc_3758, uc_3759, uc_3760, uc_3761, uc_3762, 
      uc_3763}), .c({\c5[1] [63], \c5[1] [62], \c5[1] [61], \c5[1] [60], 
      \c5[1] [59], \c5[1] [58], \c5[1] [57], \c5[1] [56], \c5[1] [55], 
      \c5[1] [54], \c5[1] [53], \c5[1] [52], \c5[1] [51], \c5[1] [50], 
      \c5[1] [49], \c5[1] [48], \c5[1] [47], \c5[1] [46], \c5[1] [45], 
      \c5[1] [44], \c5[1] [43], \c5[1] [42], \c5[1] [41], \c5[1] [40], 
      \c5[1] [39], \c5[1] [38], \c5[1] [37], \c5[1] [36], \c5[1] [35], 
      \c5[1] [34], \c5[1] [33], \c5[1] [32], \c5[1] [31], \c5[1] [30], 
      \c5[1] [29], \c5[1] [28], \c5[1] [27], \c5[1] [26], \c5[1] [25], 
      \c5[1] [24], \c5[1] [23], \c5[1] [22], uc_3764, uc_3765, uc_3766, uc_3767, 
      uc_3768, uc_3769, uc_3770, uc_3771, uc_3772, uc_3773, uc_3774, uc_3775, 
      uc_3776, uc_3777, uc_3778, uc_3779, uc_3780, uc_3781, uc_3782, uc_3783, 
      uc_3784, uc_3785}));
   CSA__4_14 A6 (.in1({\s5[0] [55], uc_3786, uc_3787, uc_3788, uc_3789, uc_3790, 
      uc_3791, uc_3792, uc_3793, \s5[0] [54], \s5[0] [53], \s5[0] [52], 
      \s5[0] [51], \s5[0] [50], \s5[0] [49], \s5[0] [48], \s5[0] [47], 
      \s5[0] [46], \s5[0] [45], \s5[0] [44], \s5[0] [43], \s5[0] [42], 
      \s5[0] [41], \s5[0] [40], \s5[0] [39], \s5[0] [38], \s5[0] [37], 
      \s5[0] [36], \s5[0] [35], \s5[0] [34], \s5[0] [33], \s5[0] [32], 
      \s5[0] [31], \s5[0] [30], \s5[0] [29], \s5[0] [28], \s5[0] [27], 
      \s5[0] [26], \s5[0] [25], \s5[0] [24], \s5[0] [23], \s5[0] [22], 
      \s5[0] [21], \s5[0] [20], \s5[0] [19], \s5[0] [18], \s5[0] [17], 
      \s5[0] [16], \s5[0] [15], \s5[0] [14], \s5[0] [13], \s5[0] [12], 
      \s5[0] [11], \s5[0] [10], \s5[0] [9], \s5[0] [8], \s5[0] [7], \s5[0] [6], 
      uc_3794, uc_3795, uc_3796, uc_3797, uc_3798, uc_3799}), .in2({\c5[0] [56], 
      uc_3800, uc_3801, uc_3802, uc_3803, uc_3804, uc_3805, uc_3806, \c5[0] [55], 
      \c5[0] [54], \c5[0] [53], \c5[0] [52], \c5[0] [51], \c5[0] [50], 
      \c5[0] [49], \c5[0] [48], \c5[0] [47], \c5[0] [46], \c5[0] [45], 
      \c5[0] [44], \c5[0] [43], \c5[0] [42], \c5[0] [41], \c5[0] [40], 
      \c5[0] [39], \c5[0] [38], \c5[0] [37], \c5[0] [36], \c5[0] [35], 
      \c5[0] [34], \c5[0] [33], \c5[0] [32], \c5[0] [31], \c5[0] [30], 
      \c5[0] [29], \c5[0] [28], \c5[0] [27], \c5[0] [26], \c5[0] [25], 
      \c5[0] [24], \c5[0] [23], \c5[0] [22], \c5[0] [21], \c5[0] [20], 
      \c5[0] [19], \c5[0] [18], \c5[0] [17], \c5[0] [16], \c5[0] [15], 
      \c5[0] [14], \c5[0] [13], \c5[0] [12], \c5[0] [11], \c5[0] [10], 
      \c5[0] [9], \c5[0] [8], \c5[0] [7], \c5[0] [6], uc_3807, uc_3808, uc_3809, 
      uc_3810, uc_3811, uc_3812}), .in3({\s5[1] [63], \s5[1] [62], \s5[1] [61], 
      \s5[1] [60], \s5[1] [59], \s5[1] [58], \s5[1] [57], \s5[1] [56], 
      \s5[1] [55], \s5[1] [54], \s5[1] [53], \s5[1] [52], \s5[1] [51], 
      \s5[1] [50], \s5[1] [49], \s5[1] [48], \s5[1] [47], \s5[1] [46], 
      \s5[1] [45], \s5[1] [44], \s5[1] [43], \s5[1] [42], \s5[1] [41], 
      \s5[1] [40], \s5[1] [39], \s5[1] [38], \s5[1] [37], \s5[1] [36], 
      \s5[1] [35], \s5[1] [34], \s5[1] [33], \s5[1] [32], \s5[1] [31], 
      \s5[1] [30], \s5[1] [29], \s5[1] [28], \s5[1] [27], \s5[1] [26], 
      \s5[1] [25], \s5[1] [24], \s5[1] [23], \s5[1] [22], \s5[1] [21], 
      \c4[1] [20], \c4[1] [19], \c4[1] [18], \c4[1] [17], \c4[1] [16], 
      \c4[1] [15], uc_3813, uc_3814, uc_3815, uc_3816, uc_3817, uc_3818, uc_3819, 
      uc_3820, uc_3821, uc_3822, uc_3823, uc_3824, uc_3825, uc_3826, uc_3827}), 
      .sum({s6[63], s6[62], s6[61], s6[60], s6[59], s6[58], s6[57], s6[56], 
      s6[55], s6[54], s6[53], s6[52], s6[51], s6[50], s6[49], s6[48], s6[47], 
      s6[46], s6[45], s6[44], s6[43], s6[42], s6[41], s6[40], s6[39], s6[38], 
      s6[37], s6[36], s6[35], s6[34], s6[33], s6[32], s6[31], s6[30], s6[29], 
      s6[28], s6[27], s6[26], s6[25], s6[24], s6[23], s6[22], s6[21], s6[20], 
      s6[19], s6[18], s6[17], s6[16], s6[15], s6[14], s6[13], s6[12], s6[11], 
      s6[10], s6[9], s6[8], s6[7], c[6], uc_3828, uc_3829, uc_3830, uc_3831, 
      uc_3832, uc_3833}), .c({c6[63], c6[62], c6[61], c6[60], c6[59], c6[58], 
      c6[57], c6[56], c6[55], c6[54], c6[53], c6[52], c6[51], c6[50], c6[49], 
      c6[48], c6[47], c6[46], c6[45], c6[44], c6[43], c6[42], c6[41], c6[40], 
      c6[39], c6[38], c6[37], c6[36], c6[35], c6[34], c6[33], c6[32], c6[31], 
      c6[30], c6[29], c6[28], c6[27], c6[26], c6[25], c6[24], c6[23], c6[22], 
      c6[21], c6[20], c6[19], c6[18], c6[17], c6[16], c6[15], c6[14], c6[13], 
      c6[12], c6[11], c6[10], c6[9], c6[8], c6[7], uc_3834, uc_3835, uc_3836, 
      uc_3837, uc_3838, uc_3839, uc_3840}));
   CSA__4_17 A7 (.in1({s6[63], s6[62], s6[61], s6[60], s6[59], s6[58], s6[57], 
      s6[56], s6[55], s6[54], s6[53], s6[52], s6[51], s6[50], s6[49], s6[48], 
      s6[47], s6[46], s6[45], s6[44], s6[43], s6[42], s6[41], s6[40], s6[39], 
      s6[38], s6[37], s6[36], s6[35], s6[34], s6[33], s6[32], s6[31], s6[30], 
      s6[29], s6[28], s6[27], s6[26], s6[25], s6[24], s6[23], s6[22], s6[21], 
      s6[20], s6[19], s6[18], s6[17], s6[16], s6[15], s6[14], s6[13], s6[12], 
      s6[11], s6[10], s6[9], s6[8], s6[7], uc_3841, uc_3842, uc_3843, uc_3844, 
      uc_3845, uc_3846, uc_3847}), .in2({c6[63], c6[62], c6[61], c6[60], c6[59], 
      c6[58], c6[57], c6[56], c6[55], c6[54], c6[53], c6[52], c6[51], c6[50], 
      c6[49], c6[48], c6[47], c6[46], c6[45], c6[44], c6[43], c6[42], c6[41], 
      c6[40], c6[39], c6[38], c6[37], c6[36], c6[35], c6[34], c6[33], c6[32], 
      c6[31], c6[30], c6[29], c6[28], c6[27], c6[26], c6[25], c6[24], c6[23], 
      c6[22], c6[21], c6[20], c6[19], c6[18], c6[17], c6[16], c6[15], c6[14], 
      c6[13], c6[12], c6[11], c6[10], c6[9], c6[8], c6[7], uc_3848, uc_3849, 
      uc_3850, uc_3851, uc_3852, uc_3853, uc_3854}), .in3({\c5[1] [63], 
      \c5[1] [62], \c5[1] [61], \c5[1] [60], \c5[1] [59], \c5[1] [58], 
      \c5[1] [57], \c5[1] [56], \c5[1] [55], \c5[1] [54], \c5[1] [53], 
      \c5[1] [52], \c5[1] [51], \c5[1] [50], \c5[1] [49], \c5[1] [48], 
      \c5[1] [47], \c5[1] [46], \c5[1] [45], \c5[1] [44], \c5[1] [43], 
      \c5[1] [42], \c5[1] [41], \c5[1] [40], \c5[1] [39], \c5[1] [38], 
      \c5[1] [37], \c5[1] [36], \c5[1] [35], \c5[1] [34], \c5[1] [33], 
      \c5[1] [32], \c5[1] [31], \c5[1] [30], \c5[1] [29], \c5[1] [28], 
      \c5[1] [27], \c5[1] [26], \c5[1] [25], \c5[1] [24], \c5[1] [23], 
      \c5[1] [22], uc_3855, uc_3856, uc_3857, uc_3858, uc_3859, uc_3860, uc_3861, 
      uc_3862, uc_3863, uc_3864, uc_3865, uc_3866, uc_3867, uc_3868, uc_3869, 
      uc_3870, uc_3871, uc_3872, uc_3873, uc_3874, uc_3875, uc_3876}), .sum({
      s7[63], s7[62], s7[61], s7[60], s7[59], s7[58], s7[57], s7[56], s7[55], 
      s7[54], s7[53], s7[52], s7[51], s7[50], s7[49], s7[48], s7[47], s7[46], 
      s7[45], s7[44], s7[43], s7[42], s7[41], s7[40], s7[39], s7[38], s7[37], 
      s7[36], s7[35], s7[34], s7[33], s7[32], s7[31], s7[30], s7[29], s7[28], 
      s7[27], s7[26], s7[25], s7[24], s7[23], s7[22], s7[21], s7[20], s7[19], 
      s7[18], s7[17], s7[16], s7[15], s7[14], s7[13], s7[12], s7[11], s7[10], 
      s7[9], s7[8], c[7], uc_3877, uc_3878, uc_3879, uc_3880, uc_3881, uc_3882, 
      uc_3883}), .c({c7[63], c7[62], c7[61], c7[60], c7[59], c7[58], c7[57], 
      c7[56], c7[55], c7[54], c7[53], c7[52], c7[51], c7[50], c7[49], c7[48], 
      c7[47], c7[46], c7[45], c7[44], c7[43], c7[42], c7[41], c7[40], c7[39], 
      c7[38], c7[37], c7[36], c7[35], c7[34], c7[33], c7[32], c7[31], c7[30], 
      c7[29], c7[28], c7[27], c7[26], c7[25], c7[24], c7[23], c7[22], c7[21], 
      c7[20], c7[19], c7[18], c7[17], c7[16], c7[15], c7[14], c7[13], c7[12], 
      c7[11], c7[10], c7[9], c7[8], uc_3884, uc_3885, uc_3886, uc_3887, uc_3888, 
      uc_3889, uc_3890, uc_3891}));
   CSA__4_20 A8 (.in1({s7[63], s7[62], s7[61], s7[60], s7[59], s7[58], s7[57], 
      s7[56], s7[55], s7[54], s7[53], s7[52], s7[51], s7[50], s7[49], s7[48], 
      s7[47], s7[46], s7[45], s7[44], s7[43], s7[42], s7[41], s7[40], s7[39], 
      s7[38], s7[37], s7[36], s7[35], s7[34], s7[33], s7[32], s7[31], s7[30], 
      s7[29], s7[28], s7[27], s7[26], s7[25], s7[24], s7[23], s7[22], s7[21], 
      s7[20], s7[19], s7[18], s7[17], s7[16], s7[15], s7[14], s7[13], s7[12], 
      s7[11], s7[10], s7[9], s7[8], uc_3892, uc_3893, uc_3894, uc_3895, uc_3896, 
      uc_3897, uc_3898, uc_3899}), .in2({c7[63], c7[62], c7[61], c7[60], c7[59], 
      c7[58], c7[57], c7[56], c7[55], c7[54], c7[53], c7[52], c7[51], c7[50], 
      c7[49], c7[48], c7[47], c7[46], c7[45], c7[44], c7[43], c7[42], c7[41], 
      c7[40], c7[39], c7[38], c7[37], c7[36], c7[35], c7[34], c7[33], c7[32], 
      c7[31], c7[30], c7[29], c7[28], c7[27], c7[26], c7[25], c7[24], c7[23], 
      c7[22], c7[21], c7[20], c7[19], c7[18], c7[17], c7[16], c7[15], c7[14], 
      c7[13], c7[12], c7[11], c7[10], c7[9], c7[8], uc_3900, uc_3901, uc_3902, 
      uc_3903, uc_3904, uc_3905, uc_3906, uc_3907}), .in3({\c3[4] [63], 
      \c3[4] [62], \c3[4] [61], \c3[4] [60], \c3[4] [59], \c3[4] [58], 
      \c3[4] [57], \c3[4] [56], \c3[4] [55], \c3[4] [54], \c3[4] [53], 
      \c3[4] [52], \c3[4] [51], \c3[4] [50], \c3[4] [49], \c3[4] [48], 
      \c3[4] [47], \c3[4] [46], \c3[4] [45], \c3[4] [44], \c3[4] [43], 
      \c3[4] [42], \c3[4] [41], \c3[4] [40], \c3[4] [39], \c3[4] [38], 
      \c3[4] [37], \c3[4] [36], \c3[4] [35], \c3[4] [34], \c3[4] [33], 
      \c3[4] [32], \c3[4] [31], uc_3908, uc_3909, uc_3910, uc_3911, uc_3912, 
      uc_3913, uc_3914, uc_3915, uc_3916, uc_3917, uc_3918, uc_3919, uc_3920, 
      uc_3921, uc_3922, uc_3923, uc_3924, uc_3925, uc_3926, uc_3927, uc_3928, 
      uc_3929, uc_3930, uc_3931, uc_3932, uc_3933, uc_3934, uc_3935, uc_3936, 
      uc_3937, uc_3938}), .sum({s8[63], s8[62], s8[61], s8[60], s8[59], s8[58], 
      s8[57], s8[56], s8[55], s8[54], s8[53], s8[52], s8[51], s8[50], s8[49], 
      s8[48], s8[47], s8[46], s8[45], s8[44], s8[43], s8[42], s8[41], s8[40], 
      s8[39], s8[38], s8[37], s8[36], s8[35], s8[34], s8[33], s8[32], s8[31], 
      s8[30], s8[29], s8[28], s8[27], s8[26], s8[25], s8[24], s8[23], s8[22], 
      s8[21], s8[20], s8[19], s8[18], s8[17], s8[16], s8[15], s8[14], s8[13], 
      s8[12], s8[11], s8[10], s8[9], c[8], uc_3939, uc_3940, uc_3941, uc_3942, 
      uc_3943, uc_3944, uc_3945, uc_3946}), .c({c8[63], c8[62], c8[61], c8[60], 
      c8[59], c8[58], c8[57], c8[56], c8[55], c8[54], c8[53], c8[52], c8[51], 
      c8[50], c8[49], c8[48], c8[47], c8[46], c8[45], c8[44], c8[43], c8[42], 
      c8[41], c8[40], c8[39], c8[38], c8[37], c8[36], c8[35], c8[34], c8[33], 
      c8[32], c8[31], c8[30], c8[29], c8[28], c8[27], c8[26], c8[25], c8[24], 
      c8[23], c8[22], c8[21], c8[20], c8[19], c8[18], c8[17], c8[16], c8[15], 
      c8[14], c8[13], c8[12], c8[11], c8[10], c8[9], uc_3947, uc_3948, uc_3949, 
      uc_3950, uc_3951, uc_3952, uc_3953, uc_3954, uc_3955}));
   CSA__4_23 A9 (.in1({s8[63], s8[62], s8[61], s8[60], s8[59], s8[58], s8[57], 
      s8[56], s8[55], s8[54], s8[53], s8[52], s8[51], s8[50], s8[49], s8[48], 
      s8[47], s8[46], s8[45], s8[44], s8[43], s8[42], s8[41], s8[40], s8[39], 
      s8[38], s8[37], s8[36], s8[35], s8[34], s8[33], s8[32], s8[31], s8[30], 
      s8[29], s8[28], s8[27], s8[26], s8[25], s8[24], s8[23], s8[22], s8[21], 
      s8[20], s8[19], s8[18], s8[17], s8[16], s8[15], s8[14], s8[13], s8[12], 
      s8[11], s8[10], s8[9], uc_3956, uc_3957, uc_3958, uc_3959, uc_3960, 
      uc_3961, uc_3962, uc_3963, uc_3964}), .in2({c8[63], c8[62], c8[61], c8[60], 
      c8[59], c8[58], c8[57], c8[56], c8[55], c8[54], c8[53], c8[52], c8[51], 
      c8[50], c8[49], c8[48], c8[47], c8[46], c8[45], c8[44], c8[43], c8[42], 
      c8[41], c8[40], c8[39], c8[38], c8[37], c8[36], c8[35], c8[34], c8[33], 
      c8[32], c8[31], c8[30], c8[29], c8[28], c8[27], c8[26], c8[25], c8[24], 
      c8[23], c8[22], c8[21], c8[20], c8[19], c8[18], c8[17], c8[16], c8[15], 
      c8[14], c8[13], c8[12], c8[11], c8[10], c8[9], uc_3965, uc_3966, uc_3967, 
      uc_3968, uc_3969, uc_3970, uc_3971, uc_3972, uc_3973}), .in3({uc_3974, 
      uc_3975, uc_3976, uc_3977, uc_3978, uc_3979, uc_3980, uc_3981, uc_3982, 
      uc_3983, uc_3984, uc_3985, uc_3986, uc_3987, uc_3988, uc_3989, uc_3990, 
      uc_3991, uc_3992, uc_3993, uc_3994, uc_3995, uc_3996, uc_3997, uc_3998, 
      uc_3999, uc_4000, uc_4001, uc_4002, uc_4003, uc_4004, uc_4005, b[31], 
      uc_4006, uc_4007, uc_4008, uc_4009, uc_4010, uc_4011, uc_4012, uc_4013, 
      uc_4014, uc_4015, uc_4016, uc_4017, uc_4018, uc_4019, uc_4020, uc_4021, 
      uc_4022, uc_4023, uc_4024, uc_4025, uc_4026, uc_4027, uc_4028, uc_4029, 
      uc_4030, uc_4031, uc_4032, uc_4033, uc_4034, uc_4035, uc_4036}), .sum({
      s9[63], s9[62], s9[61], s9[60], s9[59], s9[58], s9[57], s9[56], s9[55], 
      s9[54], s9[53], s9[52], s9[51], s9[50], s9[49], s9[48], s9[47], s9[46], 
      s9[45], s9[44], s9[43], s9[42], s9[41], s9[40], s9[39], s9[38], s9[37], 
      s9[36], s9[35], s9[34], s9[33], s9[32], s9[31], s9[30], s9[29], s9[28], 
      s9[27], s9[26], s9[25], s9[24], s9[23], s9[22], s9[21], s9[20], s9[19], 
      s9[18], s9[17], s9[16], s9[15], s9[14], s9[13], s9[12], s9[11], s9[10], 
      c[9], uc_4037, uc_4038, uc_4039, uc_4040, uc_4041, uc_4042, uc_4043, 
      uc_4044, uc_4045}), .c({c9[63], c9[62], c9[61], c9[60], c9[59], c9[58], 
      c9[57], c9[56], c9[55], c9[54], c9[53], c9[52], c9[51], c9[50], c9[49], 
      c9[48], c9[47], c9[46], c9[45], c9[44], c9[43], c9[42], c9[41], c9[40], 
      c9[39], c9[38], c9[37], c9[36], c9[35], c9[34], c9[33], c9[32], c9[31], 
      c9[30], c9[29], c9[28], c9[27], c9[26], c9[25], c9[24], c9[23], c9[22], 
      c9[21], c9[20], c9[19], c9[18], c9[17], c9[16], c9[15], c9[14], c9[13], 
      c9[12], c9[11], c9[10], uc_4046, uc_4047, uc_4048, uc_4049, uc_4050, 
      uc_4051, uc_4052, uc_4053, uc_4054, uc_4055}));
   simple_Adder RESULT (.a({s9[63], s9[62], s9[61], s9[60], s9[59], s9[58], 
      s9[57], s9[56], s9[55], s9[54], s9[53], s9[52], s9[51], s9[50], s9[49], 
      s9[48], s9[47], s9[46], s9[45], s9[44], s9[43], s9[42], s9[41], s9[40], 
      s9[39], s9[38], s9[37], s9[36], s9[35], s9[34], s9[33], s9[32], s9[31], 
      s9[30], s9[29], s9[28], s9[27], s9[26], s9[25], s9[24], s9[23], s9[22], 
      s9[21], s9[20], s9[19], s9[18], s9[17], s9[16], s9[15], s9[14], s9[13], 
      s9[12], s9[11], s9[10], uc_4056, uc_4057, uc_4058, uc_4059, uc_4060, 
      uc_4061, uc_4062, uc_4063, uc_4064, uc_4065}), .b({c9[63], c9[62], c9[61], 
      c9[60], c9[59], c9[58], c9[57], c9[56], c9[55], c9[54], c9[53], c9[52], 
      c9[51], c9[50], c9[49], c9[48], c9[47], c9[46], c9[45], c9[44], c9[43], 
      c9[42], c9[41], c9[40], c9[39], c9[38], c9[37], c9[36], c9[35], c9[34], 
      c9[33], c9[32], c9[31], c9[30], c9[29], c9[28], c9[27], c9[26], c9[25], 
      c9[24], c9[23], c9[22], c9[21], c9[20], c9[19], c9[18], c9[17], c9[16], 
      c9[15], c9[14], c9[13], c9[12], c9[11], c9[10], uc_4066, uc_4067, uc_4068, 
      uc_4069, uc_4070, uc_4071, uc_4072, uc_4073, uc_4074, uc_4075}), .cin(), 
      .S({c[63], c[62], c[61], c[60], c[59], c[58], c[57], c[56], c[55], c[54], 
      c[53], c[52], c[51], c[50], c[49], c[48], c[47], c[46], c[45], c[44], 
      c[43], c[42], c[41], c[40], c[39], c[38], c[37], c[36], c[35], c[34], 
      c[33], c[32], c[31], c[30], c[29], c[28], c[27], c[26], c[25], c[24], 
      c[23], c[22], c[21], c[20], c[19], c[18], c[17], c[16], c[15], c[14], 
      c[13], c[12], c[11], c[10], uc_4076, uc_4077, uc_4078, uc_4079, uc_4080, 
      uc_4081, uc_4082, uc_4083, uc_4084, uc_4085}));
   CSA A1_10 (.in1({n_318, uc_4086, uc_4087, uc_4088, uc_4089, uc_4090, n_317, 
      n_316, n_315, n_314, n_313, n_312, n_311, n_310, n_309, n_308, n_307, 
      n_306, n_305, n_304, n_303, n_302, n_301, n_300, n_299, n_298, n_297, 
      n_296, n_295, n_294, n_293, n_292, n_291, n_290, n_289, n_288, uc_4091, 
      uc_4092, uc_4093, uc_4094, uc_4095, uc_4096, uc_4097, uc_4098, uc_4099, 
      uc_4100, uc_4101, uc_4102, uc_4103, uc_4104, uc_4105, uc_4106, uc_4107, 
      uc_4108, uc_4109, uc_4110, uc_4111, uc_4112, uc_4113, uc_4114, uc_4115, 
      uc_4116, uc_4117, uc_4118}), .in2({n_350, uc_4119, uc_4120, uc_4121, 
      uc_4122, n_349, n_348, n_347, n_346, n_345, n_344, n_343, n_342, n_341, 
      n_340, n_339, n_338, n_337, n_336, n_335, n_334, n_333, n_332, n_331, 
      n_330, n_329, n_328, n_327, n_326, n_325, n_324, n_323, n_322, n_321, 
      n_320, n_319, uc_4123, uc_4124, uc_4125, uc_4126, uc_4127, uc_4128, 
      uc_4129, uc_4130, uc_4131, uc_4132, uc_4133, uc_4134, uc_4135, uc_4136, 
      uc_4137, uc_4138, uc_4139, uc_4140, uc_4141, uc_4142, uc_4143, uc_4144, 
      uc_4145, uc_4146, uc_4147, uc_4148, uc_4149, uc_4150}), .in3({n_382, 
      uc_4151, uc_4152, uc_4153, n_381, n_380, n_379, n_378, n_377, n_376, n_375, 
      n_374, n_373, n_372, n_371, n_370, n_369, n_368, n_367, n_366, n_365, 
      n_364, n_363, n_362, n_361, n_360, n_359, n_358, n_357, n_356, n_355, 
      n_354, n_353, n_352, n_351, uc_4154, uc_4155, uc_4156, uc_4157, uc_4158, 
      uc_4159, uc_4160, uc_4161, uc_4162, uc_4163, uc_4164, uc_4165, uc_4166, 
      uc_4167, uc_4168, uc_4169, uc_4170, uc_4171, uc_4172, uc_4173, uc_4174, 
      uc_4175, uc_4176, uc_4177, uc_4178, uc_4179, uc_4180, uc_4181, uc_4182}), 
      .sum({\s1[9] [60], uc_4183, uc_4184, uc_4185, \s1[9] [59], \s1[9] [58], 
      \s1[9] [57], \s1[9] [56], \s1[9] [55], \s1[9] [54], \s1[9] [53], 
      \s1[9] [52], \s1[9] [51], \s1[9] [50], \s1[9] [49], \s1[9] [48], 
      \s1[9] [47], \s1[9] [46], \s1[9] [45], \s1[9] [44], \s1[9] [43], 
      \s1[9] [42], \s1[9] [41], \s1[9] [40], \s1[9] [39], \s1[9] [38], 
      \s1[9] [37], \s1[9] [36], \s1[9] [35], \s1[9] [34], \s1[9] [33], 
      \s1[9] [32], \s1[9] [31], \s1[9] [30], \s1[9] [29], \s1[9] [28], uc_4186, 
      uc_4187, uc_4188, uc_4189, uc_4190, uc_4191, uc_4192, uc_4193, uc_4194, 
      uc_4195, uc_4196, uc_4197, uc_4198, uc_4199, uc_4200, uc_4201, uc_4202, 
      uc_4203, uc_4204, uc_4205, uc_4206, uc_4207, uc_4208, uc_4209, uc_4210, 
      uc_4211, uc_4212, uc_4213}), .c({\c1[9] [61], uc_4214, uc_4215, 
      \c1[9] [60], \c1[9] [59], \c1[9] [58], \c1[9] [57], \c1[9] [56], 
      \c1[9] [55], \c1[9] [54], \c1[9] [53], \c1[9] [52], \c1[9] [51], 
      \c1[9] [50], \c1[9] [49], \c1[9] [48], \c1[9] [47], \c1[9] [46], 
      \c1[9] [45], \c1[9] [44], \c1[9] [43], \c1[9] [42], \c1[9] [41], 
      \c1[9] [40], \c1[9] [39], \c1[9] [38], \c1[9] [37], \c1[9] [36], 
      \c1[9] [35], \c1[9] [34], \c1[9] [33], \c1[9] [32], \c1[9] [31], 
      \c1[9] [30], \c1[9] [29], uc_4216, uc_4217, uc_4218, uc_4219, uc_4220, 
      uc_4221, uc_4222, uc_4223, uc_4224, uc_4225, uc_4226, uc_4227, uc_4228, 
      uc_4229, uc_4230, uc_4231, uc_4232, uc_4233, uc_4234, uc_4235, uc_4236, 
      uc_4237, uc_4238, uc_4239, uc_4240, uc_4241, uc_4242, uc_4243, uc_4244}));
endmodule

module buffer__5_2(clk, rst, en, D, Q);
   input clk;
   input rst;
   input en;
   input [31:0]D;
   output [31:0]Q;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[31]  (.D(n_33), .CK(n_0), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_32), .CK(n_0), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_31), .CK(n_0), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_30), .CK(n_0), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_29), .CK(n_0), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_28), .CK(n_0), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_27), .CK(n_0), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_26), .CK(n_0), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_25), .CK(n_0), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_24), .CK(n_0), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_23), .CK(n_0), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_22), .CK(n_0), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_21), .CK(n_0), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_20), .CK(n_0), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_19), .CK(n_0), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_18), .CK(n_0), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_17), .CK(n_0), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_16), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_15), .CK(n_0), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_14), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_13), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_12), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_11), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_10), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_9), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_8), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_7), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_6), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_5), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_4), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_3), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_2), .CK(n_0), .Q(Q[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(rst), .ZN(n_1));
   INV_X1 i_0_1 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(D[31]), .ZN(n_33));
endmodule

module buffer(clk, rst, en, D, Q);
   input clk;
   input rst;
   input en;
   input [31:0]D;
   output [31:0]Q;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[31]  (.D(n_33), .CK(n_0), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_32), .CK(n_0), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_31), .CK(n_0), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_30), .CK(n_0), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_29), .CK(n_0), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_28), .CK(n_0), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_27), .CK(n_0), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_26), .CK(n_0), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_25), .CK(n_0), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_24), .CK(n_0), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_23), .CK(n_0), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_22), .CK(n_0), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_21), .CK(n_0), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_20), .CK(n_0), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_19), .CK(n_0), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_18), .CK(n_0), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_17), .CK(n_0), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_16), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_15), .CK(n_0), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_14), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_13), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_12), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_11), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_10), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_9), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_8), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_7), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_6), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_5), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_4), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_3), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_2), .CK(n_0), .Q(Q[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(rst), .ZN(n_1));
   INV_X1 i_0_1 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(D[31]), .ZN(n_33));
endmodule

module buffer__parameterized0(clk, rst, en, D, Q);
   input clk;
   input rst;
   input en;
   input [63:0]D;
   output [63:0]Q;

   wire n_0_1;
   wire n_0_0;

   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[63]  (.D(n_65), .CK(n_0), .Q(Q[63]), .QN());
   DFF_X1 \Q_reg[62]  (.D(n_64), .CK(n_0), .Q(Q[62]), .QN());
   DFF_X1 \Q_reg[61]  (.D(n_63), .CK(n_0), .Q(Q[61]), .QN());
   DFF_X1 \Q_reg[60]  (.D(n_62), .CK(n_0), .Q(Q[60]), .QN());
   DFF_X1 \Q_reg[59]  (.D(n_61), .CK(n_0), .Q(Q[59]), .QN());
   DFF_X1 \Q_reg[58]  (.D(n_60), .CK(n_0), .Q(Q[58]), .QN());
   DFF_X1 \Q_reg[57]  (.D(n_59), .CK(n_0), .Q(Q[57]), .QN());
   DFF_X1 \Q_reg[56]  (.D(n_58), .CK(n_0), .Q(Q[56]), .QN());
   DFF_X1 \Q_reg[55]  (.D(n_57), .CK(n_0), .Q(Q[55]), .QN());
   DFF_X1 \Q_reg[54]  (.D(n_56), .CK(n_0), .Q(Q[54]), .QN());
   DFF_X1 \Q_reg[53]  (.D(n_55), .CK(n_0), .Q(Q[53]), .QN());
   DFF_X1 \Q_reg[52]  (.D(n_54), .CK(n_0), .Q(Q[52]), .QN());
   DFF_X1 \Q_reg[51]  (.D(n_53), .CK(n_0), .Q(Q[51]), .QN());
   DFF_X1 \Q_reg[50]  (.D(n_52), .CK(n_0), .Q(Q[50]), .QN());
   DFF_X1 \Q_reg[49]  (.D(n_51), .CK(n_0), .Q(Q[49]), .QN());
   DFF_X1 \Q_reg[48]  (.D(n_50), .CK(n_0), .Q(Q[48]), .QN());
   DFF_X1 \Q_reg[47]  (.D(n_49), .CK(n_0), .Q(Q[47]), .QN());
   DFF_X1 \Q_reg[46]  (.D(n_48), .CK(n_0), .Q(Q[46]), .QN());
   DFF_X1 \Q_reg[45]  (.D(n_47), .CK(n_0), .Q(Q[45]), .QN());
   DFF_X1 \Q_reg[44]  (.D(n_46), .CK(n_0), .Q(Q[44]), .QN());
   DFF_X1 \Q_reg[43]  (.D(n_45), .CK(n_0), .Q(Q[43]), .QN());
   DFF_X1 \Q_reg[42]  (.D(n_44), .CK(n_0), .Q(Q[42]), .QN());
   DFF_X1 \Q_reg[41]  (.D(n_43), .CK(n_0), .Q(Q[41]), .QN());
   DFF_X1 \Q_reg[40]  (.D(n_42), .CK(n_0), .Q(Q[40]), .QN());
   DFF_X1 \Q_reg[39]  (.D(n_41), .CK(n_0), .Q(Q[39]), .QN());
   DFF_X1 \Q_reg[38]  (.D(n_40), .CK(n_0), .Q(Q[38]), .QN());
   DFF_X1 \Q_reg[37]  (.D(n_39), .CK(n_0), .Q(Q[37]), .QN());
   DFF_X1 \Q_reg[36]  (.D(n_38), .CK(n_0), .Q(Q[36]), .QN());
   DFF_X1 \Q_reg[35]  (.D(n_37), .CK(n_0), .Q(Q[35]), .QN());
   DFF_X1 \Q_reg[34]  (.D(n_36), .CK(n_0), .Q(Q[34]), .QN());
   DFF_X1 \Q_reg[33]  (.D(n_35), .CK(n_0), .Q(Q[33]), .QN());
   DFF_X1 \Q_reg[32]  (.D(n_34), .CK(n_0), .Q(Q[32]), .QN());
   DFF_X1 \Q_reg[31]  (.D(n_33), .CK(n_0), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_32), .CK(n_0), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_31), .CK(n_0), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_30), .CK(n_0), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_29), .CK(n_0), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_28), .CK(n_0), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_27), .CK(n_0), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_26), .CK(n_0), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_25), .CK(n_0), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_24), .CK(n_0), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_23), .CK(n_0), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_22), .CK(n_0), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_21), .CK(n_0), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_20), .CK(n_0), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_19), .CK(n_0), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_18), .CK(n_0), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_17), .CK(n_0), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_16), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_15), .CK(n_0), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_14), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_13), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_12), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_11), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_10), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_9), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_8), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_7), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_6), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_5), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_4), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_3), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_2), .CK(n_0), .Q(Q[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(rst), .ZN(n_1));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(D[31]), .ZN(n_33));
   AND2_X1 i_0_34 (.A1(n_0_0), .A2(D[32]), .ZN(n_34));
   AND2_X1 i_0_35 (.A1(n_0_0), .A2(D[33]), .ZN(n_35));
   AND2_X1 i_0_36 (.A1(n_0_0), .A2(D[34]), .ZN(n_36));
   AND2_X1 i_0_37 (.A1(n_0_0), .A2(D[35]), .ZN(n_37));
   AND2_X1 i_0_38 (.A1(n_0_0), .A2(D[36]), .ZN(n_38));
   AND2_X1 i_0_39 (.A1(n_0_0), .A2(D[37]), .ZN(n_39));
   AND2_X1 i_0_40 (.A1(n_0_0), .A2(D[38]), .ZN(n_40));
   AND2_X1 i_0_41 (.A1(n_0_0), .A2(D[39]), .ZN(n_41));
   AND2_X1 i_0_42 (.A1(n_0_0), .A2(D[40]), .ZN(n_42));
   AND2_X1 i_0_43 (.A1(n_0_0), .A2(D[41]), .ZN(n_43));
   AND2_X1 i_0_44 (.A1(n_0_0), .A2(D[42]), .ZN(n_44));
   AND2_X1 i_0_45 (.A1(n_0_0), .A2(D[43]), .ZN(n_45));
   AND2_X1 i_0_46 (.A1(n_0_0), .A2(D[44]), .ZN(n_46));
   AND2_X1 i_0_47 (.A1(n_0_0), .A2(D[45]), .ZN(n_47));
   AND2_X1 i_0_48 (.A1(n_0_0), .A2(D[46]), .ZN(n_48));
   AND2_X1 i_0_49 (.A1(n_0_0), .A2(D[47]), .ZN(n_49));
   AND2_X1 i_0_50 (.A1(n_0_0), .A2(D[48]), .ZN(n_50));
   AND2_X1 i_0_51 (.A1(n_0_0), .A2(D[49]), .ZN(n_51));
   AND2_X1 i_0_52 (.A1(n_0_0), .A2(D[50]), .ZN(n_52));
   AND2_X1 i_0_53 (.A1(n_0_0), .A2(D[51]), .ZN(n_53));
   AND2_X1 i_0_54 (.A1(n_0_0), .A2(D[52]), .ZN(n_54));
   AND2_X1 i_0_55 (.A1(n_0_0), .A2(D[53]), .ZN(n_55));
   AND2_X1 i_0_56 (.A1(n_0_0), .A2(D[54]), .ZN(n_56));
   AND2_X1 i_0_57 (.A1(n_0_0), .A2(D[55]), .ZN(n_57));
   AND2_X1 i_0_58 (.A1(n_0_0), .A2(D[56]), .ZN(n_58));
   AND2_X1 i_0_59 (.A1(n_0_0), .A2(D[57]), .ZN(n_59));
   AND2_X1 i_0_60 (.A1(n_0_0), .A2(D[58]), .ZN(n_60));
   AND2_X1 i_0_61 (.A1(n_0_0), .A2(D[59]), .ZN(n_61));
   AND2_X1 i_0_62 (.A1(n_0_0), .A2(D[60]), .ZN(n_62));
   AND2_X1 i_0_63 (.A1(n_0_0), .A2(D[61]), .ZN(n_63));
   AND2_X1 i_0_64 (.A1(n_0_0), .A2(D[62]), .ZN(n_64));
   INV_X1 i_0_1 (.A(rst), .ZN(n_0_1));
   AND2_X1 i_0_65 (.A1(D[63]), .A2(n_0_1), .ZN(n_65));
   BUF_X1 i_0_66 (.A(n_0_1), .Z(n_0_0));
endmodule

module multiplierTree(clk, rst, en, a, b, c);
   input clk;
   input rst;
   input en;
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   wire [63:0]c_out;
   wire [31:0]a_out;
   wire [31:0]b_out;

   wallace M64 (.a(a_out), .b(b_out), .c(c_out));
   buffer__5_2 inRegA (.clk(clk), .rst(rst), .en(en), .D(a), .Q(a_out));
   buffer inRegB (.clk(clk), .rst(rst), .en(en), .D(b), .Q(b_out));
   buffer__parameterized0 outReg (.clk(clk), .rst(rst), .en(en), .D(c_out), 
      .Q(c));
endmodule
