/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Jan  3 23:37:03 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3174960472 */

module CLA_4bit__0_53(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   AOI21_X1 i_0_0 (.A(n_0_11), .B1(n_0_10), .B2(n_0_2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(b[0]), .B(a[0]), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_6), .B(n_0_0), .ZN(sum[1]));
   XOR2_X1 i_0_3 (.A(b[1]), .B(a[1]), .Z(n_0_0));
   XNOR2_X1 i_0_4 (.A(n_0_5), .B(n_0_1), .ZN(sum[2]));
   XNOR2_X1 i_0_5 (.A(b[2]), .B(a[2]), .ZN(n_0_1));
   XNOR2_X1 i_0_6 (.A(n_0_9), .B(n_0_2), .ZN(sum[3]));
   OAI21_X1 i_0_7 (.A(n_0_3), .B1(a[2]), .B2(b[2]), .ZN(n_0_2));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_9 (.A(n_0_5), .B1(a[2]), .B2(b[2]), .ZN(n_0_4));
   OAI21_X1 i_0_10 (.A(n_0_7), .B1(n_0_8), .B2(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(b[0]), .A2(a[0]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(b[1]), .A2(a[1]), .ZN(n_0_7));
   NOR2_X1 i_0_13 (.A1(b[1]), .A2(a[1]), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[3]), .B(a[3]), .Z(n_0_9));
   NAND2_X1 i_0_15 (.A1(b[3]), .A2(a[3]), .ZN(n_0_10));
   NOR2_X1 i_0_16 (.A1(b[3]), .A2(a[3]), .ZN(n_0_11));
endmodule

module CLA_4bit__0_69(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_2), .B2(n_0_0), .ZN(cout));
   XOR2_X1 i_0_1 (.A(cin), .B(n_0_9), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_8), .B(n_0_6), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(n_0_5), .B(n_0_3), .ZN(sum[2]));
   XOR2_X1 i_0_4 (.A(n_0_2), .B(n_0_0), .Z(sum[3]));
   OAI21_X1 i_0_5 (.A(n_0_1), .B1(b[3]), .B2(a[3]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(b[3]), .A2(a[3]), .ZN(n_0_1));
   AOI22_X1 i_0_7 (.A1(b[2]), .A2(a[2]), .B1(n_0_4), .B2(n_0_3), .ZN(n_0_2));
   XOR2_X1 i_0_8 (.A(b[2]), .B(a[2]), .Z(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI22_X1 i_0_10 (.A1(b[1]), .A2(a[1]), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   XOR2_X1 i_0_11 (.A(b[1]), .B(a[1]), .Z(n_0_6));
   INV_X1 i_0_12 (.A(n_0_8), .ZN(n_0_7));
   AOI22_X1 i_0_13 (.A1(b[0]), .A2(a[0]), .B1(cin), .B2(n_0_9), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[0]), .B(a[0]), .Z(n_0_9));
endmodule

module CLA_4bit__0_77(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_2), .B2(n_0_0), .ZN(cout));
   XOR2_X1 i_0_1 (.A(cin), .B(n_0_9), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_8), .B(n_0_6), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(n_0_5), .B(n_0_3), .ZN(sum[2]));
   XOR2_X1 i_0_4 (.A(n_0_2), .B(n_0_0), .Z(sum[3]));
   OAI21_X1 i_0_5 (.A(n_0_1), .B1(b[3]), .B2(a[3]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(b[3]), .A2(a[3]), .ZN(n_0_1));
   AOI22_X1 i_0_7 (.A1(b[2]), .A2(a[2]), .B1(n_0_4), .B2(n_0_3), .ZN(n_0_2));
   XOR2_X1 i_0_8 (.A(b[2]), .B(a[2]), .Z(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI22_X1 i_0_10 (.A1(b[1]), .A2(a[1]), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   XOR2_X1 i_0_11 (.A(b[1]), .B(a[1]), .Z(n_0_6));
   INV_X1 i_0_12 (.A(n_0_8), .ZN(n_0_7));
   AOI22_X1 i_0_13 (.A1(b[0]), .A2(a[0]), .B1(cin), .B2(n_0_9), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[0]), .B(a[0]), .Z(n_0_9));
endmodule

module CLA_4bit__0_85(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_2), .B2(n_0_0), .ZN(cout));
   XOR2_X1 i_0_1 (.A(cin), .B(n_0_9), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_8), .B(n_0_6), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(n_0_5), .B(n_0_3), .ZN(sum[2]));
   XOR2_X1 i_0_4 (.A(n_0_2), .B(n_0_0), .Z(sum[3]));
   OAI21_X1 i_0_5 (.A(n_0_1), .B1(b[3]), .B2(a[3]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(b[3]), .A2(a[3]), .ZN(n_0_1));
   AOI22_X1 i_0_7 (.A1(b[2]), .A2(a[2]), .B1(n_0_4), .B2(n_0_3), .ZN(n_0_2));
   XOR2_X1 i_0_8 (.A(b[2]), .B(a[2]), .Z(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI22_X1 i_0_10 (.A1(b[1]), .A2(a[1]), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   XOR2_X1 i_0_11 (.A(b[1]), .B(a[1]), .Z(n_0_6));
   INV_X1 i_0_12 (.A(n_0_8), .ZN(n_0_7));
   AOI22_X1 i_0_13 (.A1(b[0]), .A2(a[0]), .B1(cin), .B2(n_0_9), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[0]), .B(a[0]), .Z(n_0_9));
endmodule

module CLA_4bit__0_93(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_2), .B2(n_0_0), .ZN(cout));
   XOR2_X1 i_0_1 (.A(cin), .B(n_0_9), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_8), .B(n_0_6), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(n_0_5), .B(n_0_3), .ZN(sum[2]));
   XOR2_X1 i_0_4 (.A(n_0_2), .B(n_0_0), .Z(sum[3]));
   OAI21_X1 i_0_5 (.A(n_0_1), .B1(b[3]), .B2(a[3]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(b[3]), .A2(a[3]), .ZN(n_0_1));
   AOI22_X1 i_0_7 (.A1(b[2]), .A2(a[2]), .B1(n_0_4), .B2(n_0_3), .ZN(n_0_2));
   XOR2_X1 i_0_8 (.A(b[2]), .B(a[2]), .Z(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI22_X1 i_0_10 (.A1(b[1]), .A2(a[1]), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   XOR2_X1 i_0_11 (.A(b[1]), .B(a[1]), .Z(n_0_6));
   INV_X1 i_0_12 (.A(n_0_8), .ZN(n_0_7));
   AOI22_X1 i_0_13 (.A1(b[0]), .A2(a[0]), .B1(cin), .B2(n_0_9), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[0]), .B(a[0]), .Z(n_0_9));
endmodule

module CLA_4bit__0_101(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_2), .B2(n_0_0), .ZN(cout));
   XOR2_X1 i_0_1 (.A(cin), .B(n_0_9), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_8), .B(n_0_6), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(n_0_5), .B(n_0_3), .ZN(sum[2]));
   XOR2_X1 i_0_4 (.A(n_0_2), .B(n_0_0), .Z(sum[3]));
   OAI21_X1 i_0_5 (.A(n_0_1), .B1(b[3]), .B2(a[3]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(b[3]), .A2(a[3]), .ZN(n_0_1));
   AOI22_X1 i_0_7 (.A1(b[2]), .A2(a[2]), .B1(n_0_4), .B2(n_0_3), .ZN(n_0_2));
   XOR2_X1 i_0_8 (.A(b[2]), .B(a[2]), .Z(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI22_X1 i_0_10 (.A1(b[1]), .A2(a[1]), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   XOR2_X1 i_0_11 (.A(b[1]), .B(a[1]), .Z(n_0_6));
   INV_X1 i_0_12 (.A(n_0_8), .ZN(n_0_7));
   AOI22_X1 i_0_13 (.A1(b[0]), .A2(a[0]), .B1(cin), .B2(n_0_9), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[0]), .B(a[0]), .Z(n_0_9));
endmodule

module CLA_4bit(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   XOR2_X1 i_0_0 (.A(a[3]), .B(cin), .Z(sum[0]));
endmodule

module CLA(in1, in2, cin, sum, cout, of);
   input [31:0]in1;
   input [31:0]in2;
   input cin;
   output [31:0]sum;
   output cout;
   output of;

   wire c;

   CLA_4bit__0_53 cla1 (.a({in1[3], in1[2], in1[1], in1[0]}), .b({in2[3], in2[2], 
      in2[1], in2[0]}), .cin(), .sum({sum[3], sum[2], sum[1], sum[0]}), .cout(c));
   CLA_4bit__0_69 genblk1_4_cla (.a({in1[7], in1[6], in1[5], in1[4]}), .b({
      in2[7], in2[6], in2[5], in2[4]}), .cin(c), .sum({sum[7], sum[6], sum[5], 
      sum[4]}), .cout(n_0));
   CLA_4bit__0_77 genblk1_8_cla (.a({in1[11], in1[10], in1[9], in1[8]}), 
      .b({in2[11], in2[10], in2[9], in2[8]}), .cin(n_0), .sum({sum[11], sum[10], 
      sum[9], sum[8]}), .cout(n_1));
   CLA_4bit__0_85 genblk1_12_cla (.a({in1[15], in1[14], in1[13], in1[12]}), 
      .b({in2[15], in2[14], in2[13], in2[12]}), .cin(n_1), .sum({sum[15], 
      sum[14], sum[13], sum[12]}), .cout(n_2));
   CLA_4bit__0_93 genblk1_16_cla (.a({in1[19], in1[18], in1[17], in1[16]}), 
      .b({in2[19], in2[18], in2[17], in2[16]}), .cin(n_2), .sum({sum[19], 
      sum[18], sum[17], sum[16]}), .cout(n_3));
   CLA_4bit__0_101 genblk1_20_cla (.a({in1[23], in1[22], in1[21], in1[20]}), 
      .b({in2[23], in2[22], in2[21], in2[20]}), .cin(n_3), .sum({sum[23], 
      sum[22], sum[21], sum[20]}), .cout(n_4));
   CLA_4bit genblk1_24_cla (.a({in1[31], uc_0, uc_1, uc_2}), .b(), .cin(n_4), 
      .sum({uc_3, uc_4, uc_5, sum[24]}), .cout());
endmodule

module count_leading_zeros(valueIn, result);
   input [22:0]valueIn;
   output [4:0]result;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;

   AOI21_X1 i_0_0 (.A(valueIn[22]), .B1(n_0_40), .B2(n_0_0), .ZN(result[0]));
   OAI21_X1 i_0_1 (.A(n_0_39), .B1(valueIn[19]), .B2(n_0_1), .ZN(n_0_0));
   AOI21_X1 i_0_2 (.A(valueIn[18]), .B1(n_0_38), .B2(n_0_2), .ZN(n_0_1));
   OAI21_X1 i_0_3 (.A(n_0_37), .B1(valueIn[15]), .B2(n_0_3), .ZN(n_0_2));
   AOI21_X1 i_0_4 (.A(valueIn[14]), .B1(n_0_36), .B2(n_0_4), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(n_0_35), .B1(valueIn[11]), .B2(n_0_5), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(valueIn[10]), .B1(n_0_34), .B2(n_0_6), .ZN(n_0_5));
   OAI21_X1 i_0_7 (.A(n_0_33), .B1(valueIn[7]), .B2(n_0_7), .ZN(n_0_6));
   AOI21_X1 i_0_8 (.A(valueIn[6]), .B1(n_0_32), .B2(n_0_8), .ZN(n_0_7));
   OAI21_X1 i_0_9 (.A(n_0_31), .B1(valueIn[3]), .B2(n_0_9), .ZN(n_0_8));
   AOI21_X1 i_0_10 (.A(valueIn[2]), .B1(n_0_30), .B2(valueIn[0]), .ZN(n_0_9));
   NOR3_X1 i_0_11 (.A1(valueIn[22]), .A2(valueIn[21]), .A3(n_0_10), .ZN(
      result[1]));
   NOR3_X1 i_0_12 (.A1(valueIn[20]), .A2(valueIn[19]), .A3(n_0_11), .ZN(n_0_10));
   NOR3_X1 i_0_13 (.A1(valueIn[18]), .A2(valueIn[17]), .A3(n_0_12), .ZN(n_0_11));
   NOR3_X1 i_0_14 (.A1(valueIn[16]), .A2(valueIn[15]), .A3(n_0_13), .ZN(n_0_12));
   NOR3_X1 i_0_15 (.A1(valueIn[14]), .A2(valueIn[13]), .A3(n_0_14), .ZN(n_0_13));
   AOI211_X1 i_0_16 (.A(valueIn[12]), .B(valueIn[11]), .C1(n_0_15), .C2(n_0_25), 
      .ZN(n_0_14));
   OAI21_X1 i_0_17 (.A(n_0_24), .B1(n_0_16), .B2(n_0_21), .ZN(n_0_15));
   NOR3_X1 i_0_18 (.A1(valueIn[4]), .A2(valueIn[3]), .A3(n_0_17), .ZN(n_0_16));
   NOR2_X1 i_0_19 (.A1(valueIn[2]), .A2(valueIn[1]), .ZN(n_0_17));
   AND2_X1 i_0_20 (.A1(n_0_18), .A2(n_0_29), .ZN(result[2]));
   NAND2_X1 i_0_21 (.A1(n_0_19), .A2(n_0_28), .ZN(n_0_18));
   OAI21_X1 i_0_22 (.A(n_0_26), .B1(n_0_20), .B2(n_0_23), .ZN(n_0_19));
   NOR3_X1 i_0_23 (.A1(n_0_21), .A2(valueIn[3]), .A3(valueIn[4]), .ZN(n_0_20));
   OR2_X1 i_0_24 (.A1(valueIn[6]), .A2(valueIn[5]), .ZN(n_0_21));
   AND3_X1 i_0_25 (.A1(n_0_22), .A2(n_0_28), .A3(n_0_29), .ZN(result[3]));
   NOR2_X1 i_0_26 (.A1(n_0_27), .A2(n_0_22), .ZN(result[4]));
   NAND3_X1 i_0_27 (.A1(n_0_26), .A2(n_0_25), .A3(n_0_24), .ZN(n_0_22));
   NAND2_X1 i_0_28 (.A1(n_0_25), .A2(n_0_24), .ZN(n_0_23));
   NOR2_X1 i_0_29 (.A1(valueIn[8]), .A2(valueIn[7]), .ZN(n_0_24));
   NOR2_X1 i_0_30 (.A1(valueIn[10]), .A2(valueIn[9]), .ZN(n_0_25));
   NOR4_X1 i_0_31 (.A1(valueIn[14]), .A2(valueIn[13]), .A3(valueIn[12]), 
      .A4(valueIn[11]), .ZN(n_0_26));
   NAND2_X1 i_0_32 (.A1(n_0_29), .A2(n_0_28), .ZN(n_0_27));
   NOR4_X1 i_0_33 (.A1(valueIn[18]), .A2(valueIn[17]), .A3(valueIn[16]), 
      .A4(valueIn[15]), .ZN(n_0_28));
   NOR4_X1 i_0_34 (.A1(valueIn[22]), .A2(valueIn[21]), .A3(valueIn[20]), 
      .A4(valueIn[19]), .ZN(n_0_29));
   INV_X1 i_0_35 (.A(valueIn[1]), .ZN(n_0_30));
   INV_X1 i_0_36 (.A(valueIn[4]), .ZN(n_0_31));
   INV_X1 i_0_37 (.A(valueIn[5]), .ZN(n_0_32));
   INV_X1 i_0_38 (.A(valueIn[8]), .ZN(n_0_33));
   INV_X1 i_0_39 (.A(valueIn[9]), .ZN(n_0_34));
   INV_X1 i_0_40 (.A(valueIn[12]), .ZN(n_0_35));
   INV_X1 i_0_41 (.A(valueIn[13]), .ZN(n_0_36));
   INV_X1 i_0_42 (.A(valueIn[16]), .ZN(n_0_37));
   INV_X1 i_0_43 (.A(valueIn[17]), .ZN(n_0_38));
   INV_X1 i_0_44 (.A(valueIn[20]), .ZN(n_0_39));
   INV_X1 i_0_45 (.A(valueIn[21]), .ZN(n_0_40));
endmodule

module datapath__0_23(p_0, exp_Sum, p_1);
   output p_0;
   input [7:0]exp_Sum;
   input [21:0]p_1;

   HA_X1 i_18 (.A(n_6), .B(n_4), .CO(n_18), .S());
   FA_X1 i_19 (.A(n_5), .B(n_7), .CI(n_18), .CO(n_0), .S());
   FA_X1 i_20 (.A(n_8), .B(n_11), .CI(n_0), .CO(n_1), .S());
   FA_X1 i_21 (.A(n_12), .B(n_15), .CI(n_1), .CO(n_2), .S());
   FA_X1 i_22 (.A(exp_Sum[5]), .B(n_16), .CI(n_2), .CO(n_3), .S());
   OAI21_X1 i_0 (.A(n_16), .B1(n_17), .B2(p_1[4]), .ZN(n_15));
   NAND2_X1 i_1 (.A1(n_17), .A2(p_1[4]), .ZN(n_16));
   OAI21_X1 i_2 (.A(n_12), .B1(n_14), .B2(p_1[3]), .ZN(n_11));
   NAND2_X1 i_3 (.A1(n_14), .A2(p_1[3]), .ZN(n_12));
   OAI21_X1 i_4 (.A(n_8), .B1(n_13), .B2(p_1[2]), .ZN(n_7));
   NAND2_X1 i_5 (.A1(n_13), .A2(p_1[2]), .ZN(n_8));
   OAI21_X1 i_6 (.A(n_5), .B1(n_10), .B2(p_1[1]), .ZN(n_4));
   NAND2_X1 i_7 (.A1(n_10), .A2(p_1[1]), .ZN(n_5));
   NAND2_X1 i_8 (.A1(n_9), .A2(p_1[11]), .ZN(n_6));
   NOR3_X1 i_9 (.A1(exp_Sum[7]), .A2(exp_Sum[6]), .A3(n_3), .ZN(p_0));
   INV_X1 i_10 (.A(exp_Sum[0]), .ZN(n_9));
   INV_X1 i_11 (.A(exp_Sum[1]), .ZN(n_10));
   INV_X1 i_12 (.A(exp_Sum[2]), .ZN(n_13));
   INV_X1 i_13 (.A(exp_Sum[3]), .ZN(n_14));
   INV_X1 i_14 (.A(exp_Sum[4]), .ZN(n_17));
endmodule

module datapath__0_36(p_0, p_1);
   input [21:0]p_0;
   output [10:0]p_1;

   INV_X1 i_0 (.A(p_0[11]), .ZN(p_1[0]));
   HA_X1 i_1 (.A(p_0[1]), .B(p_0[11]), .CO(n_0), .S(p_1[1]));
   HA_X1 i_2 (.A(p_0[2]), .B(n_0), .CO(n_1), .S(p_1[2]));
   HA_X1 i_3 (.A(p_0[3]), .B(n_1), .CO(n_2), .S(p_1[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_2), .CO(n_3), .S(p_1[4]));
endmodule

module datapath__0_41(mant_A, p_0);
   input [23:0]mant_A;
   output [31:0]p_0;

   XOR2_X1 i_0 (.A(mant_A[1]), .B(mant_A[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_21), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(mant_A[2]), .B1(mant_A[1]), .B2(mant_A[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(mant_A[3]), .B(n_21), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(mant_A[4]), .B(n_20), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(mant_A[5]), .B(n_19), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_18), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(mant_A[6]), .B1(n_19), .B2(mant_A[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(mant_A[7]), .B(n_18), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(mant_A[8]), .B(n_17), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_16), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(mant_A[9]), .B1(n_17), .B2(mant_A[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(mant_A[10]), .B(n_16), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(mant_A[11]), .B(n_15), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(mant_A[12]), .B(n_14), .Z(p_0[12]));
   XOR2_X1 i_15 (.A(mant_A[13]), .B(n_13), .Z(p_0[13]));
   XNOR2_X1 i_16 (.A(mant_A[14]), .B(n_12), .ZN(p_0[14]));
   XNOR2_X1 i_17 (.A(mant_A[15]), .B(n_11), .ZN(p_0[15]));
   XOR2_X1 i_18 (.A(mant_A[16]), .B(n_10), .Z(p_0[16]));
   XOR2_X1 i_19 (.A(mant_A[17]), .B(n_9), .Z(p_0[17]));
   XOR2_X1 i_20 (.A(mant_A[18]), .B(n_8), .Z(p_0[18]));
   AND2_X1 i_21 (.A1(n_7), .A2(n_3), .ZN(p_0[19]));
   OAI21_X1 i_22 (.A(mant_A[19]), .B1(n_8), .B2(mant_A[18]), .ZN(n_3));
   XOR2_X1 i_23 (.A(mant_A[20]), .B(n_7), .Z(p_0[20]));
   AND2_X1 i_24 (.A1(n_6), .A2(n_4), .ZN(p_0[21]));
   OAI21_X1 i_25 (.A(mant_A[21]), .B1(n_7), .B2(mant_A[20]), .ZN(n_4));
   XOR2_X1 i_26 (.A(mant_A[22]), .B(n_6), .Z(p_0[22]));
   AND2_X1 i_27 (.A1(p_0[31]), .A2(n_5), .ZN(p_0[23]));
   OAI21_X1 i_28 (.A(mant_A[23]), .B1(n_6), .B2(mant_A[22]), .ZN(n_5));
   OR3_X1 i_29 (.A1(n_6), .A2(mant_A[22]), .A3(mant_A[23]), .ZN(p_0[31]));
   OR3_X1 i_30 (.A1(n_7), .A2(mant_A[20]), .A3(mant_A[21]), .ZN(n_6));
   OR3_X1 i_31 (.A1(n_8), .A2(mant_A[18]), .A3(mant_A[19]), .ZN(n_7));
   OR2_X1 i_32 (.A1(n_9), .A2(mant_A[17]), .ZN(n_8));
   OR2_X1 i_33 (.A1(n_10), .A2(mant_A[16]), .ZN(n_9));
   NAND2_X1 i_34 (.A1(n_11), .A2(n_23), .ZN(n_10));
   NOR3_X1 i_35 (.A1(n_13), .A2(mant_A[13]), .A3(mant_A[14]), .ZN(n_11));
   NOR2_X1 i_36 (.A1(n_13), .A2(mant_A[13]), .ZN(n_12));
   OR2_X1 i_37 (.A1(n_14), .A2(mant_A[12]), .ZN(n_13));
   NAND2_X1 i_38 (.A1(n_15), .A2(n_22), .ZN(n_14));
   NOR2_X1 i_39 (.A1(n_16), .A2(mant_A[10]), .ZN(n_15));
   OR3_X1 i_40 (.A1(n_17), .A2(mant_A[8]), .A3(mant_A[9]), .ZN(n_16));
   OR2_X1 i_41 (.A1(n_18), .A2(mant_A[7]), .ZN(n_17));
   OR3_X1 i_42 (.A1(n_19), .A2(mant_A[5]), .A3(mant_A[6]), .ZN(n_18));
   OR2_X1 i_43 (.A1(n_20), .A2(mant_A[4]), .ZN(n_19));
   OR2_X1 i_44 (.A1(n_21), .A2(mant_A[3]), .ZN(n_20));
   OR3_X1 i_45 (.A1(mant_A[2]), .A2(mant_A[1]), .A3(mant_A[0]), .ZN(n_21));
   INV_X1 i_46 (.A(mant_A[11]), .ZN(n_22));
   INV_X1 i_47 (.A(mant_A[15]), .ZN(n_23));
endmodule

module fp_adder(A, B, Sum, overflow, underflow);
   input [31:0]A;
   input [31:0]B;
   output [31:0]Sum;
   output overflow;
   output underflow;

   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire [4:0]num_leading_zeros;
   wire n_0_30;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_0_7;
   wire n_0_0_0;
   wire n_0_0_8;
   wire n_0_0_1;
   wire n_0_0_9;
   wire n_0_0_2;
   wire n_0_0_10;
   wire n_0_0_3;
   wire n_0_0_11;
   wire n_0_0_4;
   wire n_0_0_12;
   wire n_0_0_5;
   wire n_0_0_13;
   wire n_0_0_6;
   wire [31:0]mant_A;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire [7:0]exp_Sum;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_55;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_56;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_57;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_58;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_59;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_60;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_61;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_62;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_63;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_64;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_65;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_66;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_67;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_68;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_69;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_70;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_71;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_72;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_73;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_74;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_75;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_0_369;
   wire n_0_76;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_77;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_78;
   wire n_0_0_392;
   wire n_0_79;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_80;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_81;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_82;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_83;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_416;
   wire n_0_84;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire n_0_85;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_86;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_430;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_0_433;
   wire n_0_87;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_88;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_0_439;
   wire n_0_89;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_90;
   wire n_0_0_443;
   wire n_0_0_444;
   wire n_0_0_445;
   wire n_0_91;
   wire n_0_0_446;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_92;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_0_451;
   wire n_0_93;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_94;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_462;
   wire n_0_0_463;
   wire n_0_95;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_96;
   wire n_0_0_466;
   wire n_0_0_467;
   wire n_0_97;
   wire n_0_0_468;
   wire n_0_0_469;
   wire n_0_98;
   wire n_0_0_470;
   wire n_0_0_471;
   wire n_0_0_472;
   wire n_0_0_473;
   wire n_0_99;
   wire n_0_0_474;
   wire n_0_0_475;
   wire n_0_0_476;
   wire n_0_0_477;
   wire n_0_100;
   wire n_0_0_478;
   wire n_0_0_479;
   wire n_0_0_480;
   wire n_0_0_481;
   wire n_0_0_482;
   wire n_0_0_483;
   wire n_0_0_484;
   wire n_0_101;
   wire n_0_0_485;
   wire n_0_0_486;
   wire n_0_0_487;
   wire n_0_0_488;
   wire n_0_0_489;
   wire n_0_0_490;
   wire n_0_0_491;
   wire n_0_0_492;
   wire n_0_0_493;
   wire n_0_0_494;
   wire n_0_0_495;
   wire n_0_0_496;
   wire n_0_0_497;
   wire n_0_0_498;
   wire n_0_0_499;
   wire n_0_0_500;
   wire n_0_0_501;
   wire n_0_0_502;
   wire n_0_0_503;
   wire n_0_0_504;
   wire n_0_0_505;
   wire n_0_0_506;
   wire n_0_0_507;
   wire n_0_0_508;
   wire n_0_0_509;
   wire n_0_0_510;
   wire n_0_0_511;
   wire n_0_0_512;
   wire n_0_0_513;
   wire n_0_102;
   wire n_0_0_514;
   wire n_0_0_515;
   wire n_0_0_516;
   wire n_0_0_517;
   wire n_0_0_518;
   wire n_0_0_519;
   wire n_0_0_520;
   wire n_0_0_521;
   wire n_0_0_522;
   wire n_0_0_523;
   wire n_0_0_524;
   wire n_0_0_525;
   wire n_0_0_526;
   wire n_0_0_527;
   wire n_0_0_528;
   wire n_0_0_529;
   wire n_0_0_530;
   wire n_0_0_531;
   wire n_0_0_532;
   wire n_0_0_533;
   wire n_0_0_534;
   wire n_0_0_535;
   wire n_0_0_536;
   wire n_0_0_537;
   wire n_0_0_538;
   wire n_0_0_539;
   wire n_0_0_540;
   wire n_0_0_541;
   wire n_0_0_542;
   wire n_0_0_543;
   wire n_0_0_544;
   wire n_0_0_545;
   wire n_0_0_546;
   wire n_0_0_547;
   wire n_0_0_548;
   wire n_0_0_549;
   wire n_0_0_550;
   wire n_0_0_551;
   wire n_0_0_552;
   wire n_0_0_553;
   wire n_0_0_554;
   wire n_0_0_555;
   wire n_0_0_556;
   wire n_0_0_557;
   wire n_0_0_558;
   wire n_0_0_559;
   wire n_0_0_560;
   wire n_0_0_561;
   wire n_0_0_562;
   wire n_0_0_563;
   wire n_0_0_564;
   wire n_0_0_565;
   wire n_0_0_566;
   wire n_0_0_567;
   wire n_0_0_568;
   wire n_0_0_569;
   wire n_0_0_570;
   wire n_0_0_571;
   wire n_0_0_572;
   wire n_0_0_573;
   wire n_0_0_574;
   wire n_0_0_575;
   wire n_0_0_576;
   wire n_0_0_577;
   wire n_0_0_578;
   wire n_0_0_579;
   wire n_0_0_580;
   wire n_0_0_581;
   wire n_0_0_582;
   wire n_0_0_583;
   wire n_0_0_584;
   wire n_0_0_585;
   wire n_0_0_586;
   wire n_0_0_587;
   wire n_0_0_588;
   wire n_0_0_589;
   wire n_0_0_590;
   wire n_0_0_591;
   wire n_0_0_592;
   wire n_0_0_593;
   wire n_0_0_594;
   wire n_0_0_595;
   wire n_0_0_596;
   wire n_0_0_597;
   wire n_0_0_598;
   wire n_0_0_599;
   wire n_0_0_600;

   CLA CLA_dut (.in1({mant_A[31], uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, 
      mant_A[23], mant_A[22], mant_A[21], mant_A[20], mant_A[19], mant_A[18], 
      mant_A[17], mant_A[16], mant_A[15], mant_A[14], mant_A[13], mant_A[12], 
      mant_A[11], mant_A[10], mant_A[9], mant_A[8], mant_A[7], mant_A[6], 
      mant_A[5], mant_A[4], mant_A[3], mant_A[2], mant_A[1], n_0_55}), .in2({
      uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, n_0_102, n_0_101, 
      n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, 
      n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, 
      n_0_82, n_0_81, n_0_80, n_0_79}), .cin(), .sum({uc_15, uc_16, uc_17, uc_18, 
      uc_19, uc_20, uc_21, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, 
      n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, 
      n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5}), 
      .cout(), .of());
   count_leading_zeros count_leading_zeros_instance (.valueIn({n_0_27, n_0_26, 
      n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, 
      n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, 
      n_0_7, n_0_6, n_0_5}), .result(num_leading_zeros));
   datapath__0_23 i_0_6 (.p_0(n_0_30), .exp_Sum(exp_Sum), .p_1({1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, num_leading_zeros[0], 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, num_leading_zeros[4], num_leading_zeros[3], 
      num_leading_zeros[2], num_leading_zeros[1], 1'b1}));
   datapath__0_36 i_0_18 (.p_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, num_leading_zeros[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      num_leading_zeros[4], num_leading_zeros[3], num_leading_zeros[2], 
      num_leading_zeros[1], 1'b1}), .p_1({uc_22, uc_23, uc_24, uc_25, uc_26, 
      uc_27, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0}));
   datapath__0_41 i_0_23 (.mant_A({n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, 
      n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, 
      n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, 
      n_0_55}), .p_0({n_0_54, uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, 
      n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, 
      n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, 
      n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, uc_35}));
   HA_X1 i_0_0_0 (.A(n_0_29), .B(exp_Sum[0]), .CO(n_0_0_0), .S(n_0_0_7));
   HA_X1 i_0_0_1 (.A(exp_Sum[1]), .B(n_0_0_0), .CO(n_0_0_1), .S(n_0_0_8));
   HA_X1 i_0_0_2 (.A(exp_Sum[2]), .B(n_0_0_1), .CO(n_0_0_2), .S(n_0_0_9));
   HA_X1 i_0_0_3 (.A(exp_Sum[3]), .B(n_0_0_2), .CO(n_0_0_3), .S(n_0_0_10));
   HA_X1 i_0_0_4 (.A(exp_Sum[4]), .B(n_0_0_3), .CO(n_0_0_4), .S(n_0_0_11));
   HA_X1 i_0_0_5 (.A(exp_Sum[5]), .B(n_0_0_4), .CO(n_0_0_5), .S(n_0_0_12));
   HA_X1 i_0_0_6 (.A(exp_Sum[6]), .B(n_0_0_5), .CO(n_0_0_6), .S(n_0_0_13));
   AOI21_X1 i_0_0_7 (.A(n_0_0_14), .B1(n_0_0_273), .B2(n_0_0_180), .ZN(mant_A[1]));
   NOR2_X1 i_0_0_8 (.A1(n_0_31), .A2(n_0_0_180), .ZN(n_0_0_14));
   AOI21_X1 i_0_0_9 (.A(n_0_0_15), .B1(n_0_0_277), .B2(n_0_0_180), .ZN(mant_A[2]));
   NOR2_X1 i_0_0_10 (.A1(n_0_32), .A2(n_0_0_180), .ZN(n_0_0_15));
   AOI21_X1 i_0_0_11 (.A(n_0_0_16), .B1(n_0_0_282), .B2(n_0_0_180), .ZN(
      mant_A[3]));
   NOR2_X1 i_0_0_12 (.A1(n_0_33), .A2(n_0_0_180), .ZN(n_0_0_16));
   AOI21_X1 i_0_0_13 (.A(n_0_0_17), .B1(n_0_0_288), .B2(n_0_0_180), .ZN(
      mant_A[4]));
   NOR2_X1 i_0_0_14 (.A1(n_0_34), .A2(n_0_0_180), .ZN(n_0_0_17));
   AOI21_X1 i_0_0_15 (.A(n_0_0_18), .B1(n_0_0_293), .B2(n_0_0_180), .ZN(
      mant_A[5]));
   NOR2_X1 i_0_0_16 (.A1(n_0_35), .A2(n_0_0_180), .ZN(n_0_0_18));
   AOI21_X1 i_0_0_17 (.A(n_0_0_19), .B1(n_0_0_298), .B2(n_0_0_180), .ZN(
      mant_A[6]));
   NOR2_X1 i_0_0_18 (.A1(n_0_36), .A2(n_0_0_180), .ZN(n_0_0_19));
   AOI21_X1 i_0_0_19 (.A(n_0_0_20), .B1(n_0_0_304), .B2(n_0_0_180), .ZN(
      mant_A[7]));
   NOR2_X1 i_0_0_20 (.A1(n_0_37), .A2(n_0_0_180), .ZN(n_0_0_20));
   AOI21_X1 i_0_0_21 (.A(n_0_0_21), .B1(n_0_0_308), .B2(n_0_0_180), .ZN(
      mant_A[8]));
   NOR2_X1 i_0_0_22 (.A1(n_0_38), .A2(n_0_0_180), .ZN(n_0_0_21));
   AOI21_X1 i_0_0_23 (.A(n_0_0_22), .B1(n_0_0_314), .B2(n_0_0_180), .ZN(
      mant_A[9]));
   NOR2_X1 i_0_0_24 (.A1(n_0_39), .A2(n_0_0_180), .ZN(n_0_0_22));
   AOI21_X1 i_0_0_25 (.A(n_0_0_23), .B1(n_0_0_317), .B2(n_0_0_180), .ZN(
      mant_A[10]));
   NOR2_X1 i_0_0_26 (.A1(n_0_40), .A2(n_0_0_180), .ZN(n_0_0_23));
   AOI21_X1 i_0_0_27 (.A(n_0_0_24), .B1(n_0_0_324), .B2(n_0_0_180), .ZN(
      mant_A[11]));
   NOR2_X1 i_0_0_28 (.A1(n_0_41), .A2(n_0_0_180), .ZN(n_0_0_24));
   AOI21_X1 i_0_0_29 (.A(n_0_0_25), .B1(n_0_0_329), .B2(n_0_0_180), .ZN(
      mant_A[12]));
   NOR2_X1 i_0_0_30 (.A1(n_0_42), .A2(n_0_0_180), .ZN(n_0_0_25));
   AOI21_X1 i_0_0_31 (.A(n_0_0_26), .B1(n_0_0_332), .B2(n_0_0_180), .ZN(
      mant_A[13]));
   NOR2_X1 i_0_0_32 (.A1(n_0_43), .A2(n_0_0_180), .ZN(n_0_0_26));
   AOI21_X1 i_0_0_33 (.A(n_0_0_27), .B1(n_0_0_337), .B2(n_0_0_180), .ZN(
      mant_A[14]));
   NOR2_X1 i_0_0_34 (.A1(n_0_44), .A2(n_0_0_180), .ZN(n_0_0_27));
   AOI21_X1 i_0_0_35 (.A(n_0_0_28), .B1(n_0_0_341), .B2(n_0_0_180), .ZN(
      mant_A[15]));
   NOR2_X1 i_0_0_36 (.A1(n_0_45), .A2(n_0_0_180), .ZN(n_0_0_28));
   AOI21_X1 i_0_0_37 (.A(n_0_0_29), .B1(n_0_0_349), .B2(n_0_0_180), .ZN(
      mant_A[16]));
   NOR2_X1 i_0_0_38 (.A1(n_0_46), .A2(n_0_0_180), .ZN(n_0_0_29));
   AOI21_X1 i_0_0_39 (.A(n_0_0_30), .B1(n_0_0_352), .B2(n_0_0_180), .ZN(
      mant_A[17]));
   NOR2_X1 i_0_0_40 (.A1(n_0_47), .A2(n_0_0_180), .ZN(n_0_0_30));
   AOI21_X1 i_0_0_41 (.A(n_0_0_31), .B1(n_0_0_356), .B2(n_0_0_180), .ZN(
      mant_A[18]));
   NOR2_X1 i_0_0_42 (.A1(n_0_48), .A2(n_0_0_180), .ZN(n_0_0_31));
   AOI21_X1 i_0_0_43 (.A(n_0_0_32), .B1(n_0_0_360), .B2(n_0_0_180), .ZN(
      mant_A[19]));
   NOR2_X1 i_0_0_44 (.A1(n_0_49), .A2(n_0_0_180), .ZN(n_0_0_32));
   AOI21_X1 i_0_0_45 (.A(n_0_0_33), .B1(n_0_0_367), .B2(n_0_0_180), .ZN(
      mant_A[20]));
   NOR2_X1 i_0_0_46 (.A1(n_0_50), .A2(n_0_0_180), .ZN(n_0_0_33));
   AOI21_X1 i_0_0_47 (.A(n_0_0_34), .B1(n_0_0_370), .B2(n_0_0_180), .ZN(
      mant_A[21]));
   NOR2_X1 i_0_0_48 (.A1(n_0_51), .A2(n_0_0_180), .ZN(n_0_0_34));
   AOI21_X1 i_0_0_49 (.A(n_0_0_35), .B1(n_0_0_373), .B2(n_0_0_180), .ZN(
      mant_A[22]));
   NOR2_X1 i_0_0_50 (.A1(n_0_52), .A2(n_0_0_180), .ZN(n_0_0_35));
   AOI22_X1 i_0_0_51 (.A1(n_0_0_545), .A2(n_0_0_181), .B1(n_0_0_392), .B2(
      n_0_0_214), .ZN(mant_A[23]));
   AND2_X1 i_0_0_52 (.A1(n_0_54), .A2(n_0_0_181), .ZN(mant_A[31]));
   AND2_X1 i_0_0_53 (.A1(n_0_0_214), .A2(n_0_0_154), .ZN(overflow));
   AND2_X1 i_0_0_54 (.A1(n_0_30), .A2(n_0_0_179), .ZN(underflow));
   INV_X1 i_0_0_55 (.A(n_0_0_36), .ZN(Sum[0]));
   AOI22_X1 i_0_0_56 (.A1(n_0_5), .A2(n_0_0_42), .B1(n_0_6), .B2(n_0_0_153), 
      .ZN(n_0_0_36));
   INV_X1 i_0_0_57 (.A(n_0_0_37), .ZN(Sum[1]));
   AOI221_X1 i_0_0_58 (.A(n_0_0_38), .B1(n_0_7), .B2(n_0_0_153), .C1(n_0_6), 
      .C2(n_0_0_42), .ZN(n_0_0_37));
   AND3_X1 i_0_0_59 (.A1(n_0_0_150), .A2(n_0_0_49), .A3(n_0_5), .ZN(n_0_0_38));
   NAND2_X1 i_0_0_60 (.A1(n_0_0_41), .A2(n_0_0_39), .ZN(Sum[2]));
   AOI21_X1 i_0_0_61 (.A(n_0_0_40), .B1(n_0_7), .B2(n_0_0_42), .ZN(n_0_0_39));
   AND3_X1 i_0_0_62 (.A1(n_0_0_150), .A2(n_0_0_49), .A3(n_0_6), .ZN(n_0_0_40));
   AOI22_X1 i_0_0_63 (.A1(n_0_8), .A2(n_0_0_153), .B1(n_0_0_135), .B2(n_0_0_45), 
      .ZN(n_0_0_41));
   INV_X1 i_0_0_64 (.A(n_0_0_43), .ZN(n_0_0_42));
   AOI21_X1 i_0_0_65 (.A(n_0_0_157), .B1(n_0_0_135), .B2(n_0_0_49), .ZN(n_0_0_43));
   OAI221_X1 i_0_0_66 (.A(n_0_0_46), .B1(n_0_0_151), .B2(n_0_0_44), .C1(
      n_0_0_134), .C2(n_0_0_48), .ZN(Sum[3]));
   AOI21_X1 i_0_0_67 (.A(n_0_0_45), .B1(n_0_7), .B2(n_0_0_49), .ZN(n_0_0_44));
   AND2_X1 i_0_0_68 (.A1(n_0_5), .A2(n_0_0_58), .ZN(n_0_0_45));
   AOI22_X1 i_0_0_69 (.A1(n_0_8), .A2(n_0_0_157), .B1(n_0_9), .B2(n_0_0_153), 
      .ZN(n_0_0_46));
   OAI211_X1 i_0_0_70 (.A(n_0_0_50), .B(n_0_0_47), .C1(n_0_0_151), .C2(n_0_0_48), 
      .ZN(Sum[4]));
   NAND2_X1 i_0_0_71 (.A1(n_0_9), .A2(n_0_0_157), .ZN(n_0_0_47));
   AOI22_X1 i_0_0_72 (.A1(n_0_6), .A2(n_0_0_58), .B1(n_0_8), .B2(n_0_0_49), 
      .ZN(n_0_0_48));
   AND2_X1 i_0_0_73 (.A1(n_0_0_547), .A2(n_0_0_141), .ZN(n_0_0_49));
   AOI22_X1 i_0_0_74 (.A1(n_0_0_135), .A2(n_0_0_52), .B1(n_0_10), .B2(n_0_0_153), 
      .ZN(n_0_0_50));
   NAND2_X1 i_0_0_75 (.A1(n_0_0_54), .A2(n_0_0_51), .ZN(Sum[5]));
   AOI22_X1 i_0_0_76 (.A1(n_0_0_150), .A2(n_0_0_52), .B1(n_0_10), .B2(n_0_0_157), 
      .ZN(n_0_0_51));
   OAI21_X1 i_0_0_77 (.A(n_0_0_53), .B1(n_0_1), .B2(n_0_0_62), .ZN(n_0_0_52));
   NAND2_X1 i_0_0_78 (.A1(n_0_7), .A2(n_0_0_58), .ZN(n_0_0_53));
   AOI22_X1 i_0_0_79 (.A1(n_0_0_135), .A2(n_0_0_56), .B1(n_0_11), .B2(n_0_0_153), 
      .ZN(n_0_0_54));
   NAND2_X1 i_0_0_80 (.A1(n_0_0_59), .A2(n_0_0_55), .ZN(Sum[6]));
   AOI22_X1 i_0_0_81 (.A1(n_0_0_135), .A2(n_0_0_61), .B1(n_0_0_150), .B2(
      n_0_0_56), .ZN(n_0_0_55));
   OAI21_X1 i_0_0_82 (.A(n_0_0_57), .B1(n_0_1), .B2(n_0_0_66), .ZN(n_0_0_56));
   NAND2_X1 i_0_0_83 (.A1(n_0_8), .A2(n_0_0_58), .ZN(n_0_0_57));
   AND2_X1 i_0_0_84 (.A1(n_0_1), .A2(n_0_0_141), .ZN(n_0_0_58));
   AOI22_X1 i_0_0_85 (.A1(n_0_12), .A2(n_0_0_153), .B1(n_0_11), .B2(n_0_0_157), 
      .ZN(n_0_0_59));
   NAND2_X1 i_0_0_86 (.A1(n_0_0_63), .A2(n_0_0_60), .ZN(Sum[7]));
   AOI22_X1 i_0_0_87 (.A1(n_0_0_150), .A2(n_0_0_61), .B1(n_0_12), .B2(n_0_0_157), 
      .ZN(n_0_0_60));
   OAI22_X1 i_0_0_88 (.A1(n_0_1), .A2(n_0_0_70), .B1(n_0_0_547), .B2(n_0_0_62), 
      .ZN(n_0_0_61));
   AOI22_X1 i_0_0_89 (.A1(n_0_9), .A2(n_0_0_141), .B1(n_0_5), .B2(n_0_0_108), 
      .ZN(n_0_0_62));
   AOI22_X1 i_0_0_90 (.A1(n_0_0_135), .A2(n_0_0_65), .B1(n_0_13), .B2(n_0_0_153), 
      .ZN(n_0_0_63));
   NAND2_X1 i_0_0_91 (.A1(n_0_0_67), .A2(n_0_0_64), .ZN(Sum[8]));
   AOI22_X1 i_0_0_92 (.A1(n_0_0_150), .A2(n_0_0_65), .B1(n_0_13), .B2(n_0_0_157), 
      .ZN(n_0_0_64));
   OAI22_X1 i_0_0_93 (.A1(n_0_1), .A2(n_0_0_74), .B1(n_0_0_547), .B2(n_0_0_66), 
      .ZN(n_0_0_65));
   AOI22_X1 i_0_0_94 (.A1(n_0_10), .A2(n_0_0_141), .B1(n_0_6), .B2(n_0_0_108), 
      .ZN(n_0_0_66));
   AOI22_X1 i_0_0_95 (.A1(n_0_14), .A2(n_0_0_153), .B1(n_0_0_135), .B2(n_0_0_69), 
      .ZN(n_0_0_67));
   NAND2_X1 i_0_0_96 (.A1(n_0_0_71), .A2(n_0_0_68), .ZN(Sum[9]));
   AOI22_X1 i_0_0_97 (.A1(n_0_14), .A2(n_0_0_157), .B1(n_0_0_150), .B2(n_0_0_69), 
      .ZN(n_0_0_68));
   OAI22_X1 i_0_0_98 (.A1(n_0_1), .A2(n_0_0_78), .B1(n_0_0_547), .B2(n_0_0_70), 
      .ZN(n_0_0_69));
   AOI22_X1 i_0_0_99 (.A1(n_0_11), .A2(n_0_0_141), .B1(n_0_7), .B2(n_0_0_108), 
      .ZN(n_0_0_70));
   AOI22_X1 i_0_0_100 (.A1(n_0_15), .A2(n_0_0_153), .B1(n_0_0_135), .B2(n_0_0_73), 
      .ZN(n_0_0_71));
   NAND2_X1 i_0_0_101 (.A1(n_0_0_75), .A2(n_0_0_72), .ZN(Sum[10]));
   AOI22_X1 i_0_0_102 (.A1(n_0_0_150), .A2(n_0_0_73), .B1(n_0_15), .B2(n_0_0_157), 
      .ZN(n_0_0_72));
   OAI22_X1 i_0_0_103 (.A1(n_0_1), .A2(n_0_0_82), .B1(n_0_0_547), .B2(n_0_0_74), 
      .ZN(n_0_0_73));
   AOI22_X1 i_0_0_104 (.A1(n_0_12), .A2(n_0_0_141), .B1(n_0_8), .B2(n_0_0_108), 
      .ZN(n_0_0_74));
   AOI22_X1 i_0_0_105 (.A1(n_0_0_135), .A2(n_0_0_77), .B1(n_0_16), .B2(n_0_0_153), 
      .ZN(n_0_0_75));
   NAND2_X1 i_0_0_106 (.A1(n_0_0_79), .A2(n_0_0_76), .ZN(Sum[11]));
   AOI22_X1 i_0_0_107 (.A1(n_0_0_135), .A2(n_0_0_81), .B1(n_0_0_150), .B2(
      n_0_0_77), .ZN(n_0_0_76));
   OAI22_X1 i_0_0_108 (.A1(n_0_1), .A2(n_0_0_87), .B1(n_0_0_547), .B2(n_0_0_78), 
      .ZN(n_0_0_77));
   AOI222_X1 i_0_0_109 (.A1(n_0_5), .A2(n_0_0_143), .B1(n_0_13), .B2(n_0_0_141), 
      .C1(n_0_9), .C2(n_0_0_108), .ZN(n_0_0_78));
   AOI22_X1 i_0_0_110 (.A1(n_0_16), .A2(n_0_0_157), .B1(n_0_17), .B2(n_0_0_153), 
      .ZN(n_0_0_79));
   NAND2_X1 i_0_0_111 (.A1(n_0_0_83), .A2(n_0_0_80), .ZN(Sum[12]));
   AOI22_X1 i_0_0_112 (.A1(n_0_0_150), .A2(n_0_0_81), .B1(n_0_0_135), .B2(
      n_0_0_85), .ZN(n_0_0_80));
   OAI22_X1 i_0_0_113 (.A1(n_0_0_547), .A2(n_0_0_82), .B1(n_0_1), .B2(n_0_0_92), 
      .ZN(n_0_0_81));
   AOI222_X1 i_0_0_114 (.A1(n_0_10), .A2(n_0_0_108), .B1(n_0_6), .B2(n_0_0_143), 
      .C1(n_0_14), .C2(n_0_0_141), .ZN(n_0_0_82));
   AOI22_X1 i_0_0_115 (.A1(n_0_18), .A2(n_0_0_153), .B1(n_0_17), .B2(n_0_0_157), 
      .ZN(n_0_0_83));
   NAND2_X1 i_0_0_116 (.A1(n_0_0_88), .A2(n_0_0_84), .ZN(Sum[13]));
   AOI22_X1 i_0_0_117 (.A1(n_0_0_150), .A2(n_0_0_85), .B1(n_0_0_135), .B2(
      n_0_0_90), .ZN(n_0_0_84));
   OAI21_X1 i_0_0_118 (.A(n_0_0_86), .B1(n_0_0_547), .B2(n_0_0_87), .ZN(n_0_0_85));
   NAND2_X1 i_0_0_119 (.A1(n_0_0_547), .A2(n_0_0_94), .ZN(n_0_0_86));
   AOI222_X1 i_0_0_120 (.A1(n_0_11), .A2(n_0_0_108), .B1(n_0_7), .B2(n_0_0_143), 
      .C1(n_0_15), .C2(n_0_0_141), .ZN(n_0_0_87));
   AOI22_X1 i_0_0_121 (.A1(n_0_19), .A2(n_0_0_153), .B1(n_0_18), .B2(n_0_0_157), 
      .ZN(n_0_0_88));
   OAI21_X1 i_0_0_122 (.A(n_0_0_89), .B1(n_0_0_134), .B2(n_0_0_93), .ZN(Sum[14]));
   AOI222_X1 i_0_0_123 (.A1(n_0_20), .A2(n_0_0_153), .B1(n_0_19), .B2(n_0_0_157), 
      .C1(n_0_0_150), .C2(n_0_0_90), .ZN(n_0_0_89));
   OAI21_X1 i_0_0_124 (.A(n_0_0_91), .B1(n_0_0_547), .B2(n_0_0_92), .ZN(n_0_0_90));
   NAND2_X1 i_0_0_125 (.A1(n_0_0_547), .A2(n_0_0_98), .ZN(n_0_0_91));
   AOI222_X1 i_0_0_126 (.A1(n_0_12), .A2(n_0_0_108), .B1(n_0_8), .B2(n_0_0_143), 
      .C1(n_0_16), .C2(n_0_0_141), .ZN(n_0_0_92));
   OAI221_X1 i_0_0_127 (.A(n_0_0_96), .B1(n_0_0_151), .B2(n_0_0_93), .C1(
      n_0_0_134), .C2(n_0_0_97), .ZN(Sum[15]));
   AOI22_X1 i_0_0_128 (.A1(n_0_0_547), .A2(n_0_0_102), .B1(n_0_1), .B2(n_0_0_94), 
      .ZN(n_0_0_93));
   OAI21_X1 i_0_0_129 (.A(n_0_0_95), .B1(n_0_2), .B2(n_0_0_114), .ZN(n_0_0_94));
   AOI22_X1 i_0_0_130 (.A1(n_0_5), .A2(n_0_0_109), .B1(n_0_13), .B2(n_0_0_108), 
      .ZN(n_0_0_95));
   AOI22_X1 i_0_0_131 (.A1(n_0_20), .A2(n_0_0_157), .B1(n_0_21), .B2(n_0_0_153), 
      .ZN(n_0_0_96));
   OAI221_X1 i_0_0_132 (.A(n_0_0_100), .B1(n_0_0_134), .B2(n_0_0_101), .C1(
      n_0_0_151), .C2(n_0_0_97), .ZN(Sum[16]));
   AOI22_X1 i_0_0_133 (.A1(n_0_1), .A2(n_0_0_98), .B1(n_0_0_547), .B2(n_0_0_106), 
      .ZN(n_0_0_97));
   OAI21_X1 i_0_0_134 (.A(n_0_0_99), .B1(n_0_2), .B2(n_0_0_118), .ZN(n_0_0_98));
   AOI22_X1 i_0_0_135 (.A1(n_0_6), .A2(n_0_0_109), .B1(n_0_14), .B2(n_0_0_108), 
      .ZN(n_0_0_99));
   AOI22_X1 i_0_0_136 (.A1(n_0_21), .A2(n_0_0_157), .B1(n_0_22), .B2(n_0_0_153), 
      .ZN(n_0_0_100));
   OAI221_X1 i_0_0_137 (.A(n_0_0_104), .B1(n_0_0_151), .B2(n_0_0_101), .C1(
      n_0_0_134), .C2(n_0_0_105), .ZN(Sum[17]));
   AOI22_X1 i_0_0_138 (.A1(n_0_0_547), .A2(n_0_0_113), .B1(n_0_1), .B2(n_0_0_102), 
      .ZN(n_0_0_101));
   OAI21_X1 i_0_0_139 (.A(n_0_0_103), .B1(n_0_2), .B2(n_0_0_123), .ZN(n_0_0_102));
   AOI22_X1 i_0_0_140 (.A1(n_0_7), .A2(n_0_0_109), .B1(n_0_15), .B2(n_0_0_108), 
      .ZN(n_0_0_103));
   AOI22_X1 i_0_0_141 (.A1(n_0_22), .A2(n_0_0_157), .B1(n_0_23), .B2(n_0_0_153), 
      .ZN(n_0_0_104));
   OAI221_X1 i_0_0_142 (.A(n_0_0_110), .B1(n_0_0_151), .B2(n_0_0_105), .C1(
      n_0_0_134), .C2(n_0_0_112), .ZN(Sum[18]));
   AOI22_X1 i_0_0_143 (.A1(n_0_1), .A2(n_0_0_106), .B1(n_0_0_547), .B2(n_0_0_117), 
      .ZN(n_0_0_105));
   OAI21_X1 i_0_0_144 (.A(n_0_0_107), .B1(n_0_2), .B2(n_0_0_144), .ZN(n_0_0_106));
   AOI22_X1 i_0_0_145 (.A1(n_0_8), .A2(n_0_0_109), .B1(n_0_16), .B2(n_0_0_108), 
      .ZN(n_0_0_107));
   NOR3_X1 i_0_0_146 (.A1(n_0_4), .A2(n_0_3), .A3(n_0_0_548), .ZN(n_0_0_108));
   NOR3_X1 i_0_0_147 (.A1(n_0_4), .A2(n_0_0_549), .A3(n_0_0_548), .ZN(n_0_0_109));
   AOI22_X1 i_0_0_148 (.A1(n_0_23), .A2(n_0_0_157), .B1(n_0_24), .B2(n_0_0_153), 
      .ZN(n_0_0_110));
   OAI221_X1 i_0_0_149 (.A(n_0_0_111), .B1(n_0_0_151), .B2(n_0_0_112), .C1(
      n_0_0_134), .C2(n_0_0_116), .ZN(Sum[19]));
   AOI22_X1 i_0_0_150 (.A1(n_0_25), .A2(n_0_0_153), .B1(n_0_24), .B2(n_0_0_157), 
      .ZN(n_0_0_111));
   AOI22_X1 i_0_0_151 (.A1(n_0_1), .A2(n_0_0_113), .B1(n_0_0_547), .B2(n_0_0_122), 
      .ZN(n_0_0_112));
   OAI22_X1 i_0_0_152 (.A1(n_0_2), .A2(n_0_0_133), .B1(n_0_0_548), .B2(n_0_0_114), 
      .ZN(n_0_0_113));
   AOI22_X1 i_0_0_153 (.A1(n_0_9), .A2(n_0_0_149), .B1(n_0_17), .B2(n_0_0_148), 
      .ZN(n_0_0_114));
   OAI21_X1 i_0_0_154 (.A(n_0_0_115), .B1(n_0_0_151), .B2(n_0_0_116), .ZN(
      Sum[20]));
   AOI222_X1 i_0_0_155 (.A1(n_0_26), .A2(n_0_0_153), .B1(n_0_0_135), .B2(
      n_0_0_120), .C1(n_0_25), .C2(n_0_0_157), .ZN(n_0_0_115));
   AOI22_X1 i_0_0_156 (.A1(n_0_1), .A2(n_0_0_117), .B1(n_0_0_547), .B2(n_0_0_138), 
      .ZN(n_0_0_116));
   OAI22_X1 i_0_0_157 (.A1(n_0_0_548), .A2(n_0_0_118), .B1(n_0_2), .B2(n_0_0_145), 
      .ZN(n_0_0_117));
   AOI22_X1 i_0_0_158 (.A1(n_0_10), .A2(n_0_0_149), .B1(n_0_18), .B2(n_0_0_148), 
      .ZN(n_0_0_118));
   OAI21_X1 i_0_0_159 (.A(n_0_0_119), .B1(n_0_0_136), .B2(n_0_0_134), .ZN(
      Sum[21]));
   AOI222_X1 i_0_0_160 (.A1(n_0_27), .A2(n_0_0_153), .B1(n_0_26), .B2(n_0_0_157), 
      .C1(n_0_0_150), .C2(n_0_0_120), .ZN(n_0_0_119));
   OAI21_X1 i_0_0_161 (.A(n_0_0_121), .B1(n_0_1), .B2(n_0_0_130), .ZN(n_0_0_120));
   NAND2_X1 i_0_0_162 (.A1(n_0_1), .A2(n_0_0_122), .ZN(n_0_0_121));
   OAI22_X1 i_0_0_163 (.A1(n_0_0_548), .A2(n_0_0_123), .B1(n_0_2), .B2(n_0_0_129), 
      .ZN(n_0_0_122));
   AOI22_X1 i_0_0_164 (.A1(n_0_11), .A2(n_0_0_149), .B1(n_0_19), .B2(n_0_0_148), 
      .ZN(n_0_0_123));
   OAI211_X1 i_0_0_165 (.A(n_0_0_152), .B(n_0_0_124), .C1(n_0_0_151), .C2(
      n_0_0_136), .ZN(Sum[22]));
   NAND2_X1 i_0_0_166 (.A1(n_0_0_135), .A2(n_0_0_125), .ZN(n_0_0_124));
   AOI22_X1 i_0_0_167 (.A1(n_0_1), .A2(n_0_0_130), .B1(n_0_0_547), .B2(n_0_0_126), 
      .ZN(n_0_0_125));
   AOI21_X1 i_0_0_168 (.A(n_0_0_127), .B1(n_0_27), .B2(n_0_0_141), .ZN(n_0_0_126));
   OAI21_X1 i_0_0_169 (.A(n_0_0_128), .B1(n_0_0_548), .B2(n_0_0_129), .ZN(
      n_0_0_127));
   AOI22_X1 i_0_0_170 (.A1(n_0_19), .A2(n_0_0_143), .B1(n_0_11), .B2(n_0_0_140), 
      .ZN(n_0_0_128));
   AOI222_X1 i_0_0_171 (.A1(n_0_15), .A2(n_0_0_149), .B1(n_0_7), .B2(n_0_0_147), 
      .C1(n_0_23), .C2(n_0_0_148), .ZN(n_0_0_129));
   AOI21_X1 i_0_0_172 (.A(n_0_0_131), .B1(n_0_9), .B2(n_0_0_140), .ZN(n_0_0_130));
   OAI21_X1 i_0_0_173 (.A(n_0_0_132), .B1(n_0_0_548), .B2(n_0_0_133), .ZN(
      n_0_0_131));
   AOI22_X1 i_0_0_174 (.A1(n_0_25), .A2(n_0_0_141), .B1(n_0_17), .B2(n_0_0_143), 
      .ZN(n_0_0_132));
   AOI222_X1 i_0_0_175 (.A1(n_0_21), .A2(n_0_0_148), .B1(n_0_5), .B2(n_0_0_147), 
      .C1(n_0_13), .C2(n_0_0_149), .ZN(n_0_0_133));
   INV_X1 i_0_0_176 (.A(n_0_0_135), .ZN(n_0_0_134));
   NOR2_X1 i_0_0_177 (.A1(n_0_0), .A2(n_0_0_178), .ZN(n_0_0_135));
   AOI21_X1 i_0_0_178 (.A(n_0_0_137), .B1(n_0_1), .B2(n_0_0_138), .ZN(n_0_0_136));
   AOI221_X1 i_0_0_179 (.A(n_0_1), .B1(n_0_0_548), .B2(n_0_0_146), .C1(n_0_2), 
      .C2(n_0_0_145), .ZN(n_0_0_137));
   OAI211_X1 i_0_0_180 (.A(n_0_0_142), .B(n_0_0_139), .C1(n_0_0_548), .C2(
      n_0_0_144), .ZN(n_0_0_138));
   AOI22_X1 i_0_0_181 (.A1(n_0_24), .A2(n_0_0_141), .B1(n_0_8), .B2(n_0_0_140), 
      .ZN(n_0_0_139));
   AND2_X1 i_0_0_182 (.A1(n_0_0_548), .A2(n_0_0_147), .ZN(n_0_0_140));
   NOR3_X1 i_0_0_183 (.A1(n_0_4), .A2(n_0_3), .A3(n_0_2), .ZN(n_0_0_141));
   NAND2_X1 i_0_0_184 (.A1(n_0_16), .A2(n_0_0_143), .ZN(n_0_0_142));
   NOR3_X1 i_0_0_185 (.A1(n_0_4), .A2(n_0_0_549), .A3(n_0_2), .ZN(n_0_0_143));
   AOI22_X1 i_0_0_186 (.A1(n_0_12), .A2(n_0_0_149), .B1(n_0_20), .B2(n_0_0_148), 
      .ZN(n_0_0_144));
   AOI222_X1 i_0_0_187 (.A1(n_0_14), .A2(n_0_0_149), .B1(n_0_6), .B2(n_0_0_147), 
      .C1(n_0_22), .C2(n_0_0_148), .ZN(n_0_0_145));
   AOI222_X1 i_0_0_188 (.A1(n_0_18), .A2(n_0_0_149), .B1(n_0_10), .B2(n_0_0_147), 
      .C1(n_0_26), .C2(n_0_0_148), .ZN(n_0_0_146));
   NOR2_X1 i_0_0_189 (.A1(n_0_0_550), .A2(n_0_3), .ZN(n_0_0_147));
   NOR2_X1 i_0_0_190 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_0_148));
   NOR2_X1 i_0_0_191 (.A1(n_0_4), .A2(n_0_0_549), .ZN(n_0_0_149));
   INV_X1 i_0_0_192 (.A(n_0_0_151), .ZN(n_0_0_150));
   NAND2_X1 i_0_0_193 (.A1(n_0_0), .A2(n_0_0_179), .ZN(n_0_0_151));
   AOI22_X1 i_0_0_194 (.A1(n_0_27), .A2(n_0_0_157), .B1(n_0_28), .B2(n_0_0_153), 
      .ZN(n_0_0_152));
   NOR3_X1 i_0_0_195 (.A1(n_0_0_546), .A2(n_0_0_213), .A3(n_0_0_154), .ZN(
      n_0_0_153));
   NOR4_X1 i_0_0_196 (.A1(n_0_0_546), .A2(n_0_0_543), .A3(n_0_0_267), .A4(
      n_0_0_155), .ZN(n_0_0_154));
   NAND3_X1 i_0_0_197 (.A1(exp_Sum[5]), .A2(exp_Sum[4]), .A3(n_0_0_156), 
      .ZN(n_0_0_155));
   NOR4_X1 i_0_0_198 (.A1(n_0_0_264), .A2(n_0_0_263), .A3(n_0_0_262), .A4(
      exp_Sum[0]), .ZN(n_0_0_156));
   INV_X1 i_0_0_199 (.A(n_0_0_158), .ZN(n_0_0_157));
   AOI21_X1 i_0_0_200 (.A(n_0_0_174), .B1(n_0_0_546), .B2(n_0_0_214), .ZN(
      n_0_0_158));
   INV_X1 i_0_0_201 (.A(n_0_0_159), .ZN(Sum[23]));
   AOI222_X1 i_0_0_202 (.A1(exp_Sum[0]), .A2(n_0_0_174), .B1(n_0_0_7), .B2(
      n_0_0_214), .C1(n_0_0_177), .C2(n_0_0_160), .ZN(n_0_0_159));
   OAI21_X1 i_0_0_203 (.A(n_0_0_224), .B1(n_0_0), .B2(n_0_0_261), .ZN(n_0_0_160));
   INV_X1 i_0_0_204 (.A(n_0_0_161), .ZN(Sum[24]));
   AOI222_X1 i_0_0_205 (.A1(exp_Sum[1]), .A2(n_0_0_174), .B1(n_0_0_8), .B2(
      n_0_0_214), .C1(n_0_0_177), .C2(n_0_0_162), .ZN(n_0_0_161));
   XOR2_X1 i_0_0_206 (.A(n_0_0_224), .B(n_0_0_222), .Z(n_0_0_162));
   INV_X1 i_0_0_207 (.A(n_0_0_163), .ZN(Sum[25]));
   AOI222_X1 i_0_0_208 (.A1(exp_Sum[2]), .A2(n_0_0_174), .B1(n_0_0_9), .B2(
      n_0_0_214), .C1(n_0_0_177), .C2(n_0_0_164), .ZN(n_0_0_163));
   XOR2_X1 i_0_0_209 (.A(n_0_0_226), .B(n_0_0_221), .Z(n_0_0_164));
   INV_X1 i_0_0_210 (.A(n_0_0_165), .ZN(Sum[26]));
   AOI222_X1 i_0_0_211 (.A1(exp_Sum[3]), .A2(n_0_0_174), .B1(n_0_0_10), .B2(
      n_0_0_214), .C1(n_0_0_177), .C2(n_0_0_166), .ZN(n_0_0_165));
   XNOR2_X1 i_0_0_212 (.A(n_0_0_227), .B(n_0_0_220), .ZN(n_0_0_166));
   INV_X1 i_0_0_213 (.A(n_0_0_167), .ZN(Sum[27]));
   AOI222_X1 i_0_0_214 (.A1(n_0_0_11), .A2(n_0_0_214), .B1(exp_Sum[4]), .B2(
      n_0_0_174), .C1(n_0_0_177), .C2(n_0_0_168), .ZN(n_0_0_167));
   XOR2_X1 i_0_0_215 (.A(n_0_0_228), .B(n_0_0_219), .Z(n_0_0_168));
   INV_X1 i_0_0_216 (.A(n_0_0_169), .ZN(Sum[28]));
   AOI222_X1 i_0_0_217 (.A1(n_0_0_12), .A2(n_0_0_214), .B1(n_0_0_177), .B2(
      n_0_0_170), .C1(exp_Sum[5]), .C2(n_0_0_174), .ZN(n_0_0_169));
   OAI21_X1 i_0_0_218 (.A(n_0_0_217), .B1(n_0_0_266), .B2(n_0_0_218), .ZN(
      n_0_0_170));
   OAI211_X1 i_0_0_219 (.A(n_0_0_176), .B(n_0_0_171), .C1(n_0_0_267), .C2(
      n_0_0_172), .ZN(Sum[29]));
   NAND2_X1 i_0_0_220 (.A1(n_0_0_13), .A2(n_0_0_214), .ZN(n_0_0_171));
   AOI21_X1 i_0_0_221 (.A(n_0_0_174), .B1(n_0_0_217), .B2(n_0_0_177), .ZN(
      n_0_0_172));
   AOI22_X1 i_0_0_222 (.A1(n_0_0_176), .A2(n_0_0_175), .B1(exp_Sum[7]), .B2(
      n_0_0_173), .ZN(Sum[30]));
   AOI221_X1 i_0_0_223 (.A(n_0_0_174), .B1(n_0_0_215), .B2(n_0_0_177), .C1(
      n_0_0_544), .C2(n_0_0_214), .ZN(n_0_0_173));
   AND3_X1 i_0_0_224 (.A1(num_leading_zeros[4]), .A2(num_leading_zeros[3]), 
      .A3(n_0_0_181), .ZN(n_0_0_174));
   AOI21_X1 i_0_0_225 (.A(exp_Sum[7]), .B1(n_0_0_6), .B2(n_0_0_214), .ZN(
      n_0_0_175));
   NAND2_X1 i_0_0_226 (.A1(n_0_0_216), .A2(n_0_0_177), .ZN(n_0_0_176));
   NOR2_X1 i_0_0_227 (.A1(n_0_30), .A2(n_0_0_178), .ZN(n_0_0_177));
   INV_X1 i_0_0_228 (.A(n_0_0_179), .ZN(n_0_0_178));
   AOI21_X1 i_0_0_229 (.A(n_0_0_180), .B1(num_leading_zeros[4]), .B2(
      num_leading_zeros[3]), .ZN(n_0_0_179));
   INV_X1 i_0_0_230 (.A(n_0_0_181), .ZN(n_0_0_180));
   AOI21_X1 i_0_0_231 (.A(n_0_0_214), .B1(n_0_0_194), .B2(n_0_0_182), .ZN(
      n_0_0_181));
   NOR4_X1 i_0_0_232 (.A1(n_0_0_187), .A2(n_0_0_186), .A3(n_0_0_188), .A4(
      n_0_0_183), .ZN(n_0_0_182));
   NAND4_X1 i_0_0_233 (.A1(n_0_0_185), .A2(n_0_0_184), .A3(n_0_0_211), .A4(
      n_0_0_202), .ZN(n_0_0_183));
   AOI21_X1 i_0_0_234 (.A(n_0_0_203), .B1(n_0_0_412), .B2(n_0_59), .ZN(n_0_0_184));
   AOI22_X1 i_0_0_235 (.A1(n_0_0_402), .A2(n_0_57), .B1(n_0_79), .B2(n_0_0_268), 
      .ZN(n_0_0_185));
   AOI22_X1 i_0_0_236 (.A1(n_0_0_456), .A2(n_0_0_341), .B1(n_0_94), .B2(n_0_70), 
      .ZN(n_0_0_186));
   OAI221_X1 i_0_0_237 (.A(n_0_0_208), .B1(n_0_97), .B2(n_0_0_356), .C1(n_0_84), 
      .C2(n_0_0_293), .ZN(n_0_0_187));
   NAND4_X1 i_0_0_238 (.A1(n_0_0_207), .A2(n_0_0_189), .A3(n_0_0_192), .A4(
      n_0_0_212), .ZN(n_0_0_188));
   INV_X1 i_0_0_239 (.A(n_0_0_190), .ZN(n_0_0_189));
   OAI211_X1 i_0_0_240 (.A(n_0_0_506), .B(n_0_0_191), .C1(n_0_100), .C2(
      n_0_0_370), .ZN(n_0_0_190));
   AOI221_X1 i_0_0_241 (.A(n_0_0_391), .B1(n_0_0_485), .B2(n_0_77), .C1(n_0_100), 
      .C2(n_0_0_370), .ZN(n_0_0_191));
   NOR3_X1 i_0_0_242 (.A1(n_0_0_206), .A2(n_0_0_193), .A3(n_0_0_210), .ZN(
      n_0_0_192));
   XOR2_X1 i_0_0_243 (.A(n_0_98), .B(n_0_74), .Z(n_0_0_193));
   NOR4_X1 i_0_0_244 (.A1(n_0_0_204), .A2(n_0_0_200), .A3(n_0_0_205), .A4(
      n_0_0_195), .ZN(n_0_0_194));
   NAND4_X1 i_0_0_245 (.A1(n_0_0_199), .A2(n_0_0_198), .A3(n_0_0_197), .A4(
      n_0_0_196), .ZN(n_0_0_195));
   AOI222_X1 i_0_0_246 (.A1(n_0_0_587), .A2(n_0_67), .B1(B[12]), .B2(n_0_0_329), 
      .C1(n_0_83), .C2(n_0_0_288), .ZN(n_0_0_196));
   AOI22_X1 i_0_0_247 (.A1(n_0_81), .A2(n_0_0_277), .B1(n_0_84), .B2(n_0_0_293), 
      .ZN(n_0_0_197));
   AOI221_X1 i_0_0_248 (.A(n_0_0_209), .B1(n_0_0_452), .B2(n_0_69), .C1(n_0_93), 
      .C2(n_0_0_337), .ZN(n_0_0_198));
   AOI22_X1 i_0_0_249 (.A1(n_0_80), .A2(n_0_0_273), .B1(n_0_0_397), .B2(n_0_56), 
      .ZN(n_0_0_199));
   OAI221_X1 i_0_0_250 (.A(n_0_0_201), .B1(n_0_0_443), .B2(n_0_66), .C1(n_0_89), 
      .C2(n_0_0_317), .ZN(n_0_0_200));
   AOI22_X1 i_0_0_251 (.A1(n_0_0_443), .A2(n_0_66), .B1(n_0_89), .B2(n_0_0_317), 
      .ZN(n_0_0_201));
   NAND2_X1 i_0_0_252 (.A1(n_0_0_393), .A2(n_0_55), .ZN(n_0_0_202));
   AOI22_X1 i_0_0_253 (.A1(n_0_86), .A2(n_0_62), .B1(n_0_0_428), .B2(n_0_0_304), 
      .ZN(n_0_0_203));
   AOI22_X1 i_0_0_254 (.A1(n_0_87), .A2(n_0_63), .B1(n_0_0_434), .B2(n_0_0_308), 
      .ZN(n_0_0_204));
   AOI22_X1 i_0_0_255 (.A1(n_0_92), .A2(n_0_68), .B1(n_0_0_449), .B2(n_0_0_332), 
      .ZN(n_0_0_205));
   OAI222_X1 i_0_0_256 (.A1(n_0_99), .A2(n_0_0_367), .B1(n_0_0_474), .B2(n_0_75), 
      .C1(n_0_0_485), .C2(n_0_77), .ZN(n_0_0_206));
   XNOR2_X1 i_0_0_257 (.A(n_0_95), .B(n_0_71), .ZN(n_0_0_207));
   NAND2_X1 i_0_0_258 (.A1(n_0_97), .A2(n_0_0_356), .ZN(n_0_0_208));
   AOI22_X1 i_0_0_259 (.A1(n_0_85), .A2(n_0_61), .B1(n_0_0_422), .B2(n_0_0_298), 
      .ZN(n_0_0_209));
   XNOR2_X1 i_0_0_260 (.A(n_0_96), .B(n_0_0_352), .ZN(n_0_0_210));
   AOI22_X1 i_0_0_261 (.A1(n_0_0_406), .A2(n_0_58), .B1(n_0_82), .B2(n_0_0_282), 
      .ZN(n_0_0_211));
   AOI22_X1 i_0_0_262 (.A1(n_0_88), .A2(n_0_0_314), .B1(n_0_0_437), .B2(n_0_64), 
      .ZN(n_0_0_212));
   INV_X1 i_0_0_263 (.A(n_0_0_214), .ZN(n_0_0_213));
   XNOR2_X1 i_0_0_264 (.A(B[31]), .B(A[31]), .ZN(n_0_0_214));
   INV_X1 i_0_0_265 (.A(n_0_0_216), .ZN(n_0_0_215));
   NOR2_X1 i_0_0_266 (.A1(exp_Sum[6]), .A2(n_0_0_217), .ZN(n_0_0_216));
   NAND2_X1 i_0_0_267 (.A1(n_0_0_266), .A2(n_0_0_218), .ZN(n_0_0_217));
   AOI22_X1 i_0_0_268 (.A1(n_0_0_550), .A2(exp_Sum[4]), .B1(n_0_0_228), .B2(
      n_0_0_219), .ZN(n_0_0_218));
   AOI22_X1 i_0_0_269 (.A1(n_0_3), .A2(n_0_0_264), .B1(n_0_0_227), .B2(n_0_0_220), 
      .ZN(n_0_0_219));
   OAI22_X1 i_0_0_270 (.A1(n_0_0_548), .A2(exp_Sum[2]), .B1(n_0_0_225), .B2(
      n_0_0_221), .ZN(n_0_0_220));
   AOI22_X1 i_0_0_271 (.A1(n_0_1), .A2(n_0_0_262), .B1(n_0_0_223), .B2(n_0_0_222), 
      .ZN(n_0_0_221));
   AOI22_X1 i_0_0_272 (.A1(n_0_1), .A2(n_0_0_262), .B1(n_0_0_547), .B2(
      exp_Sum[1]), .ZN(n_0_0_222));
   INV_X1 i_0_0_273 (.A(n_0_0_224), .ZN(n_0_0_223));
   NAND2_X1 i_0_0_274 (.A1(n_0_0), .A2(n_0_0_261), .ZN(n_0_0_224));
   INV_X1 i_0_0_275 (.A(n_0_0_226), .ZN(n_0_0_225));
   AOI22_X1 i_0_0_276 (.A1(n_0_2), .A2(n_0_0_263), .B1(n_0_0_548), .B2(
      exp_Sum[2]), .ZN(n_0_0_226));
   AOI22_X1 i_0_0_277 (.A1(n_0_3), .A2(n_0_0_264), .B1(n_0_0_549), .B2(
      exp_Sum[3]), .ZN(n_0_0_227));
   AOI22_X1 i_0_0_278 (.A1(n_0_0_550), .A2(exp_Sum[4]), .B1(n_0_4), .B2(
      n_0_0_265), .ZN(n_0_0_228));
   OAI21_X1 i_0_0_279 (.A(n_0_0_229), .B1(n_0_0_600), .B2(n_0_0_230), .ZN(
      Sum[31]));
   NAND2_X1 i_0_0_280 (.A1(A[31]), .A2(n_0_0_230), .ZN(n_0_0_229));
   AOI211_X1 i_0_0_281 (.A(n_0_0_392), .B(n_0_0_231), .C1(n_0_0_233), .C2(
      n_0_0_232), .ZN(n_0_0_230));
   NOR3_X1 i_0_0_282 (.A1(n_0_0_595), .A2(n_0_0_513), .A3(A[22]), .ZN(n_0_0_231));
   AOI221_X1 i_0_0_283 (.A(n_0_0_513), .B1(n_0_0_594), .B2(A[21]), .C1(n_0_0_595), 
      .C2(A[22]), .ZN(n_0_0_232));
   INV_X1 i_0_0_284 (.A(n_0_0_234), .ZN(n_0_0_233));
   AOI221_X1 i_0_0_285 (.A(n_0_0_235), .B1(B[21]), .B2(n_0_0_569), .C1(B[20]), 
      .C2(n_0_0_568), .ZN(n_0_0_234));
   AOI221_X1 i_0_0_286 (.A(n_0_0_236), .B1(n_0_0_593), .B2(A[20]), .C1(n_0_0_592), 
      .C2(A[19]), .ZN(n_0_0_235));
   AOI221_X1 i_0_0_287 (.A(n_0_0_237), .B1(B[18]), .B2(n_0_0_566), .C1(B[19]), 
      .C2(n_0_0_567), .ZN(n_0_0_236));
   AOI21_X1 i_0_0_288 (.A(n_0_0_238), .B1(n_0_0_591), .B2(A[18]), .ZN(n_0_0_237));
   AOI22_X1 i_0_0_289 (.A1(n_0_0_240), .A2(n_0_0_239), .B1(B[17]), .B2(n_0_0_565), 
      .ZN(n_0_0_238));
   AOI22_X1 i_0_0_290 (.A1(n_0_0_589), .A2(A[16]), .B1(n_0_0_590), .B2(A[17]), 
      .ZN(n_0_0_239));
   OAI221_X1 i_0_0_291 (.A(n_0_0_241), .B1(n_0_0_589), .B2(A[16]), .C1(n_0_0_588), 
      .C2(A[15]), .ZN(n_0_0_240));
   INV_X1 i_0_0_292 (.A(n_0_0_242), .ZN(n_0_0_241));
   AOI21_X1 i_0_0_293 (.A(n_0_0_243), .B1(n_0_0_588), .B2(A[15]), .ZN(n_0_0_242));
   AOI21_X1 i_0_0_294 (.A(n_0_0_244), .B1(B[14]), .B2(n_0_0_564), .ZN(n_0_0_243));
   NOR2_X1 i_0_0_295 (.A1(n_0_0_246), .A2(n_0_0_245), .ZN(n_0_0_244));
   OAI22_X1 i_0_0_296 (.A1(B[13]), .A2(n_0_0_563), .B1(B[14]), .B2(n_0_0_564), 
      .ZN(n_0_0_245));
   AOI221_X1 i_0_0_297 (.A(n_0_0_247), .B1(B[12]), .B2(n_0_0_562), .C1(B[13]), 
      .C2(n_0_0_563), .ZN(n_0_0_246));
   AOI221_X1 i_0_0_298 (.A(n_0_0_248), .B1(n_0_0_587), .B2(A[12]), .C1(n_0_0_586), 
      .C2(A[11]), .ZN(n_0_0_247));
   AOI221_X1 i_0_0_299 (.A(n_0_0_249), .B1(B[10]), .B2(n_0_0_560), .C1(B[11]), 
      .C2(n_0_0_561), .ZN(n_0_0_248));
   AOI221_X1 i_0_0_300 (.A(n_0_0_250), .B1(n_0_0_585), .B2(A[10]), .C1(n_0_0_584), 
      .C2(A[9]), .ZN(n_0_0_249));
   AOI221_X1 i_0_0_301 (.A(n_0_0_251), .B1(B[8]), .B2(n_0_0_558), .C1(B[9]), 
      .C2(n_0_0_559), .ZN(n_0_0_250));
   AOI21_X1 i_0_0_302 (.A(n_0_0_252), .B1(n_0_0_583), .B2(A[8]), .ZN(n_0_0_251));
   AOI22_X1 i_0_0_303 (.A1(B[7]), .A2(n_0_0_557), .B1(n_0_0_254), .B2(n_0_0_253), 
      .ZN(n_0_0_252));
   AOI22_X1 i_0_0_304 (.A1(n_0_0_582), .A2(A[7]), .B1(n_0_0_581), .B2(A[6]), 
      .ZN(n_0_0_253));
   INV_X1 i_0_0_305 (.A(n_0_0_255), .ZN(n_0_0_254));
   AOI221_X1 i_0_0_306 (.A(n_0_0_256), .B1(B[5]), .B2(n_0_0_555), .C1(B[6]), 
      .C2(n_0_0_556), .ZN(n_0_0_255));
   AOI221_X1 i_0_0_307 (.A(n_0_0_257), .B1(n_0_0_580), .B2(A[5]), .C1(n_0_0_579), 
      .C2(A[4]), .ZN(n_0_0_256));
   AOI221_X1 i_0_0_308 (.A(n_0_0_258), .B1(B[3]), .B2(n_0_0_553), .C1(B[4]), 
      .C2(n_0_0_554), .ZN(n_0_0_257));
   AOI221_X1 i_0_0_309 (.A(n_0_0_259), .B1(n_0_0_577), .B2(A[2]), .C1(n_0_0_578), 
      .C2(A[3]), .ZN(n_0_0_258));
   AOI221_X1 i_0_0_310 (.A(n_0_0_260), .B1(B[1]), .B2(n_0_0_551), .C1(B[2]), 
      .C2(n_0_0_552), .ZN(n_0_0_259));
   AOI22_X1 i_0_0_311 (.A1(n_0_0_576), .A2(A[1]), .B1(n_0_0_575), .B2(A[0]), 
      .ZN(n_0_0_260));
   INV_X1 i_0_0_312 (.A(n_0_0_261), .ZN(exp_Sum[0]));
   AOI22_X1 i_0_0_313 (.A1(B[23]), .A2(n_0_0_392), .B1(A[23]), .B2(n_0_78), 
      .ZN(n_0_0_261));
   INV_X1 i_0_0_314 (.A(n_0_0_262), .ZN(exp_Sum[1]));
   AOI22_X1 i_0_0_315 (.A1(B[24]), .A2(n_0_0_392), .B1(A[24]), .B2(n_0_78), 
      .ZN(n_0_0_262));
   INV_X1 i_0_0_316 (.A(n_0_0_263), .ZN(exp_Sum[2]));
   AOI22_X1 i_0_0_317 (.A1(B[25]), .A2(n_0_0_392), .B1(A[25]), .B2(n_0_78), 
      .ZN(n_0_0_263));
   INV_X1 i_0_0_318 (.A(n_0_0_264), .ZN(exp_Sum[3]));
   AOI22_X1 i_0_0_319 (.A1(A[26]), .A2(n_0_78), .B1(B[26]), .B2(n_0_0_392), 
      .ZN(n_0_0_264));
   INV_X1 i_0_0_320 (.A(n_0_0_265), .ZN(exp_Sum[4]));
   AOI22_X1 i_0_0_321 (.A1(B[27]), .A2(n_0_0_392), .B1(A[27]), .B2(n_0_78), 
      .ZN(n_0_0_265));
   INV_X1 i_0_0_322 (.A(n_0_0_266), .ZN(exp_Sum[5]));
   AOI22_X1 i_0_0_323 (.A1(B[28]), .A2(n_0_0_392), .B1(A[28]), .B2(n_0_78), 
      .ZN(n_0_0_266));
   INV_X1 i_0_0_324 (.A(n_0_0_267), .ZN(exp_Sum[6]));
   AOI22_X1 i_0_0_325 (.A1(B[29]), .A2(n_0_0_392), .B1(A[29]), .B2(n_0_78), 
      .ZN(n_0_0_267));
   INV_X1 i_0_0_326 (.A(n_0_0_268), .ZN(n_0_55));
   AOI221_X1 i_0_0_327 (.A(n_0_0_269), .B1(n_0_0_363), .B2(n_0_0_274), .C1(A[0]), 
      .C2(n_0_78), .ZN(n_0_0_268));
   AOI221_X1 i_0_0_328 (.A(n_0_0_372), .B1(n_0_0_375), .B2(n_0_0_270), .C1(
      n_0_0_376), .C2(n_0_0_279), .ZN(n_0_0_269));
   AOI222_X1 i_0_0_329 (.A1(A[0]), .A2(n_0_0_378), .B1(n_0_0_380), .B2(n_0_0_271), 
      .C1(n_0_0_381), .C2(n_0_0_291), .ZN(n_0_0_270));
   OAI21_X1 i_0_0_330 (.A(n_0_0_272), .B1(n_0_0_558), .B2(n_0_0_348), .ZN(
      n_0_0_271));
   NAND2_X1 i_0_0_331 (.A1(A[16]), .A2(n_0_0_303), .ZN(n_0_0_272));
   INV_X1 i_0_0_332 (.A(n_0_0_273), .ZN(n_0_56));
   AOI222_X1 i_0_0_333 (.A1(A[1]), .A2(n_0_78), .B1(n_0_0_371), .B2(n_0_0_274), 
      .C1(n_0_0_363), .C2(n_0_0_278), .ZN(n_0_0_273));
   AOI22_X1 i_0_0_334 (.A1(n_0_0_376), .A2(n_0_0_284), .B1(n_0_0_276), .B2(
      n_0_0_275), .ZN(n_0_0_274));
   AOI221_X1 i_0_0_335 (.A(n_0_0_376), .B1(A[1]), .B2(n_0_0_378), .C1(A[17]), 
      .C2(n_0_0_287), .ZN(n_0_0_275));
   AOI22_X1 i_0_0_336 (.A1(n_0_0_381), .A2(n_0_0_296), .B1(A[9]), .B2(n_0_0_340), 
      .ZN(n_0_0_276));
   INV_X1 i_0_0_337 (.A(n_0_0_277), .ZN(n_0_57));
   AOI222_X1 i_0_0_338 (.A1(n_0_0_363), .A2(n_0_0_283), .B1(A[2]), .B2(n_0_78), 
      .C1(n_0_0_371), .C2(n_0_0_278), .ZN(n_0_0_277));
   AOI22_X1 i_0_0_339 (.A1(n_0_0_375), .A2(n_0_0_279), .B1(n_0_0_376), .B2(
      n_0_0_290), .ZN(n_0_0_278));
   AOI221_X1 i_0_0_340 (.A(n_0_0_280), .B1(A[18]), .B2(n_0_0_287), .C1(A[2]), 
      .C2(n_0_0_378), .ZN(n_0_0_279));
   INV_X1 i_0_0_341 (.A(n_0_0_281), .ZN(n_0_0_280));
   AOI22_X1 i_0_0_342 (.A1(n_0_0_381), .A2(n_0_0_301), .B1(A[10]), .B2(n_0_0_340), 
      .ZN(n_0_0_281));
   INV_X1 i_0_0_343 (.A(n_0_0_282), .ZN(n_0_58));
   AOI222_X1 i_0_0_344 (.A1(n_0_0_363), .A2(n_0_0_289), .B1(A[3]), .B2(n_0_78), 
      .C1(n_0_0_371), .C2(n_0_0_283), .ZN(n_0_0_282));
   AOI22_X1 i_0_0_345 (.A1(n_0_0_375), .A2(n_0_0_284), .B1(n_0_0_376), .B2(
      n_0_0_295), .ZN(n_0_0_283));
   AOI221_X1 i_0_0_346 (.A(n_0_0_285), .B1(A[3]), .B2(n_0_0_378), .C1(A[19]), 
      .C2(n_0_0_287), .ZN(n_0_0_284));
   INV_X1 i_0_0_347 (.A(n_0_0_286), .ZN(n_0_0_285));
   AOI22_X1 i_0_0_348 (.A1(n_0_0_381), .A2(n_0_0_307), .B1(A[11]), .B2(n_0_0_340), 
      .ZN(n_0_0_286));
   NOR3_X1 i_0_0_349 (.A1(n_0_0_386), .A2(n_0_0_384), .A3(n_0_0_381), .ZN(
      n_0_0_287));
   INV_X1 i_0_0_350 (.A(n_0_0_288), .ZN(n_0_59));
   AOI222_X1 i_0_0_351 (.A1(n_0_0_363), .A2(n_0_0_294), .B1(A[4]), .B2(n_0_78), 
      .C1(n_0_0_371), .C2(n_0_0_289), .ZN(n_0_0_288));
   AOI22_X1 i_0_0_352 (.A1(n_0_0_375), .A2(n_0_0_290), .B1(n_0_0_376), .B2(
      n_0_0_300), .ZN(n_0_0_289));
   AOI222_X1 i_0_0_353 (.A1(A[8]), .A2(n_0_0_359), .B1(A[16]), .B2(n_0_0_323), 
      .C1(n_0_0_380), .C2(n_0_0_291), .ZN(n_0_0_290));
   OAI21_X1 i_0_0_354 (.A(n_0_0_292), .B1(n_0_0_562), .B2(n_0_0_348), .ZN(
      n_0_0_291));
   AOI22_X1 i_0_0_355 (.A1(A[20]), .A2(n_0_0_303), .B1(A[4]), .B2(n_0_0_382), 
      .ZN(n_0_0_292));
   INV_X1 i_0_0_356 (.A(n_0_0_293), .ZN(n_0_60));
   AOI222_X1 i_0_0_357 (.A1(n_0_0_371), .A2(n_0_0_294), .B1(A[5]), .B2(n_0_78), 
      .C1(n_0_0_363), .C2(n_0_0_299), .ZN(n_0_0_293));
   AOI22_X1 i_0_0_358 (.A1(n_0_0_375), .A2(n_0_0_295), .B1(n_0_0_376), .B2(
      n_0_0_306), .ZN(n_0_0_294));
   AOI222_X1 i_0_0_359 (.A1(A[9]), .A2(n_0_0_359), .B1(A[17]), .B2(n_0_0_323), 
      .C1(n_0_0_380), .C2(n_0_0_296), .ZN(n_0_0_295));
   OAI21_X1 i_0_0_360 (.A(n_0_0_297), .B1(n_0_0_555), .B2(n_0_0_383), .ZN(
      n_0_0_296));
   AOI22_X1 i_0_0_361 (.A1(A[13]), .A2(n_0_0_347), .B1(A[21]), .B2(n_0_0_303), 
      .ZN(n_0_0_297));
   INV_X1 i_0_0_362 (.A(n_0_0_298), .ZN(n_0_61));
   AOI222_X1 i_0_0_363 (.A1(n_0_0_363), .A2(n_0_0_305), .B1(A[6]), .B2(n_0_78), 
      .C1(n_0_0_371), .C2(n_0_0_299), .ZN(n_0_0_298));
   AOI22_X1 i_0_0_364 (.A1(n_0_0_375), .A2(n_0_0_300), .B1(n_0_0_376), .B2(
      n_0_0_311), .ZN(n_0_0_299));
   AOI222_X1 i_0_0_365 (.A1(A[18]), .A2(n_0_0_323), .B1(A[10]), .B2(n_0_0_359), 
      .C1(n_0_0_380), .C2(n_0_0_301), .ZN(n_0_0_300));
   OAI21_X1 i_0_0_366 (.A(n_0_0_302), .B1(n_0_0_556), .B2(n_0_0_383), .ZN(
      n_0_0_301));
   AOI22_X1 i_0_0_367 (.A1(A[14]), .A2(n_0_0_347), .B1(A[22]), .B2(n_0_0_303), 
      .ZN(n_0_0_302));
   NOR2_X1 i_0_0_368 (.A1(n_0_0_386), .A2(n_0_0_384), .ZN(n_0_0_303));
   INV_X1 i_0_0_369 (.A(n_0_0_304), .ZN(n_0_62));
   AOI222_X1 i_0_0_370 (.A1(n_0_0_371), .A2(n_0_0_305), .B1(A[7]), .B2(n_0_78), 
      .C1(n_0_0_363), .C2(n_0_0_309), .ZN(n_0_0_304));
   AOI22_X1 i_0_0_371 (.A1(n_0_0_375), .A2(n_0_0_306), .B1(n_0_0_376), .B2(
      n_0_0_316), .ZN(n_0_0_305));
   AOI22_X1 i_0_0_372 (.A1(n_0_0_380), .A2(n_0_0_307), .B1(n_0_0_381), .B2(
      n_0_0_328), .ZN(n_0_0_306));
   AOI22_X1 i_0_0_373 (.A1(n_0_0_557), .A2(n_0_0_382), .B1(n_0_0_384), .B2(
      n_0_0_346), .ZN(n_0_0_307));
   INV_X1 i_0_0_374 (.A(n_0_0_308), .ZN(n_0_63));
   AOI222_X1 i_0_0_375 (.A1(n_0_0_371), .A2(n_0_0_309), .B1(A[8]), .B2(n_0_78), 
      .C1(n_0_0_363), .C2(n_0_0_315), .ZN(n_0_0_308));
   OAI21_X1 i_0_0_376 (.A(n_0_0_310), .B1(n_0_0_376), .B2(n_0_0_311), .ZN(
      n_0_0_309));
   NAND2_X1 i_0_0_377 (.A1(n_0_0_376), .A2(n_0_0_320), .ZN(n_0_0_310));
   AOI221_X1 i_0_0_378 (.A(n_0_0_312), .B1(A[16]), .B2(n_0_0_340), .C1(A[20]), 
      .C2(n_0_0_323), .ZN(n_0_0_311));
   OAI21_X1 i_0_0_379 (.A(n_0_0_313), .B1(n_0_0_558), .B2(n_0_0_379), .ZN(
      n_0_0_312));
   NAND2_X1 i_0_0_380 (.A1(A[12]), .A2(n_0_0_359), .ZN(n_0_0_313));
   INV_X1 i_0_0_381 (.A(n_0_0_314), .ZN(n_0_64));
   AOI222_X1 i_0_0_382 (.A1(n_0_0_363), .A2(n_0_0_318), .B1(A[9]), .B2(n_0_78), 
      .C1(n_0_0_371), .C2(n_0_0_315), .ZN(n_0_0_314));
   AOI22_X1 i_0_0_383 (.A1(n_0_0_375), .A2(n_0_0_316), .B1(n_0_0_376), .B2(
      n_0_0_327), .ZN(n_0_0_315));
   AOI222_X1 i_0_0_384 (.A1(A[9]), .A2(n_0_0_378), .B1(n_0_0_354), .B2(n_0_0_347), 
      .C1(A[13]), .C2(n_0_0_359), .ZN(n_0_0_316));
   INV_X1 i_0_0_385 (.A(n_0_0_317), .ZN(n_0_65));
   AOI222_X1 i_0_0_386 (.A1(n_0_0_371), .A2(n_0_0_318), .B1(A[10]), .B2(n_0_78), 
      .C1(n_0_0_363), .C2(n_0_0_325), .ZN(n_0_0_317));
   AOI21_X1 i_0_0_387 (.A(n_0_0_319), .B1(n_0_0_376), .B2(n_0_0_331), .ZN(
      n_0_0_318));
   NOR2_X1 i_0_0_388 (.A1(n_0_0_376), .A2(n_0_0_320), .ZN(n_0_0_319));
   OAI211_X1 i_0_0_389 (.A(n_0_0_321), .B(n_0_0_322), .C1(n_0_0_560), .C2(
      n_0_0_379), .ZN(n_0_0_320));
   NAND2_X1 i_0_0_390 (.A1(A[18]), .A2(n_0_0_340), .ZN(n_0_0_321));
   AOI22_X1 i_0_0_391 (.A1(A[22]), .A2(n_0_0_323), .B1(A[14]), .B2(n_0_0_359), 
      .ZN(n_0_0_322));
   NOR2_X1 i_0_0_392 (.A1(n_0_0_380), .A2(n_0_0_348), .ZN(n_0_0_323));
   INV_X1 i_0_0_393 (.A(n_0_0_324), .ZN(n_0_66));
   AOI222_X1 i_0_0_394 (.A1(n_0_0_371), .A2(n_0_0_325), .B1(A[11]), .B2(n_0_78), 
      .C1(n_0_0_363), .C2(n_0_0_330), .ZN(n_0_0_324));
   OAI21_X1 i_0_0_395 (.A(n_0_0_326), .B1(n_0_0_376), .B2(n_0_0_327), .ZN(
      n_0_0_325));
   NAND2_X1 i_0_0_396 (.A1(n_0_0_376), .A2(n_0_0_335), .ZN(n_0_0_326));
   AOI22_X1 i_0_0_397 (.A1(n_0_0_381), .A2(n_0_0_345), .B1(n_0_0_380), .B2(
      n_0_0_328), .ZN(n_0_0_327));
   OAI22_X1 i_0_0_398 (.A1(n_0_0_561), .A2(n_0_0_383), .B1(n_0_0_567), .B2(
      n_0_0_348), .ZN(n_0_0_328));
   INV_X1 i_0_0_399 (.A(n_0_0_329), .ZN(n_0_67));
   AOI222_X1 i_0_0_400 (.A1(n_0_0_371), .A2(n_0_0_330), .B1(A[12]), .B2(n_0_78), 
      .C1(n_0_0_363), .C2(n_0_0_333), .ZN(n_0_0_329));
   OAI22_X1 i_0_0_401 (.A1(n_0_0_376), .A2(n_0_0_331), .B1(n_0_0_375), .B2(
      n_0_0_339), .ZN(n_0_0_330));
   AOI222_X1 i_0_0_402 (.A1(A[16]), .A2(n_0_0_359), .B1(A[12]), .B2(n_0_0_378), 
      .C1(A[20]), .C2(n_0_0_340), .ZN(n_0_0_331));
   INV_X1 i_0_0_403 (.A(n_0_0_332), .ZN(n_0_68));
   AOI222_X1 i_0_0_404 (.A1(n_0_0_371), .A2(n_0_0_333), .B1(A[13]), .B2(n_0_78), 
      .C1(n_0_0_363), .C2(n_0_0_338), .ZN(n_0_0_332));
   OAI21_X1 i_0_0_405 (.A(n_0_0_334), .B1(n_0_0_375), .B2(n_0_0_344), .ZN(
      n_0_0_333));
   NAND2_X1 i_0_0_406 (.A1(n_0_0_375), .A2(n_0_0_335), .ZN(n_0_0_334));
   OAI21_X1 i_0_0_407 (.A(n_0_0_336), .B1(n_0_0_563), .B2(n_0_0_379), .ZN(
      n_0_0_335));
   AOI22_X1 i_0_0_408 (.A1(A[17]), .A2(n_0_0_359), .B1(A[21]), .B2(n_0_0_340), 
      .ZN(n_0_0_336));
   INV_X1 i_0_0_409 (.A(n_0_0_337), .ZN(n_0_69));
   AOI222_X1 i_0_0_410 (.A1(n_0_0_363), .A2(n_0_0_342), .B1(A[14]), .B2(n_0_78), 
      .C1(n_0_0_371), .C2(n_0_0_338), .ZN(n_0_0_337));
   AOI22_X1 i_0_0_411 (.A1(n_0_0_376), .A2(n_0_0_351), .B1(n_0_0_375), .B2(
      n_0_0_339), .ZN(n_0_0_338));
   AOI222_X1 i_0_0_412 (.A1(A[18]), .A2(n_0_0_359), .B1(A[14]), .B2(n_0_0_378), 
      .C1(A[22]), .C2(n_0_0_340), .ZN(n_0_0_339));
   NOR2_X1 i_0_0_413 (.A1(n_0_0_381), .A2(n_0_0_348), .ZN(n_0_0_340));
   INV_X1 i_0_0_414 (.A(n_0_0_341), .ZN(n_0_70));
   AOI222_X1 i_0_0_415 (.A1(n_0_0_371), .A2(n_0_0_342), .B1(A[15]), .B2(n_0_78), 
      .C1(n_0_0_363), .C2(n_0_0_350), .ZN(n_0_0_341));
   OAI21_X1 i_0_0_416 (.A(n_0_0_343), .B1(n_0_0_376), .B2(n_0_0_344), .ZN(
      n_0_0_342));
   NAND3_X1 i_0_0_417 (.A1(n_0_0_376), .A2(n_0_0_354), .A3(n_0_0_382), .ZN(
      n_0_0_343));
   AOI22_X1 i_0_0_418 (.A1(A[19]), .A2(n_0_0_359), .B1(n_0_0_380), .B2(n_0_0_345), 
      .ZN(n_0_0_344));
   NAND2_X1 i_0_0_419 (.A1(n_0_0_348), .A2(n_0_0_346), .ZN(n_0_0_345));
   NAND2_X1 i_0_0_420 (.A1(A[15]), .A2(n_0_0_386), .ZN(n_0_0_346));
   INV_X1 i_0_0_421 (.A(n_0_0_348), .ZN(n_0_0_347));
   NAND2_X1 i_0_0_422 (.A1(n_0_0_386), .A2(n_0_0_384), .ZN(n_0_0_348));
   INV_X1 i_0_0_423 (.A(n_0_0_349), .ZN(n_0_71));
   AOI222_X1 i_0_0_424 (.A1(n_0_0_363), .A2(n_0_0_353), .B1(A[16]), .B2(n_0_78), 
      .C1(n_0_0_371), .C2(n_0_0_350), .ZN(n_0_0_349));
   AOI22_X1 i_0_0_425 (.A1(n_0_0_376), .A2(n_0_0_358), .B1(n_0_0_375), .B2(
      n_0_0_351), .ZN(n_0_0_350));
   AOI22_X1 i_0_0_426 (.A1(A[16]), .A2(n_0_0_378), .B1(A[20]), .B2(n_0_0_359), 
      .ZN(n_0_0_351));
   INV_X1 i_0_0_427 (.A(n_0_0_352), .ZN(n_0_72));
   AOI222_X1 i_0_0_428 (.A1(A[17]), .A2(n_0_78), .B1(n_0_0_371), .B2(n_0_0_353), 
      .C1(n_0_0_363), .C2(n_0_0_357), .ZN(n_0_0_352));
   AOI221_X1 i_0_0_429 (.A(n_0_0_383), .B1(n_0_0_375), .B2(n_0_0_355), .C1(
      n_0_0_376), .C2(n_0_0_365), .ZN(n_0_0_353));
   INV_X1 i_0_0_430 (.A(n_0_0_355), .ZN(n_0_0_354));
   AOI22_X1 i_0_0_431 (.A1(A[17]), .A2(n_0_0_380), .B1(A[21]), .B2(n_0_0_381), 
      .ZN(n_0_0_355));
   INV_X1 i_0_0_432 (.A(n_0_0_356), .ZN(n_0_73));
   AOI222_X1 i_0_0_433 (.A1(n_0_0_364), .A2(n_0_0_363), .B1(A[18]), .B2(n_0_78), 
      .C1(n_0_0_371), .C2(n_0_0_357), .ZN(n_0_0_356));
   OAI22_X1 i_0_0_434 (.A1(n_0_0_568), .A2(n_0_0_366), .B1(n_0_0_376), .B2(
      n_0_0_358), .ZN(n_0_0_357));
   AOI22_X1 i_0_0_435 (.A1(A[18]), .A2(n_0_0_378), .B1(A[22]), .B2(n_0_0_359), 
      .ZN(n_0_0_358));
   NOR2_X1 i_0_0_436 (.A1(n_0_0_383), .A2(n_0_0_380), .ZN(n_0_0_359));
   INV_X1 i_0_0_437 (.A(n_0_0_360), .ZN(n_0_74));
   AOI221_X1 i_0_0_438 (.A(n_0_0_361), .B1(A[19]), .B2(n_0_78), .C1(n_0_0_371), 
      .C2(n_0_0_364), .ZN(n_0_0_360));
   AND3_X1 i_0_0_439 (.A1(n_0_0_378), .A2(n_0_0_362), .A3(n_0_0_363), .ZN(
      n_0_0_361));
   OAI21_X1 i_0_0_440 (.A(n_0_0_369), .B1(n_0_0_568), .B2(n_0_0_376), .ZN(
      n_0_0_362));
   AND2_X1 i_0_0_441 (.A1(n_0_0_501), .A2(n_0_0_387), .ZN(n_0_0_363));
   OAI33_X1 i_0_0_442 (.A1(n_0_0_379), .A2(n_0_0_375), .A3(n_0_0_569), .B1(
      n_0_0_383), .B2(n_0_0_376), .B3(n_0_0_365), .ZN(n_0_0_364));
   NOR2_X1 i_0_0_443 (.A1(A[19]), .A2(n_0_0_381), .ZN(n_0_0_365));
   NAND2_X1 i_0_0_444 (.A1(n_0_0_378), .A2(n_0_0_376), .ZN(n_0_0_366));
   INV_X1 i_0_0_445 (.A(n_0_0_367), .ZN(n_0_75));
   AOI22_X1 i_0_0_446 (.A1(A[20]), .A2(n_0_78), .B1(n_0_0_377), .B2(n_0_0_368), 
      .ZN(n_0_0_367));
   AOI22_X1 i_0_0_447 (.A1(n_0_0_569), .A2(n_0_0_375), .B1(n_0_0_500), .B2(
      n_0_0_369), .ZN(n_0_0_368));
   NAND2_X1 i_0_0_448 (.A1(A[22]), .A2(n_0_0_376), .ZN(n_0_0_369));
   INV_X1 i_0_0_449 (.A(n_0_0_370), .ZN(n_0_76));
   AOI222_X1 i_0_0_450 (.A1(n_0_0_378), .A2(n_0_0_371), .B1(A[21]), .B2(n_0_78), 
      .C1(A[22]), .C2(n_0_0_374), .ZN(n_0_0_370));
   INV_X1 i_0_0_451 (.A(n_0_0_372), .ZN(n_0_0_371));
   NAND2_X1 i_0_0_452 (.A1(n_0_0_500), .A2(n_0_0_387), .ZN(n_0_0_372));
   INV_X1 i_0_0_453 (.A(n_0_0_373), .ZN(n_0_77));
   AOI21_X1 i_0_0_454 (.A(n_0_0_374), .B1(A[22]), .B2(n_0_78), .ZN(n_0_0_373));
   AND2_X1 i_0_0_455 (.A1(n_0_0_377), .A2(n_0_0_375), .ZN(n_0_0_374));
   INV_X1 i_0_0_456 (.A(n_0_0_376), .ZN(n_0_0_375));
   XNOR2_X1 i_0_0_457 (.A(n_0_0_521), .B(n_0_0_492), .ZN(n_0_0_376));
   AND2_X1 i_0_0_458 (.A1(n_0_0_387), .A2(n_0_0_378), .ZN(n_0_0_377));
   INV_X1 i_0_0_459 (.A(n_0_0_379), .ZN(n_0_0_378));
   NAND2_X1 i_0_0_460 (.A1(n_0_0_382), .A2(n_0_0_380), .ZN(n_0_0_379));
   INV_X1 i_0_0_461 (.A(n_0_0_381), .ZN(n_0_0_380));
   XNOR2_X1 i_0_0_462 (.A(n_0_0_524), .B(n_0_0_520), .ZN(n_0_0_381));
   INV_X1 i_0_0_463 (.A(n_0_0_383), .ZN(n_0_0_382));
   NAND2_X1 i_0_0_464 (.A1(n_0_0_386), .A2(n_0_0_385), .ZN(n_0_0_383));
   INV_X1 i_0_0_465 (.A(n_0_0_385), .ZN(n_0_0_384));
   AOI22_X1 i_0_0_466 (.A1(n_0_0_528), .A2(n_0_0_518), .B1(n_0_0_527), .B2(
      n_0_0_519), .ZN(n_0_0_385));
   XNOR2_X1 i_0_0_467 (.A(n_0_0_517), .B(n_0_0_515), .ZN(n_0_0_386));
   AOI21_X1 i_0_0_468 (.A(n_0_78), .B1(n_0_0_391), .B2(n_0_0_388), .ZN(n_0_0_387));
   NAND2_X1 i_0_0_469 (.A1(n_0_0_514), .A2(n_0_0_389), .ZN(n_0_0_388));
   OAI33_X1 i_0_0_470 (.A1(B[28]), .A2(n_0_0_573), .A3(n_0_0_390), .B1(n_0_0_598), 
      .B2(A[28]), .B3(n_0_0_534), .ZN(n_0_0_389));
   AOI22_X1 i_0_0_471 (.A1(n_0_0_599), .A2(A[29]), .B1(n_0_0_541), .B2(n_0_0_536), 
      .ZN(n_0_0_390));
   OR2_X1 i_0_0_472 (.A1(n_0_0_514), .A2(n_0_0_504), .ZN(n_0_0_391));
   INV_X1 i_0_0_473 (.A(n_0_0_392), .ZN(n_0_78));
   AOI21_X1 i_0_0_474 (.A(n_0_0_532), .B1(n_0_0_531), .B2(n_0_0_506), .ZN(
      n_0_0_392));
   INV_X1 i_0_0_475 (.A(n_0_0_393), .ZN(n_0_79));
   AOI221_X1 i_0_0_476 (.A(n_0_0_394), .B1(B[0]), .B2(n_0_102), .C1(n_0_0_498), 
      .C2(n_0_0_398), .ZN(n_0_0_393));
   AOI221_X1 i_0_0_477 (.A(n_0_0_484), .B1(n_0_0_396), .B2(n_0_0_395), .C1(
      n_0_0_492), .C2(n_0_0_404), .ZN(n_0_0_394));
   AOI222_X1 i_0_0_478 (.A1(B[8]), .A2(n_0_0_461), .B1(B[16]), .B2(n_0_0_411), 
      .C1(n_0_0_487), .C2(n_0_0_415), .ZN(n_0_0_395));
   AOI21_X1 i_0_0_479 (.A(n_0_0_492), .B1(B[0]), .B2(n_0_0_481), .ZN(n_0_0_396));
   INV_X1 i_0_0_480 (.A(n_0_0_397), .ZN(n_0_80));
   AOI222_X1 i_0_0_481 (.A1(n_0_0_483), .A2(n_0_0_398), .B1(B[1]), .B2(n_0_102), 
      .C1(n_0_0_498), .C2(n_0_0_403), .ZN(n_0_0_397));
   AOI22_X1 i_0_0_482 (.A1(n_0_0_490), .A2(n_0_0_408), .B1(n_0_0_491), .B2(
      n_0_0_399), .ZN(n_0_0_398));
   AOI221_X1 i_0_0_483 (.A(n_0_0_400), .B1(B[1]), .B2(n_0_0_481), .C1(B[17]), 
      .C2(n_0_0_411), .ZN(n_0_0_399));
   OAI21_X1 i_0_0_484 (.A(n_0_0_401), .B1(n_0_0_488), .B2(n_0_0_421), .ZN(
      n_0_0_400));
   NAND2_X1 i_0_0_485 (.A1(B[9]), .A2(n_0_0_461), .ZN(n_0_0_401));
   INV_X1 i_0_0_486 (.A(n_0_0_402), .ZN(n_0_81));
   AOI222_X1 i_0_0_487 (.A1(n_0_0_498), .A2(n_0_0_407), .B1(B[2]), .B2(n_0_102), 
      .C1(n_0_0_483), .C2(n_0_0_403), .ZN(n_0_0_402));
   AOI22_X1 i_0_0_488 (.A1(n_0_0_491), .A2(n_0_0_404), .B1(n_0_0_490), .B2(
      n_0_0_414), .ZN(n_0_0_403));
   AOI221_X1 i_0_0_489 (.A(n_0_0_405), .B1(B[18]), .B2(n_0_0_411), .C1(B[10]), 
      .C2(n_0_0_461), .ZN(n_0_0_404));
   OAI22_X1 i_0_0_490 (.A1(n_0_0_488), .A2(n_0_0_426), .B1(n_0_0_577), .B2(
      n_0_0_482), .ZN(n_0_0_405));
   INV_X1 i_0_0_491 (.A(n_0_0_406), .ZN(n_0_82));
   AOI222_X1 i_0_0_492 (.A1(n_0_0_483), .A2(n_0_0_407), .B1(B[3]), .B2(n_0_102), 
      .C1(n_0_0_498), .C2(n_0_0_413), .ZN(n_0_0_406));
   AOI22_X1 i_0_0_493 (.A1(n_0_0_491), .A2(n_0_0_408), .B1(n_0_0_490), .B2(
      n_0_0_419), .ZN(n_0_0_407));
   AOI221_X1 i_0_0_494 (.A(n_0_0_409), .B1(B[3]), .B2(n_0_0_481), .C1(B[11]), 
      .C2(n_0_0_461), .ZN(n_0_0_408));
   INV_X1 i_0_0_495 (.A(n_0_0_410), .ZN(n_0_0_409));
   AOI22_X1 i_0_0_496 (.A1(n_0_0_487), .A2(n_0_0_432), .B1(B[19]), .B2(n_0_0_411), 
      .ZN(n_0_0_410));
   AND2_X1 i_0_0_497 (.A1(n_0_0_488), .A2(n_0_0_427), .ZN(n_0_0_411));
   INV_X1 i_0_0_498 (.A(n_0_0_412), .ZN(n_0_83));
   AOI222_X1 i_0_0_499 (.A1(n_0_0_498), .A2(n_0_0_418), .B1(B[4]), .B2(n_0_102), 
      .C1(n_0_0_483), .C2(n_0_0_413), .ZN(n_0_0_412));
   AOI22_X1 i_0_0_500 (.A1(n_0_0_491), .A2(n_0_0_414), .B1(n_0_0_490), .B2(
      n_0_0_424), .ZN(n_0_0_413));
   AOI222_X1 i_0_0_501 (.A1(B[8]), .A2(n_0_0_460), .B1(B[16]), .B2(n_0_0_431), 
      .C1(n_0_0_488), .C2(n_0_0_415), .ZN(n_0_0_414));
   INV_X1 i_0_0_502 (.A(n_0_0_416), .ZN(n_0_0_415));
   AOI222_X1 i_0_0_503 (.A1(B[20]), .A2(n_0_0_427), .B1(B[12]), .B2(n_0_0_462), 
      .C1(B[4]), .C2(n_0_0_493), .ZN(n_0_0_416));
   OAI21_X1 i_0_0_504 (.A(n_0_0_417), .B1(n_0_0_580), .B2(n_0_0_513), .ZN(n_0_84));
   AOI22_X1 i_0_0_505 (.A1(n_0_0_483), .A2(n_0_0_418), .B1(n_0_0_498), .B2(
      n_0_0_423), .ZN(n_0_0_417));
   AOI22_X1 i_0_0_506 (.A1(n_0_0_491), .A2(n_0_0_419), .B1(n_0_0_490), .B2(
      n_0_0_430), .ZN(n_0_0_418));
   AOI222_X1 i_0_0_507 (.A1(B[17]), .A2(n_0_0_431), .B1(B[9]), .B2(n_0_0_460), 
      .C1(n_0_0_488), .C2(n_0_0_420), .ZN(n_0_0_419));
   INV_X1 i_0_0_508 (.A(n_0_0_421), .ZN(n_0_0_420));
   AOI222_X1 i_0_0_509 (.A1(B[21]), .A2(n_0_0_427), .B1(B[5]), .B2(n_0_0_493), 
      .C1(B[13]), .C2(n_0_0_462), .ZN(n_0_0_421));
   INV_X1 i_0_0_510 (.A(n_0_0_422), .ZN(n_0_85));
   AOI222_X1 i_0_0_511 (.A1(B[6]), .A2(n_0_102), .B1(n_0_0_498), .B2(n_0_0_429), 
      .C1(n_0_0_483), .C2(n_0_0_423), .ZN(n_0_0_422));
   AOI22_X1 i_0_0_512 (.A1(n_0_0_491), .A2(n_0_0_424), .B1(n_0_0_490), .B2(
      n_0_0_436), .ZN(n_0_0_423));
   AOI222_X1 i_0_0_513 (.A1(B[18]), .A2(n_0_0_431), .B1(B[10]), .B2(n_0_0_460), 
      .C1(n_0_0_488), .C2(n_0_0_425), .ZN(n_0_0_424));
   INV_X1 i_0_0_514 (.A(n_0_0_426), .ZN(n_0_0_425));
   AOI222_X1 i_0_0_515 (.A1(B[22]), .A2(n_0_0_427), .B1(B[6]), .B2(n_0_0_493), 
      .C1(B[14]), .C2(n_0_0_462), .ZN(n_0_0_426));
   NOR2_X1 i_0_0_516 (.A1(n_0_0_496), .A2(n_0_0_494), .ZN(n_0_0_427));
   INV_X1 i_0_0_517 (.A(n_0_0_428), .ZN(n_0_86));
   AOI222_X1 i_0_0_518 (.A1(B[7]), .A2(n_0_102), .B1(n_0_0_498), .B2(n_0_0_435), 
      .C1(n_0_0_483), .C2(n_0_0_429), .ZN(n_0_0_428));
   AOI22_X1 i_0_0_519 (.A1(n_0_0_491), .A2(n_0_0_430), .B1(n_0_0_490), .B2(
      n_0_0_439), .ZN(n_0_0_429));
   AOI222_X1 i_0_0_520 (.A1(B[19]), .A2(n_0_0_431), .B1(B[11]), .B2(n_0_0_460), 
      .C1(n_0_0_488), .C2(n_0_0_432), .ZN(n_0_0_430));
   NOR3_X1 i_0_0_521 (.A1(n_0_0_497), .A2(n_0_0_495), .A3(n_0_0_488), .ZN(
      n_0_0_431));
   AOI21_X1 i_0_0_522 (.A(n_0_0_433), .B1(n_0_0_582), .B2(n_0_0_493), .ZN(
      n_0_0_432));
   AOI21_X1 i_0_0_523 (.A(n_0_0_497), .B1(B[15]), .B2(n_0_0_494), .ZN(n_0_0_433));
   INV_X1 i_0_0_524 (.A(n_0_0_434), .ZN(n_0_87));
   AOI222_X1 i_0_0_525 (.A1(n_0_0_498), .A2(n_0_0_438), .B1(B[8]), .B2(n_0_102), 
      .C1(n_0_0_483), .C2(n_0_0_435), .ZN(n_0_0_434));
   AOI22_X1 i_0_0_526 (.A1(n_0_0_491), .A2(n_0_0_436), .B1(n_0_0_490), .B2(
      n_0_0_442), .ZN(n_0_0_435));
   AOI222_X1 i_0_0_527 (.A1(B[8]), .A2(n_0_0_481), .B1(n_0_0_465), .B2(n_0_0_462), 
      .C1(B[12]), .C2(n_0_0_460), .ZN(n_0_0_436));
   INV_X1 i_0_0_528 (.A(n_0_0_437), .ZN(n_0_88));
   AOI222_X1 i_0_0_529 (.A1(n_0_0_483), .A2(n_0_0_438), .B1(B[9]), .B2(n_0_102), 
      .C1(n_0_0_498), .C2(n_0_0_441), .ZN(n_0_0_437));
   AOI22_X1 i_0_0_530 (.A1(n_0_0_491), .A2(n_0_0_439), .B1(n_0_0_490), .B2(
      n_0_0_445), .ZN(n_0_0_438));
   AOI222_X1 i_0_0_531 (.A1(B[9]), .A2(n_0_0_481), .B1(n_0_0_467), .B2(n_0_0_462), 
      .C1(B[13]), .C2(n_0_0_460), .ZN(n_0_0_439));
   OAI21_X1 i_0_0_532 (.A(n_0_0_440), .B1(n_0_0_585), .B2(n_0_0_513), .ZN(n_0_89));
   AOI22_X1 i_0_0_533 (.A1(n_0_0_483), .A2(n_0_0_441), .B1(n_0_0_498), .B2(
      n_0_0_444), .ZN(n_0_0_440));
   AOI22_X1 i_0_0_534 (.A1(n_0_0_491), .A2(n_0_0_442), .B1(n_0_0_490), .B2(
      n_0_0_448), .ZN(n_0_0_441));
   AOI222_X1 i_0_0_535 (.A1(B[10]), .A2(n_0_0_481), .B1(n_0_0_469), .B2(
      n_0_0_462), .C1(B[14]), .C2(n_0_0_460), .ZN(n_0_0_442));
   INV_X1 i_0_0_536 (.A(n_0_0_443), .ZN(n_0_90));
   AOI222_X1 i_0_0_537 (.A1(n_0_0_483), .A2(n_0_0_444), .B1(B[11]), .B2(n_0_102), 
      .C1(n_0_0_498), .C2(n_0_0_447), .ZN(n_0_0_443));
   AOI22_X1 i_0_0_538 (.A1(n_0_0_491), .A2(n_0_0_445), .B1(n_0_0_490), .B2(
      n_0_0_451), .ZN(n_0_0_444));
   AOI222_X1 i_0_0_539 (.A1(B[11]), .A2(n_0_0_481), .B1(n_0_0_473), .B2(
      n_0_0_462), .C1(B[15]), .C2(n_0_0_460), .ZN(n_0_0_445));
   OAI21_X1 i_0_0_540 (.A(n_0_0_446), .B1(n_0_0_587), .B2(n_0_0_513), .ZN(n_0_91));
   AOI22_X1 i_0_0_541 (.A1(n_0_0_498), .A2(n_0_0_450), .B1(n_0_0_483), .B2(
      n_0_0_447), .ZN(n_0_0_446));
   AOI22_X1 i_0_0_542 (.A1(n_0_0_491), .A2(n_0_0_448), .B1(n_0_0_490), .B2(
      n_0_0_454), .ZN(n_0_0_447));
   AOI222_X1 i_0_0_543 (.A1(B[16]), .A2(n_0_0_460), .B1(B[12]), .B2(n_0_0_481), 
      .C1(B[20]), .C2(n_0_0_461), .ZN(n_0_0_448));
   INV_X1 i_0_0_544 (.A(n_0_0_449), .ZN(n_0_92));
   AOI222_X1 i_0_0_545 (.A1(n_0_0_498), .A2(n_0_0_453), .B1(B[13]), .B2(n_0_102), 
      .C1(n_0_0_483), .C2(n_0_0_450), .ZN(n_0_0_449));
   AOI22_X1 i_0_0_546 (.A1(n_0_0_491), .A2(n_0_0_451), .B1(n_0_0_490), .B2(
      n_0_0_459), .ZN(n_0_0_450));
   AOI222_X1 i_0_0_547 (.A1(B[17]), .A2(n_0_0_460), .B1(B[13]), .B2(n_0_0_481), 
      .C1(B[21]), .C2(n_0_0_461), .ZN(n_0_0_451));
   INV_X1 i_0_0_548 (.A(n_0_0_452), .ZN(n_0_93));
   AOI222_X1 i_0_0_549 (.A1(B[14]), .A2(n_0_102), .B1(n_0_0_483), .B2(n_0_0_453), 
      .C1(n_0_0_498), .C2(n_0_0_458), .ZN(n_0_0_452));
   OAI21_X1 i_0_0_550 (.A(n_0_0_455), .B1(n_0_0_490), .B2(n_0_0_454), .ZN(
      n_0_0_453));
   AOI222_X1 i_0_0_551 (.A1(B[22]), .A2(n_0_0_461), .B1(B[18]), .B2(n_0_0_460), 
      .C1(B[14]), .C2(n_0_0_481), .ZN(n_0_0_454));
   NAND2_X1 i_0_0_552 (.A1(n_0_0_480), .A2(n_0_0_465), .ZN(n_0_0_455));
   INV_X1 i_0_0_553 (.A(n_0_0_456), .ZN(n_0_94));
   AOI21_X1 i_0_0_554 (.A(n_0_0_457), .B1(n_0_0_483), .B2(n_0_0_458), .ZN(
      n_0_0_456));
   OAI22_X1 i_0_0_555 (.A1(n_0_0_588), .A2(n_0_0_513), .B1(n_0_0_499), .B2(
      n_0_0_464), .ZN(n_0_0_457));
   OAI21_X1 i_0_0_556 (.A(n_0_0_463), .B1(n_0_0_490), .B2(n_0_0_459), .ZN(
      n_0_0_458));
   AOI221_X1 i_0_0_557 (.A(n_0_0_461), .B1(B[19]), .B2(n_0_0_460), .C1(B[15]), 
      .C2(n_0_0_481), .ZN(n_0_0_459));
   NOR3_X1 i_0_0_558 (.A1(n_0_0_496), .A2(n_0_0_495), .A3(n_0_0_488), .ZN(
      n_0_0_460));
   NOR3_X1 i_0_0_559 (.A1(n_0_0_497), .A2(n_0_0_495), .A3(n_0_0_487), .ZN(
      n_0_0_461));
   NOR2_X1 i_0_0_560 (.A1(n_0_0_497), .A2(n_0_0_495), .ZN(n_0_0_462));
   NAND2_X1 i_0_0_561 (.A1(n_0_0_480), .A2(n_0_0_467), .ZN(n_0_0_463));
   OAI222_X1 i_0_0_562 (.A1(n_0_0_499), .A2(n_0_0_466), .B1(n_0_0_589), .B2(
      n_0_0_513), .C1(n_0_0_484), .C2(n_0_0_464), .ZN(n_0_95));
   AOI22_X1 i_0_0_563 (.A1(n_0_0_480), .A2(n_0_0_469), .B1(n_0_0_489), .B2(
      n_0_0_465), .ZN(n_0_0_464));
   OAI22_X1 i_0_0_564 (.A1(n_0_0_589), .A2(n_0_0_487), .B1(n_0_0_593), .B2(
      n_0_0_488), .ZN(n_0_0_465));
   OAI222_X1 i_0_0_565 (.A1(n_0_0_590), .A2(n_0_0_513), .B1(n_0_0_484), .B2(
      n_0_0_466), .C1(n_0_0_499), .C2(n_0_0_468), .ZN(n_0_96));
   AOI22_X1 i_0_0_566 (.A1(n_0_0_480), .A2(n_0_0_473), .B1(n_0_0_489), .B2(
      n_0_0_467), .ZN(n_0_0_466));
   OAI22_X1 i_0_0_567 (.A1(n_0_0_590), .A2(n_0_0_487), .B1(n_0_0_594), .B2(
      n_0_0_488), .ZN(n_0_0_467));
   OAI222_X1 i_0_0_568 (.A1(n_0_0_499), .A2(n_0_0_472), .B1(n_0_0_591), .B2(
      n_0_0_513), .C1(n_0_0_484), .C2(n_0_0_468), .ZN(n_0_97));
   AOI22_X1 i_0_0_569 (.A1(n_0_0_489), .A2(n_0_0_469), .B1(B[20]), .B2(n_0_0_479), 
      .ZN(n_0_0_468));
   AOI22_X1 i_0_0_570 (.A1(n_0_0_591), .A2(n_0_0_488), .B1(n_0_0_595), .B2(
      n_0_0_487), .ZN(n_0_0_469));
   OAI21_X1 i_0_0_571 (.A(n_0_0_470), .B1(n_0_0_484), .B2(n_0_0_472), .ZN(n_0_98));
   AOI21_X1 i_0_0_572 (.A(n_0_0_471), .B1(B[19]), .B2(n_0_102), .ZN(n_0_0_470));
   NOR3_X1 i_0_0_573 (.A1(n_0_0_482), .A2(n_0_0_477), .A3(n_0_0_499), .ZN(
      n_0_0_471));
   AOI22_X1 i_0_0_574 (.A1(n_0_0_489), .A2(n_0_0_473), .B1(B[21]), .B2(n_0_0_479), 
      .ZN(n_0_0_472));
   NAND2_X1 i_0_0_575 (.A1(n_0_0_592), .A2(n_0_0_488), .ZN(n_0_0_473));
   INV_X1 i_0_0_576 (.A(n_0_0_474), .ZN(n_0_99));
   AOI22_X1 i_0_0_577 (.A1(B[20]), .A2(n_0_102), .B1(n_0_0_502), .B2(n_0_0_475), 
      .ZN(n_0_0_474));
   AOI211_X1 i_0_0_578 (.A(n_0_0_482), .B(n_0_0_476), .C1(n_0_0_500), .C2(
      n_0_0_477), .ZN(n_0_0_475));
   NOR3_X1 i_0_0_579 (.A1(B[21]), .A2(n_0_0_500), .A3(n_0_0_490), .ZN(n_0_0_476));
   AOI22_X1 i_0_0_580 (.A1(B[22]), .A2(n_0_0_490), .B1(B[20]), .B2(n_0_0_491), 
      .ZN(n_0_0_477));
   OAI21_X1 i_0_0_581 (.A(n_0_0_478), .B1(n_0_0_594), .B2(n_0_0_513), .ZN(
      n_0_100));
   AOI22_X1 i_0_0_582 (.A1(B[22]), .A2(n_0_0_486), .B1(n_0_0_483), .B2(n_0_0_479), 
      .ZN(n_0_0_478));
   NOR2_X1 i_0_0_583 (.A1(n_0_0_491), .A2(n_0_0_482), .ZN(n_0_0_479));
   NOR3_X1 i_0_0_584 (.A1(n_0_0_496), .A2(n_0_0_495), .A3(n_0_0_491), .ZN(
      n_0_0_480));
   INV_X1 i_0_0_585 (.A(n_0_0_482), .ZN(n_0_0_481));
   NAND2_X1 i_0_0_586 (.A1(n_0_0_493), .A2(n_0_0_488), .ZN(n_0_0_482));
   INV_X1 i_0_0_587 (.A(n_0_0_484), .ZN(n_0_0_483));
   NAND2_X1 i_0_0_588 (.A1(n_0_0_502), .A2(n_0_0_500), .ZN(n_0_0_484));
   INV_X1 i_0_0_589 (.A(n_0_0_485), .ZN(n_0_101));
   AOI21_X1 i_0_0_590 (.A(n_0_0_486), .B1(B[22]), .B2(n_0_102), .ZN(n_0_0_485));
   AND3_X1 i_0_0_591 (.A1(n_0_0_489), .A2(n_0_0_488), .A3(n_0_0_498), .ZN(
      n_0_0_486));
   INV_X1 i_0_0_592 (.A(n_0_0_488), .ZN(n_0_0_487));
   XNOR2_X1 i_0_0_593 (.A(n_0_0_524), .B(n_0_0_510), .ZN(n_0_0_488));
   NOR3_X1 i_0_0_594 (.A1(n_0_0_496), .A2(n_0_0_495), .A3(n_0_0_490), .ZN(
      n_0_0_489));
   INV_X1 i_0_0_595 (.A(n_0_0_491), .ZN(n_0_0_490));
   XNOR2_X1 i_0_0_596 (.A(n_0_0_511), .B(n_0_0_492), .ZN(n_0_0_491));
   OAI21_X1 i_0_0_597 (.A(n_0_0_523), .B1(n_0_0_596), .B2(A[24]), .ZN(n_0_0_492));
   NOR2_X1 i_0_0_598 (.A1(n_0_0_496), .A2(n_0_0_495), .ZN(n_0_0_493));
   INV_X1 i_0_0_599 (.A(n_0_0_495), .ZN(n_0_0_494));
   XNOR2_X1 i_0_0_600 (.A(n_0_0_515), .B(n_0_0_507), .ZN(n_0_0_495));
   INV_X1 i_0_0_601 (.A(n_0_0_497), .ZN(n_0_0_496));
   XNOR2_X1 i_0_0_602 (.A(n_0_0_527), .B(n_0_0_509), .ZN(n_0_0_497));
   INV_X1 i_0_0_603 (.A(n_0_0_499), .ZN(n_0_0_498));
   NAND2_X1 i_0_0_604 (.A1(n_0_0_502), .A2(n_0_0_501), .ZN(n_0_0_499));
   INV_X1 i_0_0_605 (.A(n_0_0_501), .ZN(n_0_0_500));
   NAND2_X1 i_0_0_606 (.A1(n_0_0_521), .A2(n_0_0_512), .ZN(n_0_0_501));
   AOI221_X1 i_0_0_607 (.A(n_0_102), .B1(n_0_0_533), .B2(n_0_0_503), .C1(
      n_0_0_506), .C2(n_0_0_504), .ZN(n_0_0_502));
   AOI21_X1 i_0_0_608 (.A(n_0_0_506), .B1(n_0_0_539), .B2(n_0_0_505), .ZN(
      n_0_0_503));
   NAND3_X1 i_0_0_609 (.A1(n_0_0_537), .A2(n_0_0_533), .A3(n_0_0_531), .ZN(
      n_0_0_504));
   AOI211_X1 i_0_0_610 (.A(n_0_0_598), .B(A[28]), .C1(n_0_0_542), .C2(n_0_0_535), 
      .ZN(n_0_0_505));
   OAI21_X1 i_0_0_611 (.A(n_0_0_516), .B1(n_0_0_530), .B2(n_0_0_507), .ZN(
      n_0_0_506));
   NOR2_X1 i_0_0_612 (.A1(n_0_0_529), .A2(n_0_0_508), .ZN(n_0_0_507));
   AOI21_X1 i_0_0_613 (.A(n_0_0_509), .B1(B[26]), .B2(n_0_0_572), .ZN(n_0_0_508));
   AOI21_X1 i_0_0_614 (.A(n_0_0_526), .B1(n_0_0_525), .B2(n_0_0_510), .ZN(
      n_0_0_509));
   AOI21_X1 i_0_0_615 (.A(n_0_0_522), .B1(n_0_0_523), .B2(n_0_0_511), .ZN(
      n_0_0_510));
   INV_X1 i_0_0_616 (.A(n_0_0_512), .ZN(n_0_0_511));
   NAND2_X1 i_0_0_617 (.A1(B[23]), .A2(n_0_0_570), .ZN(n_0_0_512));
   INV_X1 i_0_0_618 (.A(n_0_102), .ZN(n_0_0_513));
   AOI21_X1 i_0_0_619 (.A(n_0_0_532), .B1(n_0_0_531), .B2(n_0_0_514), .ZN(
      n_0_102));
   AOI21_X1 i_0_0_620 (.A(n_0_0_530), .B1(n_0_0_517), .B2(n_0_0_515), .ZN(
      n_0_0_514));
   AOI21_X1 i_0_0_621 (.A(n_0_0_530), .B1(n_0_0_597), .B2(A[27]), .ZN(n_0_0_515));
   NAND2_X1 i_0_0_622 (.A1(n_0_0_597), .A2(A[27]), .ZN(n_0_0_516));
   AOI21_X1 i_0_0_623 (.A(n_0_0_529), .B1(n_0_0_528), .B2(n_0_0_518), .ZN(
      n_0_0_517));
   INV_X1 i_0_0_624 (.A(n_0_0_519), .ZN(n_0_0_518));
   AOI21_X1 i_0_0_625 (.A(n_0_0_526), .B1(n_0_0_524), .B2(n_0_0_520), .ZN(
      n_0_0_519));
   AOI21_X1 i_0_0_626 (.A(n_0_0_522), .B1(n_0_0_523), .B2(n_0_0_521), .ZN(
      n_0_0_520));
   OR2_X1 i_0_0_627 (.A1(B[23]), .A2(n_0_0_570), .ZN(n_0_0_521));
   NOR2_X1 i_0_0_628 (.A1(n_0_0_596), .A2(A[24]), .ZN(n_0_0_522));
   NAND2_X1 i_0_0_629 (.A1(n_0_0_596), .A2(A[24]), .ZN(n_0_0_523));
   AOI21_X1 i_0_0_630 (.A(n_0_0_526), .B1(B[25]), .B2(n_0_0_571), .ZN(n_0_0_524));
   NAND2_X1 i_0_0_631 (.A1(B[25]), .A2(n_0_0_571), .ZN(n_0_0_525));
   NOR2_X1 i_0_0_632 (.A1(B[25]), .A2(n_0_0_571), .ZN(n_0_0_526));
   INV_X1 i_0_0_633 (.A(n_0_0_528), .ZN(n_0_0_527));
   AOI21_X1 i_0_0_634 (.A(n_0_0_529), .B1(B[26]), .B2(n_0_0_572), .ZN(n_0_0_528));
   NOR2_X1 i_0_0_635 (.A1(B[26]), .A2(n_0_0_572), .ZN(n_0_0_529));
   NOR2_X1 i_0_0_636 (.A1(n_0_0_597), .A2(A[27]), .ZN(n_0_0_530));
   AOI221_X1 i_0_0_637 (.A(n_0_0_536), .B1(B[30]), .B2(n_0_0_574), .C1(B[28]), 
      .C2(n_0_0_573), .ZN(n_0_0_531));
   NAND2_X1 i_0_0_638 (.A1(n_0_0_537), .A2(n_0_0_533), .ZN(n_0_0_532));
   OR3_X1 i_0_0_639 (.A1(B[28]), .A2(n_0_0_573), .A3(n_0_0_534), .ZN(n_0_0_533));
   NAND2_X1 i_0_0_640 (.A1(n_0_0_540), .A2(n_0_0_535), .ZN(n_0_0_534));
   INV_X1 i_0_0_641 (.A(n_0_0_536), .ZN(n_0_0_535));
   NOR2_X1 i_0_0_642 (.A1(n_0_0_599), .A2(A[29]), .ZN(n_0_0_536));
   INV_X1 i_0_0_643 (.A(n_0_0_538), .ZN(n_0_0_537));
   AOI21_X1 i_0_0_644 (.A(n_0_0_540), .B1(B[30]), .B2(n_0_0_574), .ZN(n_0_0_538));
   INV_X1 i_0_0_645 (.A(n_0_0_540), .ZN(n_0_0_539));
   AOI21_X1 i_0_0_646 (.A(n_0_0_542), .B1(n_0_0_599), .B2(A[29]), .ZN(n_0_0_540));
   INV_X1 i_0_0_647 (.A(n_0_0_542), .ZN(n_0_0_541));
   AOI21_X1 i_0_0_648 (.A(n_0_0_543), .B1(B[30]), .B2(A[30]), .ZN(n_0_0_542));
   INV_X1 i_0_0_649 (.A(n_0_0_543), .ZN(exp_Sum[7]));
   NOR2_X1 i_0_0_650 (.A1(B[30]), .A2(A[30]), .ZN(n_0_0_543));
   INV_X1 i_0_0_651 (.A(n_0_0_6), .ZN(n_0_0_544));
   INV_X1 i_0_0_652 (.A(n_0_53), .ZN(n_0_0_545));
   INV_X1 i_0_0_653 (.A(n_0_29), .ZN(n_0_0_546));
   INV_X1 i_0_0_654 (.A(n_0_1), .ZN(n_0_0_547));
   INV_X1 i_0_0_655 (.A(n_0_2), .ZN(n_0_0_548));
   INV_X1 i_0_0_656 (.A(n_0_3), .ZN(n_0_0_549));
   INV_X1 i_0_0_657 (.A(n_0_4), .ZN(n_0_0_550));
   INV_X1 i_0_0_658 (.A(A[1]), .ZN(n_0_0_551));
   INV_X1 i_0_0_659 (.A(A[2]), .ZN(n_0_0_552));
   INV_X1 i_0_0_660 (.A(A[3]), .ZN(n_0_0_553));
   INV_X1 i_0_0_661 (.A(A[4]), .ZN(n_0_0_554));
   INV_X1 i_0_0_662 (.A(A[5]), .ZN(n_0_0_555));
   INV_X1 i_0_0_663 (.A(A[6]), .ZN(n_0_0_556));
   INV_X1 i_0_0_664 (.A(A[7]), .ZN(n_0_0_557));
   INV_X1 i_0_0_665 (.A(A[8]), .ZN(n_0_0_558));
   INV_X1 i_0_0_666 (.A(A[9]), .ZN(n_0_0_559));
   INV_X1 i_0_0_667 (.A(A[10]), .ZN(n_0_0_560));
   INV_X1 i_0_0_668 (.A(A[11]), .ZN(n_0_0_561));
   INV_X1 i_0_0_669 (.A(A[12]), .ZN(n_0_0_562));
   INV_X1 i_0_0_670 (.A(A[13]), .ZN(n_0_0_563));
   INV_X1 i_0_0_671 (.A(A[14]), .ZN(n_0_0_564));
   INV_X1 i_0_0_672 (.A(A[17]), .ZN(n_0_0_565));
   INV_X1 i_0_0_673 (.A(A[18]), .ZN(n_0_0_566));
   INV_X1 i_0_0_674 (.A(A[19]), .ZN(n_0_0_567));
   INV_X1 i_0_0_675 (.A(A[20]), .ZN(n_0_0_568));
   INV_X1 i_0_0_676 (.A(A[21]), .ZN(n_0_0_569));
   INV_X1 i_0_0_677 (.A(A[23]), .ZN(n_0_0_570));
   INV_X1 i_0_0_678 (.A(A[25]), .ZN(n_0_0_571));
   INV_X1 i_0_0_679 (.A(A[26]), .ZN(n_0_0_572));
   INV_X1 i_0_0_680 (.A(A[28]), .ZN(n_0_0_573));
   INV_X1 i_0_0_681 (.A(A[30]), .ZN(n_0_0_574));
   INV_X1 i_0_0_682 (.A(B[0]), .ZN(n_0_0_575));
   INV_X1 i_0_0_683 (.A(B[1]), .ZN(n_0_0_576));
   INV_X1 i_0_0_684 (.A(B[2]), .ZN(n_0_0_577));
   INV_X1 i_0_0_685 (.A(B[3]), .ZN(n_0_0_578));
   INV_X1 i_0_0_686 (.A(B[4]), .ZN(n_0_0_579));
   INV_X1 i_0_0_687 (.A(B[5]), .ZN(n_0_0_580));
   INV_X1 i_0_0_688 (.A(B[6]), .ZN(n_0_0_581));
   INV_X1 i_0_0_689 (.A(B[7]), .ZN(n_0_0_582));
   INV_X1 i_0_0_690 (.A(B[8]), .ZN(n_0_0_583));
   INV_X1 i_0_0_691 (.A(B[9]), .ZN(n_0_0_584));
   INV_X1 i_0_0_692 (.A(B[10]), .ZN(n_0_0_585));
   INV_X1 i_0_0_693 (.A(B[11]), .ZN(n_0_0_586));
   INV_X1 i_0_0_694 (.A(B[12]), .ZN(n_0_0_587));
   INV_X1 i_0_0_695 (.A(B[15]), .ZN(n_0_0_588));
   INV_X1 i_0_0_696 (.A(B[16]), .ZN(n_0_0_589));
   INV_X1 i_0_0_697 (.A(B[17]), .ZN(n_0_0_590));
   INV_X1 i_0_0_698 (.A(B[18]), .ZN(n_0_0_591));
   INV_X1 i_0_0_699 (.A(B[19]), .ZN(n_0_0_592));
   INV_X1 i_0_0_700 (.A(B[20]), .ZN(n_0_0_593));
   INV_X1 i_0_0_701 (.A(B[21]), .ZN(n_0_0_594));
   INV_X1 i_0_0_702 (.A(B[22]), .ZN(n_0_0_595));
   INV_X1 i_0_0_703 (.A(B[24]), .ZN(n_0_0_596));
   INV_X1 i_0_0_704 (.A(B[27]), .ZN(n_0_0_597));
   INV_X1 i_0_0_705 (.A(B[28]), .ZN(n_0_0_598));
   INV_X1 i_0_0_706 (.A(B[29]), .ZN(n_0_0_599));
   INV_X1 i_0_0_707 (.A(B[31]), .ZN(n_0_0_600));
endmodule
