
// 	Wed Jan  4 06:17:00 2023
//	vlsi
//	localhost.localdomain

module datapath__0_12 (p_0, tempResult, p_1);

output [63:0] p_1;
input [63:0] p_0;
input [63:0] tempResult;
wire n_0;
wire n_366;
wire n_1;
wire n_365;
wire n_364;
wire n_2;
wire n_369;
wire n_363;
wire n_3;
wire n_370;
wire n_376;
wire n_372;
wire n_361;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_358;
wire n_349;
wire n_11;
wire n_5;
wire n_359;
wire n_353;
wire n_8;
wire n_356;
wire n_354;
wire n_360;
wire n_351;
wire n_347;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_344;
wire n_335;
wire n_19;
wire n_13;
wire n_345;
wire n_339;
wire n_16;
wire n_342;
wire n_340;
wire n_346;
wire n_337;
wire n_333;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_330;
wire n_321;
wire n_27;
wire n_21;
wire n_331;
wire n_325;
wire n_24;
wire n_328;
wire n_326;
wire n_332;
wire n_323;
wire n_319;
wire n_34;
wire n_33;
wire n_30;
wire n_31;
wire n_28;
wire n_285;
wire n_275;
wire n_35;
wire n_29;
wire n_284;
wire n_287;
wire n_277;
wire n_32;
wire n_286;
wire n_282;
wire n_279;
wire n_289;
wire n_63;
wire n_42;
wire n_41;
wire n_38;
wire n_39;
wire n_36;
wire n_313;
wire n_257;
wire n_43;
wire n_37;
wire n_312;
wire n_315;
wire n_259;
wire n_40;
wire n_314;
wire n_318;
wire n_261;
wire n_317;
wire n_61;
wire n_50;
wire n_49;
wire n_46;
wire n_47;
wire n_44;
wire n_296;
wire n_269;
wire n_51;
wire n_45;
wire n_295;
wire n_298;
wire n_271;
wire n_48;
wire n_297;
wire n_293;
wire n_273;
wire n_300;
wire n_59;
wire n_58;
wire n_57;
wire n_54;
wire n_55;
wire n_52;
wire n_305;
wire n_263;
wire n_65;
wire n_53;
wire n_304;
wire n_307;
wire n_266;
wire n_56;
wire n_306;
wire n_302;
wire n_267;
wire n_60;
wire n_268;
wire n_292;
wire n_62;
wire n_256;
wire n_310;
wire n_64;
wire n_274;
wire n_281;
wire n_308;
wire n_377;
wire n_373;
wire n_254;
wire n_72;
wire n_71;
wire n_68;
wire n_69;
wire n_66;
wire n_223;
wire n_213;
wire n_73;
wire n_67;
wire n_222;
wire n_225;
wire n_215;
wire n_70;
wire n_224;
wire n_220;
wire n_217;
wire n_227;
wire n_101;
wire n_80;
wire n_79;
wire n_76;
wire n_77;
wire n_74;
wire n_248;
wire n_206;
wire n_81;
wire n_75;
wire n_247;
wire n_250;
wire n_208;
wire n_78;
wire n_249;
wire n_253;
wire n_210;
wire n_252;
wire n_99;
wire n_88;
wire n_87;
wire n_84;
wire n_85;
wire n_82;
wire n_234;
wire n_192;
wire n_89;
wire n_83;
wire n_233;
wire n_236;
wire n_194;
wire n_86;
wire n_235;
wire n_231;
wire n_196;
wire n_238;
wire n_98;
wire n_97;
wire n_95;
wire n_94;
wire n_91;
wire n_90;
wire n_202;
wire n_242;
wire n_199;
wire n_103;
wire n_92;
wire n_93;
wire n_241;
wire n_200;
wire n_96;
wire n_243;
wire n_203;
wire n_204;
wire n_191;
wire n_230;
wire n_100;
wire n_205;
wire n_245;
wire n_102;
wire n_212;
wire n_219;
wire n_244;
wire n_189;
wire n_110;
wire n_109;
wire n_106;
wire n_107;
wire n_104;
wire n_186;
wire n_177;
wire n_111;
wire n_105;
wire n_187;
wire n_181;
wire n_108;
wire n_184;
wire n_182;
wire n_188;
wire n_179;
wire n_175;
wire n_118;
wire n_117;
wire n_114;
wire n_115;
wire n_112;
wire n_164;
wire n_154;
wire n_119;
wire n_113;
wire n_163;
wire n_166;
wire n_156;
wire n_116;
wire n_165;
wire n_161;
wire n_158;
wire n_168;
wire n_128;
wire n_127;
wire n_125;
wire n_124;
wire n_121;
wire n_120;
wire n_149;
wire n_172;
wire n_145;
wire n_129;
wire n_122;
wire n_123;
wire n_171;
wire n_146;
wire n_126;
wire n_173;
wire n_150;
wire n_151;
wire n_153;
wire n_160;
wire n_174;
wire n_143;
wire n_142;
wire n_140;
wire n_136;
wire n_141;
wire n_135;
wire n_131;
wire n_130;
wire n_137;
wire n_139;
wire n_133;
wire n_132;
wire n_134;
wire n_138;
wire n_379;
wire n_375;
wire n_371;
wire n_147;
wire n_144;
wire n_152;
wire n_159;
wire n_378;
wire n_374;
wire n_148;
wire n_170;
wire n_169;
wire n_155;
wire n_167;
wire n_162;
wire n_157;
wire n_176;
wire n_180;
wire n_183;
wire n_178;
wire n_185;
wire n_211;
wire n_190;
wire n_218;
wire n_197;
wire n_239;
wire n_229;
wire n_193;
wire n_237;
wire n_232;
wire n_195;
wire n_198;
wire n_201;
wire n_240;
wire n_207;
wire n_251;
wire n_246;
wire n_209;
wire n_228;
wire n_214;
wire n_226;
wire n_221;
wire n_216;
wire n_262;
wire n_255;
wire n_280;
wire n_290;
wire n_291;
wire n_301;
wire n_258;
wire n_316;
wire n_311;
wire n_260;
wire n_303;
wire n_265;
wire n_309;
wire n_264;
wire n_270;
wire n_299;
wire n_294;
wire n_272;
wire n_276;
wire n_288;
wire n_283;
wire n_278;
wire n_320;
wire n_324;
wire n_327;
wire n_322;
wire n_329;
wire n_334;
wire n_338;
wire n_341;
wire n_336;
wire n_343;
wire n_348;
wire n_352;
wire n_355;
wire n_350;
wire n_357;
wire n_362;
wire n_368;
wire n_367;


INV_X1 i_443 (.ZN (n_379), .A (p_0[61]));
INV_X1 i_442 (.ZN (n_378), .A (p_0[59]));
INV_X1 i_441 (.ZN (n_377), .A (p_0[31]));
INV_X1 i_440 (.ZN (n_376), .A (p_0[3]));
INV_X1 i_439 (.ZN (n_375), .A (tempResult[61]));
INV_X1 i_438 (.ZN (n_374), .A (tempResult[59]));
INV_X1 i_437 (.ZN (n_373), .A (tempResult[31]));
INV_X1 i_436 (.ZN (n_372), .A (tempResult[3]));
NOR2_X1 i_435 (.ZN (n_371), .A1 (p_0[60]), .A2 (tempResult[60]));
NAND2_X1 i_434 (.ZN (n_370), .A1 (n_376), .A2 (n_372));
NAND2_X1 i_433 (.ZN (n_369), .A1 (p_0[2]), .A2 (tempResult[2]));
INV_X1 i_432 (.ZN (n_368), .A (n_369));
NOR2_X1 i_431 (.ZN (n_367), .A1 (p_0[1]), .A2 (tempResult[1]));
NAND2_X1 i_430 (.ZN (n_366), .A1 (p_0[0]), .A2 (tempResult[0]));
NAND2_X1 i_429 (.ZN (n_365), .A1 (p_0[1]), .A2 (tempResult[1]));
AOI21_X1 i_428 (.ZN (n_364), .A (n_367), .B1 (n_366), .B2 (n_365));
OAI22_X2 i_427 (.ZN (n_363), .A1 (p_0[2]), .A2 (tempResult[2]), .B1 (n_368), .B2 (n_364));
OAI21_X1 i_426 (.ZN (n_362), .A (n_363), .B1 (n_376), .B2 (n_372));
NAND2_X1 i_425 (.ZN (n_361), .A1 (n_370), .A2 (n_362));
NOR2_X2 i_424 (.ZN (n_360), .A1 (p_0[7]), .A2 (tempResult[7]));
NOR2_X2 i_423 (.ZN (n_359), .A1 (p_0[5]), .A2 (tempResult[5]));
NOR2_X1 i_422 (.ZN (n_358), .A1 (p_0[6]), .A2 (tempResult[6]));
OR3_X1 i_421 (.ZN (n_357), .A1 (n_360), .A2 (n_358), .A3 (n_359));
NOR2_X1 i_420 (.ZN (n_356), .A1 (p_0[4]), .A2 (tempResult[4]));
NOR3_X1 i_419 (.ZN (n_355), .A1 (n_357), .A2 (n_356), .A3 (n_361));
NAND2_X1 i_418 (.ZN (n_354), .A1 (p_0[4]), .A2 (tempResult[4]));
NAND2_X1 i_417 (.ZN (n_353), .A1 (p_0[5]), .A2 (tempResult[5]));
AOI21_X1 i_416 (.ZN (n_352), .A (n_357), .B1 (n_354), .B2 (n_353));
AND2_X1 i_415 (.ZN (n_351), .A1 (p_0[7]), .A2 (tempResult[7]));
NAND2_X1 i_414 (.ZN (n_350), .A1 (p_0[6]), .A2 (tempResult[6]));
INV_X1 i_413 (.ZN (n_349), .A (n_350));
NOR2_X1 i_412 (.ZN (n_348), .A1 (n_360), .A2 (n_350));
NOR4_X2 i_411 (.ZN (n_347), .A1 (n_351), .A2 (n_348), .A3 (n_352), .A4 (n_355));
NOR2_X1 i_410 (.ZN (n_346), .A1 (p_0[11]), .A2 (tempResult[11]));
NOR2_X1 i_409 (.ZN (n_345), .A1 (p_0[9]), .A2 (tempResult[9]));
NOR2_X1 i_408 (.ZN (n_344), .A1 (p_0[10]), .A2 (tempResult[10]));
OR3_X1 i_407 (.ZN (n_343), .A1 (n_346), .A2 (n_344), .A3 (n_345));
NOR2_X1 i_406 (.ZN (n_342), .A1 (p_0[8]), .A2 (tempResult[8]));
NOR3_X1 i_405 (.ZN (n_341), .A1 (n_343), .A2 (n_342), .A3 (n_347));
NAND2_X1 i_404 (.ZN (n_340), .A1 (p_0[8]), .A2 (tempResult[8]));
NAND2_X1 i_403 (.ZN (n_339), .A1 (p_0[9]), .A2 (tempResult[9]));
AOI21_X1 i_402 (.ZN (n_338), .A (n_343), .B1 (n_340), .B2 (n_339));
AND2_X1 i_401 (.ZN (n_337), .A1 (p_0[11]), .A2 (tempResult[11]));
NAND2_X1 i_400 (.ZN (n_336), .A1 (p_0[10]), .A2 (tempResult[10]));
INV_X1 i_399 (.ZN (n_335), .A (n_336));
NOR2_X1 i_398 (.ZN (n_334), .A1 (n_346), .A2 (n_336));
NOR4_X2 i_397 (.ZN (n_333), .A1 (n_337), .A2 (n_334), .A3 (n_338), .A4 (n_341));
NOR2_X1 i_396 (.ZN (n_332), .A1 (p_0[15]), .A2 (tempResult[15]));
NOR2_X1 i_395 (.ZN (n_331), .A1 (p_0[13]), .A2 (tempResult[13]));
NOR2_X1 i_394 (.ZN (n_330), .A1 (p_0[14]), .A2 (tempResult[14]));
OR3_X1 i_393 (.ZN (n_329), .A1 (n_332), .A2 (n_330), .A3 (n_331));
NOR2_X1 i_392 (.ZN (n_328), .A1 (p_0[12]), .A2 (tempResult[12]));
NOR3_X1 i_391 (.ZN (n_327), .A1 (n_329), .A2 (n_328), .A3 (n_333));
NAND2_X1 i_390 (.ZN (n_326), .A1 (p_0[12]), .A2 (tempResult[12]));
NAND2_X1 i_389 (.ZN (n_325), .A1 (p_0[13]), .A2 (tempResult[13]));
AOI21_X1 i_388 (.ZN (n_324), .A (n_329), .B1 (n_326), .B2 (n_325));
AND2_X1 i_387 (.ZN (n_323), .A1 (p_0[15]), .A2 (tempResult[15]));
NAND2_X1 i_386 (.ZN (n_322), .A1 (p_0[14]), .A2 (tempResult[14]));
INV_X1 i_385 (.ZN (n_321), .A (n_322));
NOR2_X1 i_384 (.ZN (n_320), .A1 (n_332), .A2 (n_322));
NOR4_X4 i_383 (.ZN (n_319), .A1 (n_323), .A2 (n_320), .A3 (n_324), .A4 (n_327));
NOR2_X1 i_382 (.ZN (n_318), .A1 (p_0[20]), .A2 (tempResult[20]));
NOR2_X1 i_381 (.ZN (n_317), .A1 (p_0[23]), .A2 (tempResult[23]));
INV_X1 i_380 (.ZN (n_316), .A (n_317));
NOR2_X1 i_379 (.ZN (n_315), .A1 (p_0[21]), .A2 (tempResult[21]));
INV_X1 i_378 (.ZN (n_314), .A (n_315));
NOR2_X1 i_377 (.ZN (n_313), .A1 (p_0[22]), .A2 (tempResult[22]));
INV_X1 i_376 (.ZN (n_312), .A (n_313));
NAND3_X1 i_375 (.ZN (n_311), .A1 (n_316), .A2 (n_312), .A3 (n_314));
OR2_X1 i_374 (.ZN (n_310), .A1 (n_318), .A2 (n_311));
NOR2_X1 i_373 (.ZN (n_309), .A1 (p_0[31]), .A2 (tempResult[31]));
INV_X1 i_372 (.ZN (n_308), .A (n_309));
NOR2_X1 i_371 (.ZN (n_307), .A1 (p_0[29]), .A2 (tempResult[29]));
INV_X1 i_370 (.ZN (n_306), .A (n_307));
NOR2_X1 i_369 (.ZN (n_305), .A1 (p_0[30]), .A2 (tempResult[30]));
INV_X1 i_368 (.ZN (n_304), .A (n_305));
NAND3_X1 i_367 (.ZN (n_303), .A1 (n_308), .A2 (n_304), .A3 (n_306));
NOR2_X1 i_366 (.ZN (n_302), .A1 (p_0[28]), .A2 (tempResult[28]));
OR2_X1 i_365 (.ZN (n_301), .A1 (n_303), .A2 (n_302));
NOR2_X1 i_364 (.ZN (n_300), .A1 (p_0[27]), .A2 (tempResult[27]));
INV_X1 i_363 (.ZN (n_299), .A (n_300));
NOR2_X1 i_362 (.ZN (n_298), .A1 (p_0[25]), .A2 (tempResult[25]));
INV_X1 i_361 (.ZN (n_297), .A (n_298));
NOR2_X1 i_360 (.ZN (n_296), .A1 (p_0[26]), .A2 (tempResult[26]));
INV_X1 i_359 (.ZN (n_295), .A (n_296));
NAND3_X1 i_358 (.ZN (n_294), .A1 (n_299), .A2 (n_295), .A3 (n_297));
NOR2_X1 i_357 (.ZN (n_293), .A1 (p_0[24]), .A2 (tempResult[24]));
OR2_X1 i_356 (.ZN (n_292), .A1 (n_294), .A2 (n_293));
OR2_X1 i_355 (.ZN (n_291), .A1 (n_301), .A2 (n_292));
OR2_X1 i_354 (.ZN (n_290), .A1 (n_310), .A2 (n_291));
NOR2_X1 i_353 (.ZN (n_289), .A1 (p_0[19]), .A2 (tempResult[19]));
INV_X1 i_352 (.ZN (n_288), .A (n_289));
NOR2_X1 i_351 (.ZN (n_287), .A1 (p_0[17]), .A2 (tempResult[17]));
INV_X1 i_350 (.ZN (n_286), .A (n_287));
NOR2_X1 i_349 (.ZN (n_285), .A1 (p_0[18]), .A2 (tempResult[18]));
INV_X1 i_348 (.ZN (n_284), .A (n_285));
NAND3_X1 i_347 (.ZN (n_283), .A1 (n_288), .A2 (n_284), .A3 (n_286));
NOR2_X1 i_346 (.ZN (n_282), .A1 (p_0[16]), .A2 (tempResult[16]));
OR2_X1 i_345 (.ZN (n_281), .A1 (n_283), .A2 (n_282));
NOR3_X1 i_344 (.ZN (n_280), .A1 (n_290), .A2 (n_281), .A3 (n_319));
NAND2_X1 i_343 (.ZN (n_279), .A1 (p_0[16]), .A2 (tempResult[16]));
NAND2_X1 i_342 (.ZN (n_278), .A1 (p_0[17]), .A2 (tempResult[17]));
INV_X1 i_341 (.ZN (n_277), .A (n_278));
AOI21_X1 i_340 (.ZN (n_276), .A (n_283), .B1 (n_279), .B2 (n_278));
AND2_X1 i_339 (.ZN (n_275), .A1 (p_0[18]), .A2 (tempResult[18]));
AOI221_X1 i_338 (.ZN (n_274), .A (n_276), .B1 (p_0[19]), .B2 (tempResult[19]), .C1 (n_288), .C2 (n_275));
NAND2_X1 i_337 (.ZN (n_273), .A1 (p_0[24]), .A2 (tempResult[24]));
NAND2_X1 i_336 (.ZN (n_272), .A1 (p_0[25]), .A2 (tempResult[25]));
INV_X1 i_335 (.ZN (n_271), .A (n_272));
AOI21_X1 i_334 (.ZN (n_270), .A (n_294), .B1 (n_273), .B2 (n_272));
AND2_X1 i_333 (.ZN (n_269), .A1 (p_0[26]), .A2 (tempResult[26]));
AOI221_X1 i_332 (.ZN (n_268), .A (n_270), .B1 (p_0[27]), .B2 (tempResult[27]), .C1 (n_299), .C2 (n_269));
NAND2_X1 i_331 (.ZN (n_267), .A1 (p_0[28]), .A2 (tempResult[28]));
AND2_X1 i_330 (.ZN (n_266), .A1 (p_0[29]), .A2 (tempResult[29]));
AOI21_X1 i_329 (.ZN (n_265), .A (n_266), .B1 (p_0[28]), .B2 (tempResult[28]));
NAND2_X1 i_328 (.ZN (n_264), .A1 (p_0[30]), .A2 (tempResult[30]));
INV_X1 i_327 (.ZN (n_263), .A (n_264));
OAI222_X1 i_326 (.ZN (n_262), .A1 (n_303), .A2 (n_265), .B1 (n_309), .B2 (n_264), .C1 (n_377), .C2 (n_373));
NAND2_X1 i_325 (.ZN (n_261), .A1 (p_0[20]), .A2 (tempResult[20]));
NAND2_X1 i_324 (.ZN (n_260), .A1 (p_0[21]), .A2 (tempResult[21]));
INV_X1 i_323 (.ZN (n_259), .A (n_260));
AOI21_X1 i_322 (.ZN (n_258), .A (n_311), .B1 (n_261), .B2 (n_260));
AND2_X1 i_321 (.ZN (n_257), .A1 (p_0[22]), .A2 (tempResult[22]));
AOI221_X1 i_320 (.ZN (n_256), .A (n_258), .B1 (p_0[23]), .B2 (tempResult[23]), .C1 (n_316), .C2 (n_257));
OAI222_X1 i_319 (.ZN (n_255), .A1 (n_290), .A2 (n_274), .B1 (n_291), .B2 (n_256), .C1 (n_301), .C2 (n_268));
NOR3_X2 i_318 (.ZN (n_254), .A1 (n_262), .A2 (n_255), .A3 (n_280));
NOR2_X1 i_317 (.ZN (n_253), .A1 (p_0[36]), .A2 (tempResult[36]));
NOR2_X1 i_316 (.ZN (n_252), .A1 (p_0[39]), .A2 (tempResult[39]));
INV_X1 i_315 (.ZN (n_251), .A (n_252));
NOR2_X1 i_314 (.ZN (n_250), .A1 (p_0[37]), .A2 (tempResult[37]));
INV_X1 i_313 (.ZN (n_249), .A (n_250));
NOR2_X1 i_312 (.ZN (n_248), .A1 (p_0[38]), .A2 (tempResult[38]));
INV_X1 i_311 (.ZN (n_247), .A (n_248));
NAND3_X1 i_310 (.ZN (n_246), .A1 (n_251), .A2 (n_247), .A3 (n_249));
OR2_X1 i_309 (.ZN (n_245), .A1 (n_253), .A2 (n_246));
NOR2_X1 i_308 (.ZN (n_244), .A1 (p_0[47]), .A2 (tempResult[47]));
NOR2_X1 i_307 (.ZN (n_243), .A1 (p_0[45]), .A2 (tempResult[45]));
NOR2_X1 i_306 (.ZN (n_242), .A1 (p_0[46]), .A2 (tempResult[46]));
NOR2_X1 i_305 (.ZN (n_241), .A1 (n_243), .A2 (n_242));
NOR3_X1 i_304 (.ZN (n_240), .A1 (n_244), .A2 (n_242), .A3 (n_243));
OAI21_X1 i_303 (.ZN (n_239), .A (n_240), .B1 (p_0[44]), .B2 (tempResult[44]));
NOR2_X1 i_302 (.ZN (n_238), .A1 (p_0[43]), .A2 (tempResult[43]));
INV_X1 i_301 (.ZN (n_237), .A (n_238));
NOR2_X1 i_300 (.ZN (n_236), .A1 (p_0[41]), .A2 (tempResult[41]));
INV_X1 i_299 (.ZN (n_235), .A (n_236));
NOR2_X1 i_298 (.ZN (n_234), .A1 (p_0[42]), .A2 (tempResult[42]));
INV_X1 i_297 (.ZN (n_233), .A (n_234));
NAND3_X1 i_296 (.ZN (n_232), .A1 (n_237), .A2 (n_233), .A3 (n_235));
NOR2_X1 i_295 (.ZN (n_231), .A1 (p_0[40]), .A2 (tempResult[40]));
OR2_X1 i_294 (.ZN (n_230), .A1 (n_232), .A2 (n_231));
OR2_X1 i_293 (.ZN (n_229), .A1 (n_239), .A2 (n_230));
OR2_X1 i_292 (.ZN (n_228), .A1 (n_245), .A2 (n_229));
NOR2_X1 i_291 (.ZN (n_227), .A1 (p_0[35]), .A2 (tempResult[35]));
INV_X1 i_290 (.ZN (n_226), .A (n_227));
NOR2_X1 i_289 (.ZN (n_225), .A1 (p_0[33]), .A2 (tempResult[33]));
INV_X1 i_288 (.ZN (n_224), .A (n_225));
NOR2_X1 i_287 (.ZN (n_223), .A1 (p_0[34]), .A2 (tempResult[34]));
INV_X1 i_286 (.ZN (n_222), .A (n_223));
NAND3_X1 i_285 (.ZN (n_221), .A1 (n_226), .A2 (n_222), .A3 (n_224));
NOR2_X1 i_284 (.ZN (n_220), .A1 (p_0[32]), .A2 (tempResult[32]));
OR2_X1 i_283 (.ZN (n_219), .A1 (n_221), .A2 (n_220));
NOR3_X1 i_282 (.ZN (n_218), .A1 (n_228), .A2 (n_219), .A3 (n_254));
NAND2_X1 i_281 (.ZN (n_217), .A1 (p_0[32]), .A2 (tempResult[32]));
NAND2_X1 i_280 (.ZN (n_216), .A1 (p_0[33]), .A2 (tempResult[33]));
INV_X1 i_279 (.ZN (n_215), .A (n_216));
AOI21_X1 i_278 (.ZN (n_214), .A (n_221), .B1 (n_217), .B2 (n_216));
AND2_X1 i_277 (.ZN (n_213), .A1 (p_0[34]), .A2 (tempResult[34]));
AOI221_X1 i_276 (.ZN (n_212), .A (n_214), .B1 (p_0[35]), .B2 (tempResult[35]), .C1 (n_226), .C2 (n_213));
NOR2_X1 i_275 (.ZN (n_211), .A1 (n_228), .A2 (n_212));
NAND2_X1 i_274 (.ZN (n_210), .A1 (p_0[36]), .A2 (tempResult[36]));
NAND2_X1 i_273 (.ZN (n_209), .A1 (p_0[37]), .A2 (tempResult[37]));
INV_X1 i_272 (.ZN (n_208), .A (n_209));
AOI21_X1 i_271 (.ZN (n_207), .A (n_246), .B1 (n_210), .B2 (n_209));
AND2_X1 i_270 (.ZN (n_206), .A1 (p_0[38]), .A2 (tempResult[38]));
AOI221_X1 i_269 (.ZN (n_205), .A (n_207), .B1 (p_0[39]), .B2 (tempResult[39]), .C1 (n_251), .C2 (n_206));
NAND2_X1 i_268 (.ZN (n_204), .A1 (p_0[44]), .A2 (tempResult[44]));
INV_X1 i_267 (.ZN (n_203), .A (n_204));
AND2_X1 i_266 (.ZN (n_202), .A1 (p_0[45]), .A2 (tempResult[45]));
OAI21_X1 i_265 (.ZN (n_201), .A (n_240), .B1 (n_203), .B2 (n_202));
NAND2_X1 i_264 (.ZN (n_200), .A1 (p_0[46]), .A2 (tempResult[46]));
INV_X1 i_263 (.ZN (n_199), .A (n_200));
OAI21_X1 i_262 (.ZN (n_198), .A (n_201), .B1 (n_244), .B2 (n_200));
AOI21_X1 i_261 (.ZN (n_197), .A (n_198), .B1 (p_0[47]), .B2 (tempResult[47]));
NAND2_X1 i_260 (.ZN (n_196), .A1 (p_0[40]), .A2 (tempResult[40]));
NAND2_X1 i_259 (.ZN (n_195), .A1 (p_0[41]), .A2 (tempResult[41]));
INV_X1 i_258 (.ZN (n_194), .A (n_195));
AOI21_X1 i_257 (.ZN (n_193), .A (n_232), .B1 (n_196), .B2 (n_195));
AND2_X1 i_256 (.ZN (n_192), .A1 (p_0[42]), .A2 (tempResult[42]));
AOI221_X1 i_255 (.ZN (n_191), .A (n_193), .B1 (p_0[43]), .B2 (tempResult[43]), .C1 (n_237), .C2 (n_192));
OAI221_X1 i_254 (.ZN (n_190), .A (n_197), .B1 (n_239), .B2 (n_191), .C1 (n_229), .C2 (n_205));
NOR3_X2 i_253 (.ZN (n_189), .A1 (n_211), .A2 (n_190), .A3 (n_218));
NOR2_X1 i_252 (.ZN (n_188), .A1 (p_0[51]), .A2 (tempResult[51]));
NOR2_X1 i_251 (.ZN (n_187), .A1 (p_0[49]), .A2 (tempResult[49]));
NOR2_X1 i_250 (.ZN (n_186), .A1 (p_0[50]), .A2 (tempResult[50]));
OR3_X1 i_249 (.ZN (n_185), .A1 (n_188), .A2 (n_186), .A3 (n_187));
NOR2_X1 i_248 (.ZN (n_184), .A1 (p_0[48]), .A2 (tempResult[48]));
NOR3_X1 i_247 (.ZN (n_183), .A1 (n_185), .A2 (n_184), .A3 (n_189));
NAND2_X1 i_246 (.ZN (n_182), .A1 (p_0[48]), .A2 (tempResult[48]));
NAND2_X1 i_245 (.ZN (n_181), .A1 (p_0[49]), .A2 (tempResult[49]));
AOI21_X1 i_244 (.ZN (n_180), .A (n_185), .B1 (n_182), .B2 (n_181));
AND2_X1 i_243 (.ZN (n_179), .A1 (p_0[51]), .A2 (tempResult[51]));
NAND2_X1 i_242 (.ZN (n_178), .A1 (p_0[50]), .A2 (tempResult[50]));
INV_X1 i_241 (.ZN (n_177), .A (n_178));
NOR2_X1 i_240 (.ZN (n_176), .A1 (n_188), .A2 (n_178));
NOR4_X2 i_239 (.ZN (n_175), .A1 (n_179), .A2 (n_176), .A3 (n_180), .A4 (n_183));
NOR2_X1 i_238 (.ZN (n_174), .A1 (p_0[59]), .A2 (tempResult[59]));
NOR2_X1 i_237 (.ZN (n_173), .A1 (p_0[57]), .A2 (tempResult[57]));
NOR2_X1 i_236 (.ZN (n_172), .A1 (p_0[58]), .A2 (tempResult[58]));
NOR2_X1 i_235 (.ZN (n_171), .A1 (n_173), .A2 (n_172));
NOR3_X1 i_234 (.ZN (n_170), .A1 (n_174), .A2 (n_172), .A3 (n_173));
OAI21_X1 i_233 (.ZN (n_169), .A (n_170), .B1 (p_0[56]), .B2 (tempResult[56]));
NOR2_X1 i_232 (.ZN (n_168), .A1 (p_0[55]), .A2 (tempResult[55]));
INV_X1 i_231 (.ZN (n_167), .A (n_168));
NOR2_X1 i_230 (.ZN (n_166), .A1 (p_0[53]), .A2 (tempResult[53]));
INV_X1 i_229 (.ZN (n_165), .A (n_166));
NOR2_X1 i_228 (.ZN (n_164), .A1 (p_0[54]), .A2 (tempResult[54]));
INV_X1 i_227 (.ZN (n_163), .A (n_164));
NAND3_X1 i_226 (.ZN (n_162), .A1 (n_167), .A2 (n_163), .A3 (n_165));
NOR2_X1 i_225 (.ZN (n_161), .A1 (p_0[52]), .A2 (tempResult[52]));
OR2_X1 i_224 (.ZN (n_160), .A1 (n_162), .A2 (n_161));
NOR3_X1 i_223 (.ZN (n_159), .A1 (n_169), .A2 (n_160), .A3 (n_175));
NAND2_X1 i_222 (.ZN (n_158), .A1 (p_0[52]), .A2 (tempResult[52]));
NAND2_X1 i_221 (.ZN (n_157), .A1 (p_0[53]), .A2 (tempResult[53]));
INV_X1 i_220 (.ZN (n_156), .A (n_157));
AOI21_X1 i_219 (.ZN (n_155), .A (n_162), .B1 (n_158), .B2 (n_157));
AND2_X1 i_218 (.ZN (n_154), .A1 (p_0[54]), .A2 (tempResult[54]));
AOI221_X1 i_217 (.ZN (n_153), .A (n_155), .B1 (p_0[55]), .B2 (tempResult[55]), .C1 (n_167), .C2 (n_154));
NOR2_X1 i_216 (.ZN (n_152), .A1 (n_169), .A2 (n_153));
NAND2_X1 i_215 (.ZN (n_151), .A1 (p_0[56]), .A2 (tempResult[56]));
INV_X1 i_214 (.ZN (n_150), .A (n_151));
AND2_X1 i_213 (.ZN (n_149), .A1 (p_0[57]), .A2 (tempResult[57]));
OAI21_X1 i_212 (.ZN (n_148), .A (n_170), .B1 (n_150), .B2 (n_149));
INV_X1 i_211 (.ZN (n_147), .A (n_148));
NAND2_X1 i_210 (.ZN (n_146), .A1 (p_0[58]), .A2 (tempResult[58]));
INV_X1 i_209 (.ZN (n_145), .A (n_146));
OAI22_X1 i_208 (.ZN (n_144), .A1 (n_378), .A2 (n_374), .B1 (n_174), .B2 (n_146));
NOR4_X2 i_207 (.ZN (n_143), .A1 (n_147), .A2 (n_144), .A3 (n_152), .A4 (n_159));
AOI21_X1 i_206 (.ZN (n_142), .A (n_371), .B1 (p_0[60]), .B2 (tempResult[60]));
AOI21_X1 i_205 (.ZN (n_141), .A (n_371), .B1 (n_143), .B2 (n_142));
INV_X1 i_204 (.ZN (n_140), .A (n_141));
NAND2_X1 i_203 (.ZN (n_139), .A1 (p_0[62]), .A2 (tempResult[62]));
INV_X1 i_202 (.ZN (n_138), .A (n_139));
NAND2_X1 i_201 (.ZN (n_137), .A1 (n_379), .A2 (n_375));
OAI21_X1 i_200 (.ZN (n_136), .A (n_137), .B1 (n_379), .B2 (n_375));
INV_X1 i_199 (.ZN (n_135), .A (n_136));
NAND3_X1 i_198 (.ZN (n_134), .A1 (n_139), .A2 (n_135), .A3 (n_140));
OAI221_X1 i_197 (.ZN (n_133), .A (n_134), .B1 (p_0[62]), .B2 (tempResult[62]), .C1 (n_138), .C2 (n_137));
XNOR2_X1 i_196 (.ZN (n_132), .A (p_0[63]), .B (tempResult[63]));
XOR2_X1 i_195 (.Z (p_1[63]), .A (n_133), .B (n_132));
OAI21_X1 i_194 (.ZN (n_131), .A (n_139), .B1 (p_0[62]), .B2 (tempResult[62]));
AOI22_X1 i_193 (.ZN (n_130), .A1 (p_0[61]), .A2 (tempResult[61]), .B1 (n_141), .B2 (n_137));
XOR2_X1 i_192 (.Z (p_1[62]), .A (n_131), .B (n_130));
AOI22_X1 i_191 (.ZN (p_1[61]), .A1 (n_140), .A2 (n_136), .B1 (n_141), .B2 (n_135));
XNOR2_X1 i_190 (.ZN (p_1[60]), .A (n_143), .B (n_142));
AOI21_X1 i_189 (.ZN (n_129), .A (n_174), .B1 (p_0[59]), .B2 (tempResult[59]));
OAI21_X1 i_188 (.ZN (n_128), .A (n_153), .B1 (n_175), .B2 (n_160));
OAI21_X1 i_187 (.ZN (n_127), .A (n_151), .B1 (p_0[56]), .B2 (tempResult[56]));
OAI22_X1 i_186 (.ZN (n_126), .A1 (p_0[56]), .A2 (tempResult[56]), .B1 (n_150), .B2 (n_128));
INV_X1 i_185 (.ZN (n_125), .A (n_126));
NOR2_X1 i_184 (.ZN (n_124), .A1 (n_173), .A2 (n_149));
NAND3_X1 i_183 (.ZN (n_123), .A1 (n_146), .A2 (n_124), .A3 (n_126));
OAI21_X1 i_182 (.ZN (n_122), .A (n_123), .B1 (n_171), .B2 (n_145));
XNOR2_X1 i_181 (.ZN (p_1[59]), .A (n_129), .B (n_122));
NOR2_X1 i_180 (.ZN (n_121), .A1 (n_172), .A2 (n_145));
OAI22_X1 i_179 (.ZN (n_120), .A1 (p_0[57]), .A2 (tempResult[57]), .B1 (n_149), .B2 (n_125));
XNOR2_X1 i_178 (.ZN (p_1[58]), .A (n_121), .B (n_120));
XOR2_X1 i_177 (.Z (p_1[57]), .A (n_125), .B (n_124));
XNOR2_X1 i_176 (.ZN (p_1[56]), .A (n_128), .B (n_127));
AOI21_X1 i_175 (.ZN (n_119), .A (n_168), .B1 (p_0[55]), .B2 (tempResult[55]));
OAI21_X1 i_174 (.ZN (n_118), .A (n_158), .B1 (p_0[52]), .B2 (tempResult[52]));
AOI21_X1 i_173 (.ZN (n_117), .A (n_161), .B1 (n_175), .B2 (n_158));
OAI21_X1 i_172 (.ZN (n_116), .A (n_165), .B1 (n_156), .B2 (n_117));
INV_X1 i_171 (.ZN (n_115), .A (n_116));
NOR2_X1 i_170 (.ZN (n_114), .A1 (n_166), .A2 (n_156));
OAI21_X1 i_169 (.ZN (n_113), .A (n_163), .B1 (n_154), .B2 (n_115));
XNOR2_X1 i_168 (.ZN (p_1[55]), .A (n_119), .B (n_113));
NOR2_X1 i_167 (.ZN (n_112), .A1 (n_164), .A2 (n_154));
XOR2_X1 i_166 (.Z (p_1[54]), .A (n_115), .B (n_112));
XOR2_X1 i_165 (.Z (p_1[53]), .A (n_117), .B (n_114));
XOR2_X1 i_164 (.Z (p_1[52]), .A (n_175), .B (n_118));
NOR2_X1 i_163 (.ZN (n_111), .A1 (n_188), .A2 (n_179));
OAI21_X1 i_162 (.ZN (n_110), .A (n_182), .B1 (p_0[48]), .B2 (tempResult[48]));
AOI21_X1 i_161 (.ZN (n_109), .A (n_184), .B1 (n_189), .B2 (n_182));
INV_X1 i_160 (.ZN (n_108), .A (n_109));
AOI21_X1 i_159 (.ZN (n_107), .A (n_187), .B1 (n_181), .B2 (n_108));
AOI21_X1 i_158 (.ZN (n_106), .A (n_187), .B1 (p_0[49]), .B2 (tempResult[49]));
OAI22_X1 i_157 (.ZN (n_105), .A1 (p_0[50]), .A2 (tempResult[50]), .B1 (n_177), .B2 (n_107));
XNOR2_X1 i_156 (.ZN (p_1[51]), .A (n_111), .B (n_105));
NOR2_X1 i_155 (.ZN (n_104), .A1 (n_186), .A2 (n_177));
XOR2_X1 i_154 (.Z (p_1[50]), .A (n_107), .B (n_104));
XOR2_X1 i_153 (.Z (p_1[49]), .A (n_109), .B (n_106));
XOR2_X1 i_152 (.Z (p_1[48]), .A (n_189), .B (n_110));
AOI21_X1 i_151 (.ZN (n_103), .A (n_244), .B1 (p_0[47]), .B2 (tempResult[47]));
OAI21_X1 i_150 (.ZN (n_102), .A (n_212), .B1 (n_254), .B2 (n_219));
INV_X1 i_149 (.ZN (n_101), .A (n_102));
OAI21_X1 i_148 (.ZN (n_100), .A (n_205), .B1 (n_245), .B2 (n_101));
INV_X1 i_147 (.ZN (n_99), .A (n_100));
OAI21_X1 i_146 (.ZN (n_98), .A (n_191), .B1 (n_230), .B2 (n_99));
OAI21_X1 i_145 (.ZN (n_97), .A (n_204), .B1 (p_0[44]), .B2 (tempResult[44]));
OAI22_X1 i_144 (.ZN (n_96), .A1 (p_0[44]), .A2 (tempResult[44]), .B1 (n_203), .B2 (n_98));
INV_X1 i_143 (.ZN (n_95), .A (n_96));
NOR2_X1 i_142 (.ZN (n_94), .A1 (n_243), .A2 (n_202));
NAND3_X1 i_141 (.ZN (n_93), .A1 (n_200), .A2 (n_94), .A3 (n_96));
OAI21_X1 i_140 (.ZN (n_92), .A (n_93), .B1 (n_241), .B2 (n_199));
XNOR2_X1 i_139 (.ZN (p_1[47]), .A (n_103), .B (n_92));
NOR2_X1 i_138 (.ZN (n_91), .A1 (n_242), .A2 (n_199));
OAI22_X1 i_137 (.ZN (n_90), .A1 (p_0[45]), .A2 (tempResult[45]), .B1 (n_202), .B2 (n_95));
XNOR2_X1 i_136 (.ZN (p_1[46]), .A (n_91), .B (n_90));
XOR2_X1 i_135 (.Z (p_1[45]), .A (n_95), .B (n_94));
XNOR2_X1 i_134 (.ZN (p_1[44]), .A (n_98), .B (n_97));
AOI21_X1 i_133 (.ZN (n_89), .A (n_238), .B1 (p_0[43]), .B2 (tempResult[43]));
OAI21_X1 i_132 (.ZN (n_88), .A (n_196), .B1 (p_0[40]), .B2 (tempResult[40]));
AOI21_X1 i_131 (.ZN (n_87), .A (n_231), .B1 (n_196), .B2 (n_99));
OAI21_X1 i_130 (.ZN (n_86), .A (n_235), .B1 (n_194), .B2 (n_87));
INV_X1 i_129 (.ZN (n_85), .A (n_86));
NOR2_X1 i_128 (.ZN (n_84), .A1 (n_236), .A2 (n_194));
OAI21_X1 i_127 (.ZN (n_83), .A (n_233), .B1 (n_192), .B2 (n_85));
XNOR2_X1 i_126 (.ZN (p_1[43]), .A (n_89), .B (n_83));
NOR2_X1 i_125 (.ZN (n_82), .A1 (n_234), .A2 (n_192));
XOR2_X1 i_124 (.Z (p_1[42]), .A (n_85), .B (n_82));
XOR2_X1 i_123 (.Z (p_1[41]), .A (n_87), .B (n_84));
XOR2_X1 i_122 (.Z (p_1[40]), .A (n_99), .B (n_88));
AOI21_X1 i_121 (.ZN (n_81), .A (n_252), .B1 (p_0[39]), .B2 (tempResult[39]));
OAI21_X1 i_120 (.ZN (n_80), .A (n_210), .B1 (p_0[36]), .B2 (tempResult[36]));
AOI21_X1 i_119 (.ZN (n_79), .A (n_253), .B1 (n_210), .B2 (n_101));
OAI21_X1 i_118 (.ZN (n_78), .A (n_249), .B1 (n_208), .B2 (n_79));
INV_X1 i_117 (.ZN (n_77), .A (n_78));
NOR2_X1 i_116 (.ZN (n_76), .A1 (n_250), .A2 (n_208));
OAI21_X1 i_115 (.ZN (n_75), .A (n_247), .B1 (n_206), .B2 (n_77));
XNOR2_X1 i_114 (.ZN (p_1[39]), .A (n_81), .B (n_75));
NOR2_X1 i_113 (.ZN (n_74), .A1 (n_248), .A2 (n_206));
XOR2_X1 i_112 (.Z (p_1[38]), .A (n_77), .B (n_74));
XOR2_X1 i_111 (.Z (p_1[37]), .A (n_79), .B (n_76));
XOR2_X1 i_110 (.Z (p_1[36]), .A (n_101), .B (n_80));
AOI21_X1 i_109 (.ZN (n_73), .A (n_227), .B1 (p_0[35]), .B2 (tempResult[35]));
OAI21_X1 i_108 (.ZN (n_72), .A (n_217), .B1 (p_0[32]), .B2 (tempResult[32]));
AOI21_X1 i_107 (.ZN (n_71), .A (n_220), .B1 (n_254), .B2 (n_217));
OAI21_X1 i_106 (.ZN (n_70), .A (n_224), .B1 (n_215), .B2 (n_71));
INV_X1 i_105 (.ZN (n_69), .A (n_70));
NOR2_X1 i_104 (.ZN (n_68), .A1 (n_225), .A2 (n_215));
OAI21_X1 i_103 (.ZN (n_67), .A (n_222), .B1 (n_213), .B2 (n_69));
XNOR2_X1 i_102 (.ZN (p_1[35]), .A (n_73), .B (n_67));
NOR2_X1 i_101 (.ZN (n_66), .A1 (n_223), .A2 (n_213));
XOR2_X1 i_100 (.Z (p_1[34]), .A (n_69), .B (n_66));
XOR2_X1 i_99 (.Z (p_1[33]), .A (n_71), .B (n_68));
XOR2_X1 i_98 (.Z (p_1[32]), .A (n_254), .B (n_72));
OAI21_X1 i_97 (.ZN (n_65), .A (n_308), .B1 (n_377), .B2 (n_373));
OAI21_X1 i_96 (.ZN (n_64), .A (n_274), .B1 (n_319), .B2 (n_281));
INV_X1 i_95 (.ZN (n_63), .A (n_64));
OAI21_X1 i_94 (.ZN (n_62), .A (n_256), .B1 (n_310), .B2 (n_63));
INV_X1 i_93 (.ZN (n_61), .A (n_62));
OAI21_X1 i_92 (.ZN (n_60), .A (n_268), .B1 (n_292), .B2 (n_61));
INV_X1 i_91 (.ZN (n_59), .A (n_60));
OAI21_X1 i_90 (.ZN (n_58), .A (n_267), .B1 (p_0[28]), .B2 (tempResult[28]));
AOI21_X1 i_89 (.ZN (n_57), .A (n_302), .B1 (n_267), .B2 (n_59));
OAI21_X1 i_88 (.ZN (n_56), .A (n_306), .B1 (n_266), .B2 (n_57));
INV_X1 i_87 (.ZN (n_55), .A (n_56));
NOR2_X1 i_86 (.ZN (n_54), .A1 (n_307), .A2 (n_266));
OAI21_X1 i_85 (.ZN (n_53), .A (n_304), .B1 (n_263), .B2 (n_55));
XOR2_X1 i_84 (.Z (p_1[31]), .A (n_65), .B (n_53));
NOR2_X1 i_83 (.ZN (n_52), .A1 (n_305), .A2 (n_263));
XOR2_X1 i_82 (.Z (p_1[30]), .A (n_55), .B (n_52));
XOR2_X1 i_81 (.Z (p_1[29]), .A (n_57), .B (n_54));
XOR2_X1 i_80 (.Z (p_1[28]), .A (n_59), .B (n_58));
AOI21_X1 i_79 (.ZN (n_51), .A (n_300), .B1 (p_0[27]), .B2 (tempResult[27]));
OAI21_X1 i_78 (.ZN (n_50), .A (n_273), .B1 (p_0[24]), .B2 (tempResult[24]));
AOI21_X1 i_77 (.ZN (n_49), .A (n_293), .B1 (n_273), .B2 (n_61));
OAI21_X1 i_76 (.ZN (n_48), .A (n_297), .B1 (n_271), .B2 (n_49));
INV_X1 i_75 (.ZN (n_47), .A (n_48));
NOR2_X1 i_74 (.ZN (n_46), .A1 (n_298), .A2 (n_271));
OAI21_X1 i_73 (.ZN (n_45), .A (n_295), .B1 (n_269), .B2 (n_47));
XNOR2_X1 i_72 (.ZN (p_1[27]), .A (n_51), .B (n_45));
NOR2_X1 i_71 (.ZN (n_44), .A1 (n_296), .A2 (n_269));
XOR2_X1 i_70 (.Z (p_1[26]), .A (n_47), .B (n_44));
XOR2_X1 i_69 (.Z (p_1[25]), .A (n_49), .B (n_46));
XOR2_X1 i_68 (.Z (p_1[24]), .A (n_61), .B (n_50));
AOI21_X1 i_67 (.ZN (n_43), .A (n_317), .B1 (p_0[23]), .B2 (tempResult[23]));
OAI21_X1 i_66 (.ZN (n_42), .A (n_261), .B1 (p_0[20]), .B2 (tempResult[20]));
AOI21_X1 i_65 (.ZN (n_41), .A (n_318), .B1 (n_261), .B2 (n_63));
OAI21_X1 i_64 (.ZN (n_40), .A (n_314), .B1 (n_259), .B2 (n_41));
INV_X1 i_63 (.ZN (n_39), .A (n_40));
NOR2_X1 i_62 (.ZN (n_38), .A1 (n_315), .A2 (n_259));
OAI21_X1 i_61 (.ZN (n_37), .A (n_312), .B1 (n_257), .B2 (n_39));
XNOR2_X1 i_60 (.ZN (p_1[23]), .A (n_43), .B (n_37));
NOR2_X1 i_59 (.ZN (n_36), .A1 (n_313), .A2 (n_257));
XOR2_X1 i_58 (.Z (p_1[22]), .A (n_39), .B (n_36));
XOR2_X1 i_57 (.Z (p_1[21]), .A (n_41), .B (n_38));
XOR2_X1 i_56 (.Z (p_1[20]), .A (n_63), .B (n_42));
AOI21_X1 i_55 (.ZN (n_35), .A (n_289), .B1 (p_0[19]), .B2 (tempResult[19]));
OAI21_X1 i_54 (.ZN (n_34), .A (n_279), .B1 (p_0[16]), .B2 (tempResult[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_282), .B1 (n_319), .B2 (n_279));
OAI21_X1 i_52 (.ZN (n_32), .A (n_286), .B1 (n_277), .B2 (n_33));
INV_X1 i_51 (.ZN (n_31), .A (n_32));
NOR2_X1 i_50 (.ZN (n_30), .A1 (n_287), .A2 (n_277));
OAI21_X1 i_49 (.ZN (n_29), .A (n_284), .B1 (n_275), .B2 (n_31));
XNOR2_X1 i_48 (.ZN (p_1[19]), .A (n_35), .B (n_29));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_285), .A2 (n_275));
XOR2_X1 i_46 (.Z (p_1[18]), .A (n_31), .B (n_28));
XOR2_X1 i_45 (.Z (p_1[17]), .A (n_33), .B (n_30));
XOR2_X1 i_44 (.Z (p_1[16]), .A (n_319), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_332), .A2 (n_323));
OAI21_X1 i_42 (.ZN (n_26), .A (n_326), .B1 (p_0[12]), .B2 (tempResult[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_328), .B1 (n_333), .B2 (n_326));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_331), .B1 (n_325), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_331), .B1 (p_0[13]), .B2 (tempResult[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (p_0[14]), .A2 (tempResult[14]), .B1 (n_321), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (p_1[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_330), .A2 (n_321));
XOR2_X1 i_34 (.Z (p_1[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (p_1[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (p_1[12]), .A (n_333), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_346), .A2 (n_337));
AOI21_X1 i_30 (.ZN (n_18), .A (n_342), .B1 (p_0[8]), .B2 (tempResult[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_342), .B1 (n_347), .B2 (n_340));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_345), .B1 (n_339), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_345), .B1 (p_0[9]), .B2 (tempResult[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (p_0[10]), .A2 (tempResult[10]), .B1 (n_335), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (p_1[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_344), .A2 (n_335));
XOR2_X1 i_22 (.Z (p_1[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (p_1[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (p_1[8]), .A (n_347), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_360), .A2 (n_351));
OAI21_X1 i_18 (.ZN (n_10), .A (n_354), .B1 (p_0[4]), .B2 (tempResult[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_356), .B1 (n_361), .B2 (n_354));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_359), .B1 (n_353), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_359), .B1 (p_0[5]), .B2 (tempResult[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (p_0[6]), .A2 (tempResult[6]), .B1 (n_349), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (p_1[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_358), .A2 (n_349));
XOR2_X1 i_10 (.Z (p_1[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (p_1[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (p_1[4]), .A (n_361), .B (n_10));
OAI21_X1 i_7 (.ZN (n_3), .A (n_370), .B1 (n_376), .B2 (n_372));
XOR2_X1 i_6 (.Z (p_1[3]), .A (n_363), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_369), .B1 (p_0[2]), .B2 (tempResult[2]));
XNOR2_X1 i_4 (.ZN (p_1[2]), .A (n_364), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_365), .B1 (p_0[1]), .B2 (tempResult[1]));
XOR2_X1 i_2 (.Z (p_1[1]), .A (n_366), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_366), .B1 (p_0[0]), .B2 (tempResult[0]));
INV_X1 i_0 (.ZN (p_1[0]), .A (n_0));

endmodule //datapath__0_12

module datapath__0_0 (p_0, p_1);

output [32:0] p_0;
input [32:0] p_1;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (p_1[26]));
INV_X1 i_63 (.ZN (n_32), .A (p_1[22]));
INV_X1 i_62 (.ZN (n_31), .A (p_1[15]));
INV_X1 i_61 (.ZN (n_30), .A (p_1[12]));
OR3_X1 i_60 (.ZN (n_29), .A1 (p_1[3]), .A2 (p_1[2]), .A3 (p_1[1]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (p_1[4]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (p_1[5]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (p_1[6]), .A3 (p_1[7]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (p_1[8]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (p_1[9]), .A3 (p_1[10]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (p_1[11]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (p_1[13]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (p_1[13]), .A3 (p_1[14]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (p_1[16]), .A3 (p_1[17]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (p_1[18]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (p_1[19]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (p_1[19]), .A3 (p_1[20]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (p_1[19]), .A3 (p_1[20]), .A4 (p_1[21]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (p_1[23]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (p_1[24]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (p_1[24]), .A3 (p_1[25]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (p_1[27]), .A3 (p_1[28]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (p_1[29]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (p_1[29]), .A3 (p_1[30]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (p_1[29]), .A3 (p_1[30]), .A4 (p_1[31]));
XNOR2_X1 i_35 (.ZN (p_0[32]), .A (p_1[32]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[31]), .A (p_1[31]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[30]), .A (p_1[30]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[29]), .A (p_1[29]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (p_1[28]), .B1 (n_9), .B2 (p_1[27]));
AND2_X1 i_30 (.ZN (p_0[28]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[27]), .A (p_1[27]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[26]), .A (p_1[26]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[25]), .A (p_1[25]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[24]), .A (p_1[24]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[23]), .A (p_1[23]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[22]), .A (p_1[22]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[21]), .A (p_1[21]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[20]), .A (p_1[20]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[19]), .A (p_1[19]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[18]), .A (p_1[18]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (p_1[17]), .B1 (n_19), .B2 (p_1[16]));
AND2_X1 i_18 (.ZN (p_0[17]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[16]), .A (p_1[16]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[15]), .A (p_1[15]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[14]), .A (p_1[14]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[13]), .A (p_1[13]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[12]), .A (p_1[12]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[11]), .A (p_1[11]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (p_1[10]), .B1 (n_25), .B2 (p_1[9]));
AND2_X1 i_10 (.ZN (p_0[10]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[9]), .A (p_1[9]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[8]), .A (p_1[8]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (p_1[7]), .B1 (n_27), .B2 (p_1[6]));
AND2_X1 i_6 (.ZN (p_0[7]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[6]), .A (p_1[6]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[5]), .A (p_1[5]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[4]), .A (p_1[4]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (p_1[3]), .B1 (p_1[2]), .B2 (p_1[1]));
AND2_X1 i_1 (.ZN (p_0[3]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[2]), .A (p_1[2]), .B (p_1[1]));

endmodule //datapath__0_0

module Noaman_4_Booth (clk_CTS_1_PP_2, CTSclk_CTS_1_PP_2PP_0, start, clk, in1, in2, 
    result);

output [63:0] result;
input clk;
input [31:0] in1;
input [31:0] in2;
input start;
input clk_CTS_1_PP_2;
input CTSclk_CTS_1_PP_2PP_0;
wire CLOCK_slh_n239;
wire n_0_3;
wire n_0_0;
wire n_0_4;
wire n_0_1;
wire n_0_5;
wire n_0_2;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_316__0;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_318__0;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_320__0;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_321__0;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_322__0;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_323__0;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_324__0;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_325__0;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_326__0;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_327__0;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_328__0;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_329__0;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_330__0;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_331__0;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_332__0;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_333__0;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_334__0;
wire n_0_185;
wire n_0_186;
wire n_0_187;
wire n_0_188;
wire n_0_189;
wire n_0_190;
wire n_0_335__0;
wire n_0_191;
wire n_0_192;
wire n_0_193;
wire n_0_194;
wire n_0_195;
wire n_0_196;
wire n_0_336__0;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_201;
wire n_0_202;
wire n_0_337__0;
wire n_0_203;
wire n_0_204;
wire n_0_205;
wire n_0_206;
wire n_0_207;
wire n_0_208;
wire n_0_338__0;
wire n_0_209;
wire n_0_210;
wire n_0_211;
wire n_0_212;
wire n_0_213;
wire n_0_214;
wire n_0_339__0;
wire n_0_215;
wire n_0_216;
wire n_0_217;
wire n_0_218;
wire n_0_219;
wire n_0_220;
wire n_0_340__0;
wire n_0_221;
wire n_0_222;
wire n_0_223;
wire n_0_224;
wire n_0_225;
wire n_0_226;
wire n_0_341__0;
wire n_0_227;
wire n_0_228;
wire n_0_229;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_342__0;
wire n_0_233;
wire n_0_234;
wire n_0_235;
wire n_0_236;
wire n_0_237;
wire n_0_238;
wire n_0_343__0;
wire n_0_239;
wire n_0_240;
wire n_0_241;
wire n_0_242;
wire n_0_243;
wire n_0_244;
wire n_0_344__0;
wire n_0_245;
wire n_0_246;
wire n_0_247;
wire n_0_248;
wire n_0_249;
wire n_0_250;
wire n_0_345__0;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_346__0;
wire n_0_257;
wire n_0_258;
wire n_0_259;
wire n_0_260;
wire n_0_261;
wire n_0_262;
wire n_0_347__0;
wire n_0_263;
wire n_0_264;
wire n_0_265;
wire n_0_266;
wire n_0_267;
wire n_0_268;
wire n_0_348__0;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_272;
wire n_0_273;
wire n_0_274;
wire n_0_349__0;
wire n_0_275;
wire n_0_276;
wire n_0_277;
wire n_0_278;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_350__0;
wire n_0_282;
wire n_0_283;
wire n_0_284;
wire n_0_351__0;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_288;
wire n_0_352__0;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_353__0;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_354__0;
wire n_0_296;
wire n_0_297;
wire n_0_298;
wire n_0_355__0;
wire n_0_299;
wire n_0_300;
wire n_0_301;
wire n_0_302;
wire n_0_356__0;
wire n_0_303;
wire n_0_304;
wire n_0_305;
wire n_0_306;
wire n_0_357__0;
wire n_0_307;
wire n_0_308;
wire n_0_309;
wire n_0_358__0;
wire n_0_310;
wire n_0_311;
wire n_0_312;
wire n_0_359__0;
wire n_0_313;
wire n_0_314;
wire n_0_315;
wire n_0_360__0;
wire n_0_316__1;
wire n_0_317;
wire n_0_318__1;
wire n_0_361__0;
wire n_0_319;
wire n_0_320__1;
wire n_0_321__1;
wire n_0_362__0;
wire n_0_322__1;
wire n_0_323__1;
wire n_0_324__1;
wire n_0_363__0;
wire n_0_325__1;
wire n_0_326__1;
wire n_0_327__1;
wire n_0_364__0;
wire n_0_328__1;
wire n_0_329__1;
wire n_0_330__1;
wire n_0_365__0;
wire n_0_331__1;
wire n_0_332__1;
wire n_0_333__1;
wire n_0_334__1;
wire n_0_335__1;
wire n_0_366__0;
wire n_0_336__1;
wire n_0_337__1;
wire n_0_338__1;
wire n_0_367__0;
wire n_0_339__1;
wire n_0_340__1;
wire n_0_341__1;
wire n_0_368__0;
wire n_0_342__1;
wire n_0_343__1;
wire n_0_344__1;
wire n_0_369__0;
wire n_0_345__1;
wire n_0_346__1;
wire n_0_347__1;
wire n_0_370__0;
wire n_0_348__1;
wire n_0_349__1;
wire n_0_350__1;
wire n_0_371__0;
wire n_0_351__1;
wire n_0_352__1;
wire n_0_353__1;
wire n_0_372;
wire n_0_354__1;
wire n_0_355__1;
wire n_0_356__1;
wire n_0_373;
wire n_0_357__1;
wire n_0_358__1;
wire n_0_359__1;
wire n_0_374;
wire n_0_360__1;
wire n_0_361__1;
wire n_0_362__1;
wire n_0_375;
wire n_0_363__1;
wire n_0_364__1;
wire n_0_365__1;
wire n_0_376;
wire n_0_366__1;
wire n_0_367__1;
wire n_0_368__1;
wire n_0_377;
wire n_0_369__1;
wire n_0_381;
wire n_0_370__1;
wire n_0_378;
wire n_0_379;
wire n_0_371__1;
wire n_0_380;
wire \tempResult[63] ;
wire \tempResult[62] ;
wire \tempResult[61] ;
wire \tempResult[60] ;
wire \tempResult[59] ;
wire \tempResult[58] ;
wire \tempResult[57] ;
wire \tempResult[56] ;
wire \tempResult[55] ;
wire \tempResult[54] ;
wire \tempResult[53] ;
wire \tempResult[52] ;
wire \tempResult[51] ;
wire \tempResult[50] ;
wire \tempResult[49] ;
wire \tempResult[48] ;
wire \tempResult[47] ;
wire \tempResult[46] ;
wire \tempResult[45] ;
wire \tempResult[44] ;
wire \tempResult[43] ;
wire \tempResult[42] ;
wire \tempResult[41] ;
wire \tempResult[40] ;
wire \tempResult[39] ;
wire \tempResult[38] ;
wire \tempResult[37] ;
wire \tempResult[36] ;
wire \tempResult[35] ;
wire \tempResult[34] ;
wire \tempResult[33] ;
wire \tempResult[32] ;
wire \tempResult[31] ;
wire \tempResult[30] ;
wire \tempResult[29] ;
wire \tempResult[28] ;
wire \tempResult[27] ;
wire \tempResult[26] ;
wire \tempResult[25] ;
wire \tempResult[24] ;
wire \tempResult[23] ;
wire \tempResult[22] ;
wire \tempResult[21] ;
wire \tempResult[20] ;
wire \tempResult[19] ;
wire \tempResult[18] ;
wire \tempResult[17] ;
wire \tempResult[16] ;
wire \tempResult[15] ;
wire \tempResult[14] ;
wire \tempResult[13] ;
wire \tempResult[12] ;
wire \tempResult[11] ;
wire \tempResult[10] ;
wire \tempResult[9] ;
wire \tempResult[8] ;
wire \tempResult[7] ;
wire \tempResult[6] ;
wire \tempResult[5] ;
wire \tempResult[4] ;
wire \tempResult[3] ;
wire \tempResult[2] ;
wire \tempResult[1] ;
wire \tempResult[0] ;
wire \shiftingAmount[5] ;
wire \shiftingAmount[4] ;
wire \shiftingAmount[3] ;
wire \shiftingAmount[2] ;
wire \shiftingAmount[1] ;
wire \newB[34] ;
wire \newB[31] ;
wire \newB[30] ;
wire \newB[29] ;
wire \newB[28] ;
wire \newB[27] ;
wire \newB[26] ;
wire \newB[25] ;
wire \newB[24] ;
wire \newB[23] ;
wire \newB[22] ;
wire \newB[21] ;
wire \newB[20] ;
wire \newB[19] ;
wire \newB[18] ;
wire \newB[17] ;
wire \newB[16] ;
wire \newB[15] ;
wire \newB[14] ;
wire \newB[13] ;
wire \newB[12] ;
wire \newB[11] ;
wire \newB[10] ;
wire \newB[9] ;
wire \newB[8] ;
wire \newB[7] ;
wire \newB[6] ;
wire \newB[5] ;
wire \newB[4] ;
wire \newB[3] ;
wire \newB[2] ;
wire \newB[1] ;
wire \Input1_1_Negative[63] ;
wire \Input1_1_Negative[29] ;
wire \Input1_1_Negative[27] ;
wire \Input1_1_Negative[25] ;
wire \Input1_1_Negative[23] ;
wire \Input1_1_Negative[21] ;
wire \Input1_1_Negative[19] ;
wire \Input1_1_Negative[17] ;
wire \Input1_1_Negative[15] ;
wire \Input1_1_Negative[13] ;
wire \Input1_1_Negative[11] ;
wire \Input1_1_Negative[9] ;
wire \Input1_1_Negative[7] ;
wire \Input1_1_Negative[5] ;
wire \Input1_1_Negative[3] ;
wire \Input1_1_Negative[1] ;
wire \Input1_1_Positive[63] ;
wire \Input1_1_Positive[29] ;
wire \Input1_1_Positive[27] ;
wire \Input1_1_Positive[25] ;
wire \Input1_1_Positive[23] ;
wire \Input1_1_Positive[21] ;
wire \Input1_1_Positive[19] ;
wire \Input1_1_Positive[17] ;
wire \Input1_1_Positive[15] ;
wire \Input1_1_Positive[13] ;
wire \Input1_1_Positive[11] ;
wire \Input1_1_Positive[9] ;
wire \Input1_1_Positive[7] ;
wire \Input1_1_Positive[5] ;
wire \Input1_1_Positive[3] ;
wire \Input1_1_Positive[1] ;
wire \Input1_2_Negative[31] ;
wire \Input1_2_Negative[29] ;
wire \Input1_2_Negative[27] ;
wire \Input1_2_Negative[25] ;
wire \Input1_2_Negative[23] ;
wire \Input1_2_Negative[21] ;
wire \Input1_2_Negative[19] ;
wire \Input1_2_Negative[17] ;
wire \Input1_2_Negative[15] ;
wire \Input1_2_Negative[13] ;
wire \Input1_2_Negative[11] ;
wire \Input1_2_Negative[9] ;
wire \Input1_2_Negative[7] ;
wire \Input1_2_Negative[5] ;
wire \Input1_2_Negative[3] ;
wire n_tid1_233;
wire CTS_n_tid1_133;
wire CTS_n_tid0_105;
wire \Input1_2_Positive[31] ;
wire CTS_n_tid0_143;
wire \Input1_2_Positive[29] ;
wire \Input1_2_Positive[27] ;
wire \Input1_2_Positive[25] ;
wire CTS_n_tid1_42;
wire \Input1_2_Positive[23] ;
wire drc_ipo_n34;
wire \Input1_2_Positive[21] ;
wire CTS_n_tid1_41;
wire \Input1_2_Positive[19] ;
wire drc_ipo_n33;
wire \Input1_2_Positive[17] ;
wire hfn_ipo_n30;
wire \Input1_2_Positive[15] ;
wire hfn_ipo_n29;
wire \Input1_2_Positive[13] ;
wire hfn_ipo_n26;
wire \Input1_2_Positive[11] ;
wire hfn_ipo_n32;
wire \Input1_2_Positive[9] ;
wire hfn_ipo_n31;
wire \Input1_2_Positive[7] ;
wire hfn_ipo_n28;
wire \Input1_2_Positive[5] ;
wire hfn_ipo_n27;
wire \Input1_2_Positive[3] ;
wire hfn_ipo_n24;
wire \Input1_2_Positive[1] ;
wire hfn_ipo_n23;
wire n_168;
wire CTS_n_tid0_142;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire uc_0;
wire uc_1;
wire n_95;
wire n_94;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire CTS_n_tid0_40;
wire CTS_n_tid0_39;
wire n_147;


INV_X1 i_14 (.ZN (n_147), .A (n_168));
DFF_X1 \Input1_1_Positive_reg[63]  (.Q (\Input1_1_Positive[63] ), .CK (CTS_n_tid1_42), .D (in1[31]));
DFF_X1 \Input1_2_Positive_reg[1]  (.Q (\Input1_2_Positive[1] ), .CK (CTS_n_tid1_41), .D (in1[0]));
DFF_X1 \Input1_2_Positive_reg[31]  (.Q (\Input1_2_Positive[31] ), .CK (CTS_n_tid1_42), .D (in1[30]));
DFF_X1 \Input1_2_Negative_reg[31]  (.Q (\Input1_2_Negative[31] ), .CK (CTS_n_tid1_42), .D (n_62));
DFF_X1 \Input1_1_Positive_reg[29]  (.Q (\Input1_1_Positive[29] ), .CK (CTS_n_tid1_42), .D (in1[29]));
DFF_X1 \Input1_1_Negative_reg[29]  (.Q (\Input1_1_Negative[29] ), .CK (CTS_n_tid1_42), .D (n_61));
DFF_X1 \Input1_2_Positive_reg[15]  (.Q (\Input1_2_Positive[15] ), .CK (CTS_n_tid1_42), .D (in1[14]));
DFF_X1 \Input1_2_Negative_reg[15]  (.Q (\Input1_2_Negative[15] ), .CK (CTS_n_tid1_42), .D (n_46));
DFF_X1 \Input1_1_Positive_reg[13]  (.Q (\Input1_1_Positive[13] ), .CK (CTS_n_tid1_42), .D (in1[13]));
DFF_X1 \Input1_1_Negative_reg[13]  (.Q (\Input1_1_Negative[13] ), .CK (CTS_n_tid1_42), .D (n_45));
DFF_X1 \Input1_2_Positive_reg[23]  (.Q (\Input1_2_Positive[23] ), .CK (CTS_n_tid1_42), .D (in1[22]));
DFF_X1 \Input1_2_Negative_reg[23]  (.Q (\Input1_2_Negative[23] ), .CK (CTS_n_tid1_42), .D (n_54));
DFF_X1 \Input1_1_Positive_reg[21]  (.Q (\Input1_1_Positive[21] ), .CK (CTS_n_tid1_42), .D (in1[21]));
DFF_X1 \Input1_1_Negative_reg[21]  (.Q (\Input1_1_Negative[21] ), .CK (CTS_n_tid1_42), .D (n_53));
DFF_X1 \Input1_2_Positive_reg[7]  (.Q (\Input1_2_Positive[7] ), .CK (CTS_n_tid1_41), .D (in1[6]));
DFF_X1 \Input1_2_Negative_reg[7]  (.Q (\Input1_2_Negative[7] ), .CK (CTS_n_tid1_41), .D (n_38));
DFF_X1 \Input1_1_Positive_reg[5]  (.Q (\Input1_1_Positive[5] ), .CK (CTS_n_tid1_41), .D (in1[5]));
DFF_X1 \Input1_1_Negative_reg[5]  (.Q (\Input1_1_Negative[5] ), .CK (CTS_n_tid1_41), .D (n_37));
DFF_X1 \Input1_2_Positive_reg[27]  (.Q (\Input1_2_Positive[27] ), .CK (CTS_n_tid1_42), .D (in1[26]));
DFF_X1 \Input1_2_Negative_reg[27]  (.Q (\Input1_2_Negative[27] ), .CK (CTS_n_tid1_42), .D (n_58));
DFF_X1 \Input1_1_Positive_reg[25]  (.Q (\Input1_1_Positive[25] ), .CK (CTS_n_tid1_42), .D (in1[25]));
DFF_X1 \Input1_1_Negative_reg[25]  (.Q (\Input1_1_Negative[25] ), .CK (CTS_n_tid1_42), .D (n_57));
DFF_X1 \Input1_2_Positive_reg[11]  (.Q (\Input1_2_Positive[11] ), .CK (CTS_n_tid1_42), .D (in1[10]));
DFF_X1 \Input1_2_Negative_reg[11]  (.Q (\Input1_2_Negative[11] ), .CK (CTS_n_tid1_42), .D (n_42));
DFF_X1 \Input1_1_Positive_reg[9]  (.Q (\Input1_1_Positive[9] ), .CK (CTS_n_tid1_42), .D (in1[9]));
DFF_X1 \Input1_1_Negative_reg[9]  (.Q (\Input1_1_Negative[9] ), .CK (CTS_n_tid1_42), .D (n_41));
DFF_X1 \Input1_2_Positive_reg[19]  (.Q (\Input1_2_Positive[19] ), .CK (CTS_n_tid1_42), .D (in1[18]));
DFF_X1 \Input1_2_Negative_reg[19]  (.Q (\Input1_2_Negative[19] ), .CK (CTS_n_tid1_42), .D (n_50));
DFF_X1 \Input1_1_Positive_reg[17]  (.Q (\Input1_1_Positive[17] ), .CK (CTS_n_tid1_42), .D (in1[17]));
DFF_X1 \Input1_1_Negative_reg[17]  (.Q (\Input1_1_Negative[17] ), .CK (CTS_n_tid1_42), .D (n_49));
DFF_X1 \Input1_2_Positive_reg[3]  (.Q (\Input1_2_Positive[3] ), .CK (CTS_n_tid1_41), .D (in1[2]));
DFF_X1 \Input1_2_Negative_reg[3]  (.Q (\Input1_2_Negative[3] ), .CK (CTS_n_tid1_41), .D (n_34));
DFF_X1 \Input1_1_Positive_reg[1]  (.Q (\Input1_1_Positive[1] ), .CK (CTS_n_tid1_41), .D (in1[1]));
DFF_X1 \Input1_1_Negative_reg[1]  (.Q (\Input1_1_Negative[1] ), .CK (CTS_n_tid1_41), .D (n_33));
DFF_X1 \Input1_2_Positive_reg[29]  (.Q (\Input1_2_Positive[29] ), .CK (CTS_n_tid1_42), .D (in1[28]));
DFF_X1 \Input1_2_Negative_reg[29]  (.Q (\Input1_2_Negative[29] ), .CK (CTS_n_tid1_42), .D (n_60));
DFF_X1 \Input1_1_Positive_reg[27]  (.Q (\Input1_1_Positive[27] ), .CK (CTS_n_tid1_42), .D (in1[27]));
DFF_X1 \Input1_1_Negative_reg[27]  (.Q (\Input1_1_Negative[27] ), .CK (CTS_n_tid1_42), .D (n_59));
DFF_X1 \Input1_2_Positive_reg[13]  (.Q (\Input1_2_Positive[13] ), .CK (CTS_n_tid1_42), .D (in1[12]));
DFF_X1 \Input1_2_Negative_reg[13]  (.Q (\Input1_2_Negative[13] ), .CK (CTS_n_tid1_42), .D (n_44));
DFF_X1 \Input1_1_Positive_reg[11]  (.Q (\Input1_1_Positive[11] ), .CK (CTS_n_tid1_42), .D (in1[11]));
DFF_X1 \Input1_1_Negative_reg[11]  (.Q (\Input1_1_Negative[11] ), .CK (CTS_n_tid1_42), .D (n_43));
DFF_X1 \Input1_2_Positive_reg[21]  (.Q (\Input1_2_Positive[21] ), .CK (CTS_n_tid1_42), .D (in1[20]));
DFF_X1 \Input1_2_Negative_reg[21]  (.Q (\Input1_2_Negative[21] ), .CK (CTS_n_tid1_42), .D (n_52));
DFF_X1 \Input1_1_Positive_reg[19]  (.Q (\Input1_1_Positive[19] ), .CK (CTS_n_tid1_42), .D (in1[19]));
DFF_X1 \Input1_1_Negative_reg[19]  (.Q (\Input1_1_Negative[19] ), .CK (CTS_n_tid1_42), .D (n_51));
DFF_X1 \Input1_2_Positive_reg[5]  (.Q (\Input1_2_Positive[5] ), .CK (CTS_n_tid1_41), .D (in1[4]));
DFF_X1 \Input1_2_Negative_reg[5]  (.Q (\Input1_2_Negative[5] ), .CK (CTS_n_tid1_41), .D (n_36));
DFF_X1 \Input1_1_Positive_reg[3]  (.Q (\Input1_1_Positive[3] ), .CK (CTS_n_tid1_41), .D (in1[3]));
DFF_X1 \Input1_1_Negative_reg[3]  (.Q (\Input1_1_Negative[3] ), .CK (CTS_n_tid1_41), .D (n_35));
DFF_X1 \Input1_2_Positive_reg[25]  (.Q (\Input1_2_Positive[25] ), .CK (CTS_n_tid1_42), .D (in1[24]));
DFF_X1 \Input1_2_Negative_reg[25]  (.Q (\Input1_2_Negative[25] ), .CK (CTS_n_tid1_42), .D (n_56));
DFF_X1 \Input1_1_Positive_reg[23]  (.Q (\Input1_1_Positive[23] ), .CK (CTS_n_tid1_42), .D (in1[23]));
DFF_X1 \Input1_1_Negative_reg[23]  (.Q (\Input1_1_Negative[23] ), .CK (CTS_n_tid1_42), .D (n_55));
DFF_X1 \Input1_2_Positive_reg[9]  (.Q (\Input1_2_Positive[9] ), .CK (CTS_n_tid1_42), .D (in1[8]));
DFF_X1 \Input1_2_Negative_reg[9]  (.Q (\Input1_2_Negative[9] ), .CK (CTS_n_tid1_42), .D (n_40));
DFF_X1 \Input1_1_Positive_reg[7]  (.Q (\Input1_1_Positive[7] ), .CK (CTS_n_tid1_42), .D (in1[7]));
DFF_X1 \Input1_1_Negative_reg[7]  (.Q (\Input1_1_Negative[7] ), .CK (CTS_n_tid1_42), .D (n_39));
DFF_X1 \Input1_2_Positive_reg[17]  (.Q (\Input1_2_Positive[17] ), .CK (CTS_n_tid1_42), .D (in1[16]));
DFF_X1 \Input1_2_Negative_reg[17]  (.Q (\Input1_2_Negative[17] ), .CK (CTS_n_tid1_42), .D (n_48));
DFF_X1 \Input1_1_Positive_reg[15]  (.Q (\Input1_1_Positive[15] ), .CK (CTS_n_tid1_42), .D (in1[15]));
DFF_X1 \Input1_1_Negative_reg[15]  (.Q (\Input1_1_Negative[15] ), .CK (CTS_n_tid1_42), .D (n_47));
DFF_X1 \Input1_1_Negative_reg[63]  (.Q (\Input1_1_Negative[63] ), .CK (CTS_n_tid1_42), .D (n_63));
CLKGATETST_X8 clk_gate_Input1_1_Positive_reg (.GCK (CTS_n_tid1_133), .CK (clk_CTS_1_PP_2)
    , .E (start), .SE (1'b0 ));
CLKGATETST_X8 clk_gate_tempResult_reg (.GCK (CTS_n_tid0_105), .CK (n_tid1_233), .E (n_147), .SE (1'b0 ));
DFF_X1 \newB_reg[1]  (.Q (\newB[1] ), .CK (CTS_n_tid1_41), .D (in2[0]));
DFF_X1 \newB_reg[2]  (.Q (\newB[2] ), .CK (CTS_n_tid1_41), .D (in2[1]));
DFF_X1 \newB_reg[3]  (.Q (\newB[3] ), .CK (CTS_n_tid1_41), .D (in2[2]));
DFF_X1 \newB_reg[4]  (.Q (\newB[4] ), .CK (CTS_n_tid1_41), .D (in2[3]));
DFF_X1 \newB_reg[5]  (.Q (\newB[5] ), .CK (CTS_n_tid1_41), .D (in2[4]));
DFF_X1 \newB_reg[6]  (.Q (\newB[6] ), .CK (CTS_n_tid1_41), .D (in2[5]));
DFF_X1 \newB_reg[7]  (.Q (\newB[7] ), .CK (CTS_n_tid1_41), .D (in2[6]));
DFF_X1 \newB_reg[8]  (.Q (\newB[8] ), .CK (CTS_n_tid1_41), .D (in2[7]));
DFF_X1 \newB_reg[9]  (.Q (\newB[9] ), .CK (CTS_n_tid1_41), .D (in2[8]));
DFF_X1 \newB_reg[10]  (.Q (\newB[10] ), .CK (CTS_n_tid1_41), .D (in2[9]));
DFF_X1 \newB_reg[11]  (.Q (\newB[11] ), .CK (CTS_n_tid1_41), .D (in2[10]));
DFF_X1 \newB_reg[12]  (.Q (\newB[12] ), .CK (CTS_n_tid1_41), .D (in2[11]));
DFF_X1 \newB_reg[13]  (.Q (\newB[13] ), .CK (CTS_n_tid1_41), .D (in2[12]));
DFF_X1 \newB_reg[14]  (.Q (\newB[14] ), .CK (CTS_n_tid1_41), .D (in2[13]));
DFF_X1 \newB_reg[15]  (.Q (\newB[15] ), .CK (CTS_n_tid1_41), .D (in2[14]));
DFF_X1 \newB_reg[16]  (.Q (\newB[16] ), .CK (CTS_n_tid1_41), .D (in2[15]));
DFF_X1 \newB_reg[17]  (.Q (\newB[17] ), .CK (CTS_n_tid1_41), .D (in2[16]));
DFF_X1 \newB_reg[18]  (.Q (\newB[18] ), .CK (CTS_n_tid1_41), .D (in2[17]));
DFF_X1 \newB_reg[19]  (.Q (\newB[19] ), .CK (CTS_n_tid1_41), .D (in2[18]));
DFF_X1 \newB_reg[20]  (.Q (\newB[20] ), .CK (CTS_n_tid1_41), .D (in2[19]));
DFF_X1 \newB_reg[21]  (.Q (\newB[21] ), .CK (CTS_n_tid1_41), .D (in2[20]));
DFF_X1 \newB_reg[22]  (.Q (\newB[22] ), .CK (CTS_n_tid1_41), .D (in2[21]));
DFF_X1 \newB_reg[23]  (.Q (\newB[23] ), .CK (CTS_n_tid1_41), .D (in2[22]));
DFF_X1 \newB_reg[24]  (.Q (\newB[24] ), .CK (CTS_n_tid1_41), .D (in2[23]));
DFF_X1 \newB_reg[25]  (.Q (\newB[25] ), .CK (CTS_n_tid1_41), .D (in2[24]));
DFF_X1 \newB_reg[26]  (.Q (\newB[26] ), .CK (CTS_n_tid1_41), .D (in2[25]));
DFF_X1 \newB_reg[27]  (.Q (\newB[27] ), .CK (CTS_n_tid1_41), .D (in2[26]));
DFF_X1 \newB_reg[28]  (.Q (\newB[28] ), .CK (CTS_n_tid1_41), .D (in2[27]));
DFF_X1 \newB_reg[29]  (.Q (\newB[29] ), .CK (CTS_n_tid1_41), .D (in2[28]));
DFF_X1 \newB_reg[30]  (.Q (\newB[30] ), .CK (CTS_n_tid1_41), .D (in2[29]));
DFF_X1 \newB_reg[31]  (.Q (\newB[31] ), .CK (CTS_n_tid1_41), .D (in2[30]));
DFF_X1 \newB_reg[34]  (.Q (\newB[34] ), .CK (CTS_n_tid1_41), .D (in2[31]));
DFF_X1 \shiftingAmount_reg[1]  (.Q (\shiftingAmount[1] ), .CK (CTS_n_tid0_39), .D (n_163));
DFF_X1 \shiftingAmount_reg[2]  (.Q (\shiftingAmount[2] ), .CK (CTS_n_tid0_39), .D (n_164));
DFF_X1 \shiftingAmount_reg[3]  (.Q (\shiftingAmount[3] ), .CK (CTS_n_tid0_40), .D (n_165));
DFF_X1 \shiftingAmount_reg[4]  (.Q (\shiftingAmount[4] ), .CK (CTS_n_tid0_39), .D (n_166));
DFF_X1 \shiftingAmount_reg[5]  (.Q (\shiftingAmount[5] ), .CK (CTS_n_tid0_40), .D (n_167));
DFF_X1 \tempResult_reg[0]  (.Q (\tempResult[0] ), .CK (CTS_n_tid0_39), .D (n_96));
DFF_X1 \tempResult_reg[1]  (.Q (\tempResult[1] ), .CK (CTS_n_tid0_39), .D (n_97));
DFF_X1 \tempResult_reg[2]  (.Q (\tempResult[2] ), .CK (CTS_n_tid0_39), .D (n_98));
DFF_X1 \tempResult_reg[3]  (.Q (\tempResult[3] ), .CK (CTS_n_tid0_39), .D (n_99));
DFF_X1 \tempResult_reg[4]  (.Q (\tempResult[4] ), .CK (CTS_n_tid0_39), .D (n_100));
DFF_X1 \tempResult_reg[5]  (.Q (\tempResult[5] ), .CK (CTS_n_tid0_39), .D (n_101));
DFF_X1 \tempResult_reg[6]  (.Q (\tempResult[6] ), .CK (CTS_n_tid0_39), .D (n_102));
DFF_X1 \tempResult_reg[7]  (.Q (\tempResult[7] ), .CK (CTS_n_tid0_39), .D (n_103));
DFF_X1 \tempResult_reg[8]  (.Q (\tempResult[8] ), .CK (CTS_n_tid0_39), .D (n_104));
DFF_X1 \tempResult_reg[9]  (.Q (\tempResult[9] ), .CK (CTS_n_tid0_39), .D (n_105));
DFF_X1 \tempResult_reg[10]  (.Q (\tempResult[10] ), .CK (CTS_n_tid0_39), .D (n_106));
DFF_X1 \tempResult_reg[11]  (.Q (\tempResult[11] ), .CK (CTS_n_tid0_39), .D (n_107));
DFF_X1 \tempResult_reg[12]  (.Q (\tempResult[12] ), .CK (CTS_n_tid0_39), .D (n_108));
DFF_X1 \tempResult_reg[13]  (.Q (\tempResult[13] ), .CK (CTS_n_tid0_39), .D (n_109));
DFF_X1 \tempResult_reg[14]  (.Q (\tempResult[14] ), .CK (CTS_n_tid0_39), .D (n_110));
DFF_X1 \tempResult_reg[15]  (.Q (\tempResult[15] ), .CK (CTS_n_tid0_39), .D (n_111));
DFF_X1 \tempResult_reg[16]  (.Q (\tempResult[16] ), .CK (CTS_n_tid0_39), .D (n_112));
DFF_X1 \tempResult_reg[17]  (.Q (\tempResult[17] ), .CK (CTS_n_tid0_39), .D (n_113));
DFF_X1 \tempResult_reg[18]  (.Q (\tempResult[18] ), .CK (CTS_n_tid0_39), .D (n_114));
DFF_X1 \tempResult_reg[19]  (.Q (\tempResult[19] ), .CK (CTS_n_tid0_39), .D (n_115));
DFF_X1 \tempResult_reg[20]  (.Q (\tempResult[20] ), .CK (CTS_n_tid0_40), .D (n_116));
DFF_X1 \tempResult_reg[21]  (.Q (\tempResult[21] ), .CK (CTS_n_tid0_40), .D (n_117));
DFF_X1 \tempResult_reg[22]  (.Q (\tempResult[22] ), .CK (CTS_n_tid0_40), .D (n_118));
DFF_X1 \tempResult_reg[23]  (.Q (\tempResult[23] ), .CK (CTS_n_tid0_40), .D (n_119));
DFF_X1 \tempResult_reg[24]  (.Q (\tempResult[24] ), .CK (CTS_n_tid0_40), .D (n_120));
DFF_X1 \tempResult_reg[25]  (.Q (\tempResult[25] ), .CK (CTS_n_tid0_40), .D (n_121));
DFF_X1 \tempResult_reg[26]  (.Q (\tempResult[26] ), .CK (CTS_n_tid0_40), .D (n_122));
DFF_X1 \tempResult_reg[27]  (.Q (\tempResult[27] ), .CK (CTS_n_tid0_40), .D (n_123));
DFF_X1 \tempResult_reg[28]  (.Q (\tempResult[28] ), .CK (CTS_n_tid0_40), .D (n_124));
DFF_X1 \tempResult_reg[29]  (.Q (\tempResult[29] ), .CK (CTS_n_tid0_40), .D (n_125));
DFF_X1 \tempResult_reg[30]  (.Q (\tempResult[30] ), .CK (CTS_n_tid0_40), .D (n_126));
DFF_X1 \tempResult_reg[31]  (.Q (\tempResult[31] ), .CK (CTS_n_tid0_40), .D (n_127));
DFF_X1 \tempResult_reg[32]  (.Q (\tempResult[32] ), .CK (CTS_n_tid0_40), .D (n_128));
DFF_X1 \tempResult_reg[33]  (.Q (\tempResult[33] ), .CK (CTS_n_tid0_40), .D (n_129));
DFF_X1 \tempResult_reg[34]  (.Q (\tempResult[34] ), .CK (CTS_n_tid0_39), .D (n_130));
DFF_X1 \tempResult_reg[35]  (.Q (\tempResult[35] ), .CK (CTS_n_tid0_39), .D (n_131));
DFF_X1 \tempResult_reg[36]  (.Q (\tempResult[36] ), .CK (CTS_n_tid0_39), .D (n_132));
DFF_X1 \tempResult_reg[37]  (.Q (\tempResult[37] ), .CK (CTS_n_tid0_39), .D (n_133));
DFF_X1 \tempResult_reg[38]  (.Q (\tempResult[38] ), .CK (CTS_n_tid0_39), .D (n_134));
DFF_X1 \tempResult_reg[39]  (.Q (\tempResult[39] ), .CK (CTS_n_tid0_39), .D (n_135));
DFF_X1 \tempResult_reg[40]  (.Q (\tempResult[40] ), .CK (CTS_n_tid0_39), .D (n_136));
DFF_X1 \tempResult_reg[41]  (.Q (\tempResult[41] ), .CK (CTS_n_tid0_39), .D (n_137));
DFF_X1 \tempResult_reg[42]  (.Q (\tempResult[42] ), .CK (CTS_n_tid0_39), .D (n_138));
DFF_X1 \tempResult_reg[43]  (.Q (\tempResult[43] ), .CK (CTS_n_tid0_39), .D (n_139));
DFF_X1 \tempResult_reg[44]  (.Q (\tempResult[44] ), .CK (CTS_n_tid0_39), .D (n_140));
DFF_X1 \tempResult_reg[45]  (.Q (\tempResult[45] ), .CK (CTS_n_tid0_39), .D (n_141));
DFF_X1 \tempResult_reg[46]  (.Q (\tempResult[46] ), .CK (CTS_n_tid0_39), .D (n_142));
DFF_X1 \tempResult_reg[47]  (.Q (\tempResult[47] ), .CK (CTS_n_tid0_39), .D (n_143));
DFF_X1 \tempResult_reg[48]  (.Q (\tempResult[48] ), .CK (CTS_n_tid0_40), .D (n_144));
DFF_X1 \tempResult_reg[49]  (.Q (\tempResult[49] ), .CK (CTS_n_tid0_40), .D (n_148));
DFF_X1 \tempResult_reg[50]  (.Q (\tempResult[50] ), .CK (CTS_n_tid0_40), .D (n_149));
DFF_X1 \tempResult_reg[51]  (.Q (\tempResult[51] ), .CK (CTS_n_tid0_40), .D (n_150));
DFF_X1 \tempResult_reg[52]  (.Q (\tempResult[52] ), .CK (CTS_n_tid0_40), .D (n_151));
DFF_X1 \tempResult_reg[53]  (.Q (\tempResult[53] ), .CK (CTS_n_tid0_40), .D (n_152));
DFF_X1 \tempResult_reg[54]  (.Q (\tempResult[54] ), .CK (CTS_n_tid0_40), .D (n_153));
DFF_X1 \tempResult_reg[55]  (.Q (\tempResult[55] ), .CK (CTS_n_tid0_40), .D (n_154));
DFF_X1 \tempResult_reg[56]  (.Q (\tempResult[56] ), .CK (CTS_n_tid0_40), .D (n_155));
DFF_X1 \tempResult_reg[57]  (.Q (\tempResult[57] ), .CK (CTS_n_tid0_40), .D (n_156));
DFF_X1 \tempResult_reg[58]  (.Q (\tempResult[58] ), .CK (CTS_n_tid0_40), .D (n_157));
DFF_X1 \tempResult_reg[59]  (.Q (\tempResult[59] ), .CK (CTS_n_tid0_40), .D (n_158));
DFF_X1 \tempResult_reg[60]  (.Q (\tempResult[60] ), .CK (CTS_n_tid0_40), .D (n_159));
DFF_X1 \tempResult_reg[61]  (.Q (\tempResult[61] ), .CK (CTS_n_tid0_40), .D (n_160));
DFF_X1 \tempResult_reg[62]  (.Q (\tempResult[62] ), .CK (CTS_n_tid0_40), .D (n_161));
DFF_X1 \tempResult_reg[63]  (.Q (\tempResult[63] ), .CK (CTS_n_tid0_40), .D (n_162));
OAI21_X1 i_0_502 (.ZN (n_0_380), .A (n_0_331__1), .B1 (n_0_8), .B2 (n_0_371__1));
INV_X1 i_0_501 (.ZN (n_0_371__1), .A (n_0_253));
AOI21_X1 i_0_500 (.ZN (n_0_379), .A (n_0_370__1), .B1 (n_0_368__1), .B2 (hfn_ipo_n32));
AOI21_X1 i_0_499 (.ZN (n_0_378), .A (n_0_370__1), .B1 (n_0_365__1), .B2 (hfn_ipo_n32));
NOR2_X1 i_0_498 (.ZN (n_0_370__1), .A1 (n_0_381), .A2 (hfn_ipo_n32));
OAI21_X1 i_0_497 (.ZN (n_0_381), .A (n_0_331__1), .B1 (n_0_8), .B2 (n_0_369__1));
INV_X1 i_0_496 (.ZN (n_0_369__1), .A (n_0_259));
OAI22_X1 i_0_495 (.ZN (n_0_377), .A1 (n_0_362__1), .A2 (hfn_ipo_n28), .B1 (n_0_368__1), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_494 (.ZN (n_0_368__1), .A1 (n_0_355__1), .A2 (hfn_ipo_n30), .B1 (n_0_367__1), .B2 (hfn_ipo_n26));
OAI21_X1 i_0_493 (.ZN (n_0_367__1), .A (n_0_331__1), .B1 (n_0_8), .B2 (n_0_366__1));
INV_X1 i_0_492 (.ZN (n_0_366__1), .A (n_0_247));
OAI22_X1 i_0_491 (.ZN (n_0_376), .A1 (n_0_359__1), .A2 (hfn_ipo_n28), .B1 (n_0_365__1), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_490 (.ZN (n_0_365__1), .A1 (n_0_352__1), .A2 (hfn_ipo_n30), .B1 (n_0_364__1), .B2 (hfn_ipo_n26));
OAI21_X1 i_0_489 (.ZN (n_0_364__1), .A (n_0_331__1), .B1 (n_0_8), .B2 (n_0_363__1));
INV_X1 i_0_488 (.ZN (n_0_363__1), .A (n_0_241));
OAI22_X1 i_0_487 (.ZN (n_0_375), .A1 (n_0_356__1), .A2 (hfn_ipo_n28), .B1 (n_0_362__1), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_486 (.ZN (n_0_362__1), .A1 (n_0_349__1), .A2 (hfn_ipo_n30), .B1 (hfn_ipo_n26), .B2 (n_0_361__1));
OAI21_X1 i_0_485 (.ZN (n_0_361__1), .A (n_0_331__1), .B1 (n_0_8), .B2 (n_0_360__1));
INV_X1 i_0_484 (.ZN (n_0_360__1), .A (n_0_235));
OAI22_X1 i_0_483 (.ZN (n_0_374), .A1 (n_0_353__1), .A2 (hfn_ipo_n28), .B1 (n_0_359__1), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_482 (.ZN (n_0_359__1), .A1 (n_0_346__1), .A2 (hfn_ipo_n30), .B1 (hfn_ipo_n26), .B2 (n_0_358__1));
OAI21_X1 i_0_481 (.ZN (n_0_358__1), .A (n_0_331__1), .B1 (n_0_8), .B2 (n_0_357__1));
INV_X1 i_0_480 (.ZN (n_0_357__1), .A (n_0_229));
OAI22_X1 i_0_479 (.ZN (n_0_373), .A1 (n_0_350__1), .A2 (hfn_ipo_n28), .B1 (n_0_356__1), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_478 (.ZN (n_0_356__1), .A1 (n_0_355__1), .A2 (hfn_ipo_n26), .B1 (n_0_343__1), .B2 (hfn_ipo_n30));
AOI21_X1 i_0_477 (.ZN (n_0_355__1), .A (n_0_354__1), .B1 (n_0_328__1), .B2 (drc_ipo_n33));
AOI21_X1 i_0_476 (.ZN (n_0_354__1), .A (n_0_332__1), .B1 (drc_ipo_n34), .B2 (n_0_223));
OAI22_X1 i_0_475 (.ZN (n_0_372), .A1 (n_0_347__1), .A2 (hfn_ipo_n28), .B1 (n_0_353__1), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_474 (.ZN (n_0_353__1), .A1 (n_0_340__1), .A2 (hfn_ipo_n30), .B1 (n_0_352__1), .B2 (hfn_ipo_n26));
AOI21_X1 i_0_473 (.ZN (n_0_352__1), .A (n_0_351__1), .B1 (n_0_325__1), .B2 (drc_ipo_n33));
AOI21_X1 i_0_472 (.ZN (n_0_351__1), .A (n_0_332__1), .B1 (drc_ipo_n34), .B2 (n_0_217));
OAI22_X1 i_0_471 (.ZN (n_0_371__0), .A1 (n_0_350__1), .A2 (hfn_ipo_n32), .B1 (n_0_344__1), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_470 (.ZN (n_0_350__1), .A1 (n_0_337__1), .A2 (hfn_ipo_n30), .B1 (n_0_349__1), .B2 (hfn_ipo_n26));
AOI21_X1 i_0_469 (.ZN (n_0_349__1), .A (n_0_348__1), .B1 (n_0_322__1), .B2 (drc_ipo_n33));
AOI21_X1 i_0_468 (.ZN (n_0_348__1), .A (n_0_332__1), .B1 (drc_ipo_n34), .B2 (n_0_211));
OAI22_X1 i_0_467 (.ZN (n_0_370__0), .A1 (n_0_347__1), .A2 (hfn_ipo_n32), .B1 (n_0_341__1), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_466 (.ZN (n_0_347__1), .A1 (n_0_334__1), .A2 (hfn_ipo_n30), .B1 (n_0_346__1), .B2 (hfn_ipo_n26));
AOI21_X1 i_0_465 (.ZN (n_0_346__1), .A (n_0_345__1), .B1 (n_0_319), .B2 (drc_ipo_n33));
AOI21_X1 i_0_464 (.ZN (n_0_345__1), .A (n_0_332__1), .B1 (drc_ipo_n34), .B2 (n_0_205));
OAI22_X1 i_0_463 (.ZN (n_0_369__0), .A1 (n_0_338__1), .A2 (hfn_ipo_n28), .B1 (n_0_344__1), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_462 (.ZN (n_0_344__1), .A1 (n_0_329__1), .A2 (hfn_ipo_n30), .B1 (n_0_343__1), .B2 (hfn_ipo_n26));
AOI21_X1 i_0_461 (.ZN (n_0_343__1), .A (n_0_342__1), .B1 (n_0_316__1), .B2 (drc_ipo_n33));
AOI21_X1 i_0_460 (.ZN (n_0_342__1), .A (n_0_332__1), .B1 (drc_ipo_n34), .B2 (n_0_199));
OAI22_X1 i_0_459 (.ZN (n_0_368__0), .A1 (n_0_335__1), .A2 (hfn_ipo_n28), .B1 (n_0_341__1), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_458 (.ZN (n_0_341__1), .A1 (n_0_326__1), .A2 (hfn_ipo_n30), .B1 (n_0_340__1), .B2 (hfn_ipo_n26));
AOI21_X1 i_0_457 (.ZN (n_0_340__1), .A (n_0_339__1), .B1 (n_0_313), .B2 (drc_ipo_n33));
AOI21_X1 i_0_456 (.ZN (n_0_339__1), .A (n_0_332__1), .B1 (drc_ipo_n34), .B2 (n_0_193));
OAI22_X1 i_0_455 (.ZN (n_0_367__0), .A1 (n_0_338__1), .A2 (hfn_ipo_n32), .B1 (n_0_330__1), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_454 (.ZN (n_0_338__1), .A1 (n_0_323__1), .A2 (hfn_ipo_n30), .B1 (n_0_337__1), .B2 (hfn_ipo_n26));
AOI21_X1 i_0_453 (.ZN (n_0_337__1), .A (n_0_336__1), .B1 (n_0_310), .B2 (drc_ipo_n33));
AOI21_X1 i_0_452 (.ZN (n_0_336__1), .A (n_0_332__1), .B1 (drc_ipo_n34), .B2 (n_0_187));
OAI22_X1 i_0_451 (.ZN (n_0_366__0), .A1 (n_0_335__1), .A2 (hfn_ipo_n32), .B1 (n_0_327__1), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_450 (.ZN (n_0_335__1), .A1 (n_0_320__1), .A2 (hfn_ipo_n30), .B1 (n_0_334__1), .B2 (hfn_ipo_n26));
AOI21_X1 i_0_449 (.ZN (n_0_334__1), .A (n_0_333__1), .B1 (n_0_307), .B2 (drc_ipo_n33));
AOI21_X1 i_0_448 (.ZN (n_0_333__1), .A (n_0_332__1), .B1 (drc_ipo_n34), .B2 (n_0_181));
NAND2_X1 i_0_447 (.ZN (n_0_332__1), .A1 (n_0_331__1), .A2 (n_0_17));
NAND2_X1 i_0_446 (.ZN (n_0_331__1), .A1 (n_0_276), .A2 (n_0_8));
OAI22_X1 i_0_445 (.ZN (n_0_365__0), .A1 (n_0_324__1), .A2 (hfn_ipo_n27), .B1 (n_0_330__1), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_444 (.ZN (n_0_330__1), .A1 (n_0_317), .A2 (hfn_ipo_n30), .B1 (n_0_329__1), .B2 (hfn_ipo_n26));
OAI22_X1 i_0_443 (.ZN (n_0_329__1), .A1 (n_0_328__1), .A2 (drc_ipo_n33), .B1 (n_0_304), .B2 (n_0_17));
AOI221_X1 i_0_442 (.ZN (n_0_328__1), .A (n_0_278), .B1 (drc_ipo_n34), .B2 (n_0_175)
    , .C1 (n_0_16), .C2 (n_0_271));
OAI22_X1 i_0_441 (.ZN (n_0_364__0), .A1 (n_0_321__1), .A2 (hfn_ipo_n28), .B1 (n_0_327__1), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_440 (.ZN (n_0_327__1), .A1 (n_0_314), .A2 (hfn_ipo_n30), .B1 (n_0_326__1), .B2 (hfn_ipo_n26));
OAI22_X1 i_0_439 (.ZN (n_0_326__1), .A1 (n_0_325__1), .A2 (drc_ipo_n33), .B1 (n_0_300), .B2 (n_0_17));
AOI221_X1 i_0_438 (.ZN (n_0_325__1), .A (n_0_278), .B1 (n_0_16), .B2 (n_0_265), .C1 (drc_ipo_n34), .C2 (n_0_168));
OAI22_X1 i_0_437 (.ZN (n_0_363__0), .A1 (n_0_324__1), .A2 (hfn_ipo_n31), .B1 (hfn_ipo_n27), .B2 (n_0_318__1));
AOI22_X1 i_0_436 (.ZN (n_0_324__1), .A1 (n_0_311), .A2 (hfn_ipo_n29), .B1 (n_0_323__1), .B2 (n_0_20));
AOI22_X1 i_0_435 (.ZN (n_0_323__1), .A1 (n_0_296), .A2 (drc_ipo_n33), .B1 (n_0_322__1), .B2 (n_0_17));
AOI221_X1 i_0_434 (.ZN (n_0_322__1), .A (n_0_278), .B1 (n_0_16), .B2 (n_0_259), .C1 (drc_ipo_n34), .C2 (n_0_161));
OAI22_X1 i_0_433 (.ZN (n_0_362__0), .A1 (n_0_321__1), .A2 (hfn_ipo_n31), .B1 (hfn_ipo_n27), .B2 (n_0_315));
AOI22_X1 i_0_432 (.ZN (n_0_321__1), .A1 (n_0_308), .A2 (hfn_ipo_n30), .B1 (n_0_320__1), .B2 (hfn_ipo_n26));
OAI22_X1 i_0_431 (.ZN (n_0_320__1), .A1 (n_0_293), .A2 (n_0_17), .B1 (n_0_319), .B2 (drc_ipo_n33));
AOI221_X1 i_0_430 (.ZN (n_0_319), .A (n_0_278), .B1 (drc_ipo_n34), .B2 (n_0_155), .C1 (n_0_16), .C2 (n_0_253));
OAI22_X1 i_0_429 (.ZN (n_0_361__0), .A1 (n_0_312), .A2 (hfn_ipo_n27), .B1 (n_0_318__1), .B2 (hfn_ipo_n31));
AOI22_X1 i_0_428 (.ZN (n_0_318__1), .A1 (n_0_317), .A2 (hfn_ipo_n26), .B1 (hfn_ipo_n30), .B2 (n_0_305));
OAI22_X1 i_0_427 (.ZN (n_0_317), .A1 (n_0_316__1), .A2 (drc_ipo_n33), .B1 (n_0_290), .B2 (n_0_17));
AOI221_X1 i_0_426 (.ZN (n_0_316__1), .A (n_0_278), .B1 (n_0_16), .B2 (n_0_247), .C1 (drc_ipo_n34), .C2 (n_0_148));
OAI22_X1 i_0_425 (.ZN (n_0_360__0), .A1 (n_0_309), .A2 (hfn_ipo_n27), .B1 (n_0_315), .B2 (hfn_ipo_n31));
AOI22_X1 i_0_424 (.ZN (n_0_315), .A1 (n_0_314), .A2 (hfn_ipo_n26), .B1 (hfn_ipo_n30), .B2 (n_0_301));
OAI22_X1 i_0_423 (.ZN (n_0_314), .A1 (n_0_313), .A2 (drc_ipo_n33), .B1 (n_0_286), .B2 (n_0_17));
AOI221_X1 i_0_422 (.ZN (n_0_313), .A (n_0_278), .B1 (n_0_16), .B2 (n_0_241), .C1 (drc_ipo_n34), .C2 (n_0_142));
OAI22_X1 i_0_421 (.ZN (n_0_359__0), .A1 (n_0_312), .A2 (hfn_ipo_n31), .B1 (hfn_ipo_n27), .B2 (n_0_306));
AOI22_X1 i_0_420 (.ZN (n_0_312), .A1 (n_0_311), .A2 (n_0_20), .B1 (n_0_297), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_419 (.ZN (n_0_311), .A1 (n_0_282), .A2 (drc_ipo_n33), .B1 (n_0_310), .B2 (n_0_17));
AOI221_X1 i_0_418 (.ZN (n_0_310), .A (n_0_278), .B1 (drc_ipo_n34), .B2 (n_0_136), .C1 (n_0_16), .C2 (n_0_235));
OAI22_X1 i_0_417 (.ZN (n_0_358__0), .A1 (n_0_309), .A2 (hfn_ipo_n31), .B1 (hfn_ipo_n27), .B2 (n_0_302));
AOI22_X1 i_0_416 (.ZN (n_0_309), .A1 (n_0_308), .A2 (n_0_20), .B1 (n_0_294), .B2 (hfn_ipo_n29));
AOI22_X1 i_0_415 (.ZN (n_0_308), .A1 (n_0_279), .A2 (drc_ipo_n33), .B1 (n_0_307), .B2 (n_0_17));
AOI221_X1 i_0_414 (.ZN (n_0_307), .A (n_0_278), .B1 (drc_ipo_n34), .B2 (n_0_129), .C1 (n_0_16), .C2 (n_0_229));
OAI22_X1 i_0_413 (.ZN (n_0_357__0), .A1 (n_0_298), .A2 (hfn_ipo_n27), .B1 (n_0_306), .B2 (hfn_ipo_n31));
AOI22_X1 i_0_412 (.ZN (n_0_306), .A1 (n_0_291), .A2 (hfn_ipo_n29), .B1 (n_0_305), .B2 (n_0_20));
OAI22_X1 i_0_411 (.ZN (n_0_305), .A1 (n_0_304), .A2 (drc_ipo_n33), .B1 (n_0_17), .B2 (n_0_272));
AOI21_X1 i_0_410 (.ZN (n_0_304), .A (n_0_303), .B1 (n_0_16), .B2 (n_0_223));
OAI21_X1 i_0_409 (.ZN (n_0_303), .A (n_0_277), .B1 (n_0_8), .B2 (n_0_172));
OAI22_X1 i_0_408 (.ZN (n_0_356__0), .A1 (n_0_295), .A2 (hfn_ipo_n27), .B1 (n_0_302), .B2 (hfn_ipo_n31));
AOI22_X1 i_0_407 (.ZN (n_0_302), .A1 (n_0_287), .A2 (hfn_ipo_n30), .B1 (n_0_301), .B2 (hfn_ipo_n26));
OAI22_X1 i_0_406 (.ZN (n_0_301), .A1 (n_0_300), .A2 (drc_ipo_n33), .B1 (n_0_17), .B2 (n_0_266));
AOI21_X1 i_0_405 (.ZN (n_0_300), .A (n_0_299), .B1 (n_0_16), .B2 (n_0_217));
OAI21_X1 i_0_404 (.ZN (n_0_299), .A (n_0_277), .B1 (n_0_8), .B2 (n_0_120));
OAI22_X1 i_0_403 (.ZN (n_0_355__0), .A1 (n_0_298), .A2 (hfn_ipo_n31), .B1 (hfn_ipo_n27), .B2 (n_0_292));
AOI22_X1 i_0_402 (.ZN (n_0_298), .A1 (n_0_283), .A2 (hfn_ipo_n29), .B1 (n_0_297), .B2 (n_0_20));
OAI22_X1 i_0_401 (.ZN (n_0_297), .A1 (n_0_296), .A2 (drc_ipo_n33), .B1 (n_0_17), .B2 (n_0_260));
AOI221_X1 i_0_400 (.ZN (n_0_296), .A (n_0_278), .B1 (n_0_16), .B2 (n_0_211), .C1 (drc_ipo_n34), .C2 (n_0_115));
OAI22_X1 i_0_399 (.ZN (n_0_354__0), .A1 (n_0_295), .A2 (hfn_ipo_n31), .B1 (hfn_ipo_n27), .B2 (n_0_288));
AOI22_X1 i_0_398 (.ZN (n_0_295), .A1 (n_0_280), .A2 (hfn_ipo_n29), .B1 (n_0_294), .B2 (n_0_20));
OAI22_X1 i_0_397 (.ZN (n_0_294), .A1 (n_0_293), .A2 (drc_ipo_n33), .B1 (n_0_17), .B2 (n_0_254));
AOI221_X1 i_0_396 (.ZN (n_0_293), .A (n_0_278), .B1 (n_0_16), .B2 (n_0_205), .C1 (drc_ipo_n34), .C2 (n_0_105));
OAI22_X1 i_0_395 (.ZN (n_0_353__0), .A1 (n_0_284), .A2 (hfn_ipo_n28), .B1 (hfn_ipo_n32), .B2 (n_0_292));
AOI22_X1 i_0_394 (.ZN (n_0_292), .A1 (n_0_291), .A2 (n_0_20), .B1 (hfn_ipo_n29), .B2 (n_0_273));
OAI22_X1 i_0_393 (.ZN (n_0_291), .A1 (n_0_290), .A2 (drc_ipo_n33), .B1 (n_0_17), .B2 (n_0_248));
AOI21_X1 i_0_392 (.ZN (n_0_290), .A (n_0_289), .B1 (n_0_16), .B2 (n_0_199));
OAI21_X1 i_0_391 (.ZN (n_0_289), .A (n_0_277), .B1 (n_0_8), .B2 (n_0_102));
OAI22_X1 i_0_390 (.ZN (n_0_352__0), .A1 (n_0_281), .A2 (hfn_ipo_n28), .B1 (n_0_288), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_389 (.ZN (n_0_288), .A1 (n_0_287), .A2 (hfn_ipo_n26), .B1 (hfn_ipo_n30), .B2 (n_0_267));
OAI22_X1 i_0_388 (.ZN (n_0_287), .A1 (n_0_286), .A2 (drc_ipo_n33), .B1 (n_0_17), .B2 (n_0_242));
AOI21_X1 i_0_387 (.ZN (n_0_286), .A (n_0_285), .B1 (n_0_16), .B2 (n_0_193));
OAI21_X1 i_0_386 (.ZN (n_0_285), .A (n_0_277), .B1 (n_0_8), .B2 (n_0_97));
OAI22_X1 i_0_385 (.ZN (n_0_351__0), .A1 (n_0_284), .A2 (hfn_ipo_n32), .B1 (hfn_ipo_n28), .B2 (n_0_274));
AOI22_X1 i_0_384 (.ZN (n_0_284), .A1 (n_0_283), .A2 (n_0_20), .B1 (hfn_ipo_n29), .B2 (n_0_261));
OAI22_X1 i_0_383 (.ZN (n_0_283), .A1 (n_0_282), .A2 (drc_ipo_n33), .B1 (n_0_17), .B2 (n_0_236));
AOI221_X1 i_0_382 (.ZN (n_0_282), .A (n_0_278), .B1 (n_0_16), .B2 (n_0_187), .C1 (n_0_112), .C2 (drc_ipo_n34));
OAI22_X1 i_0_381 (.ZN (n_0_350__0), .A1 (n_0_281), .A2 (hfn_ipo_n32), .B1 (hfn_ipo_n28), .B2 (n_0_268));
AOI22_X1 i_0_380 (.ZN (n_0_281), .A1 (n_0_280), .A2 (hfn_ipo_n26), .B1 (hfn_ipo_n30), .B2 (n_0_255));
OAI22_X1 i_0_379 (.ZN (n_0_280), .A1 (n_0_279), .A2 (drc_ipo_n33), .B1 (n_0_17), .B2 (n_0_230));
AOI221_X1 i_0_378 (.ZN (n_0_279), .A (n_0_278), .B1 (drc_ipo_n34), .B2 (n_0_108), .C1 (n_0_16), .C2 (n_0_181));
INV_X1 i_0_377 (.ZN (n_0_278), .A (n_0_277));
NAND2_X2 i_0_376 (.ZN (n_0_277), .A1 (n_0_276), .A2 (n_0_109));
NAND2_X1 i_0_375 (.ZN (n_0_276), .A1 (n_0_269), .A2 (n_0_275));
AOI22_X1 i_0_374 (.ZN (n_0_275), .A1 (n_0_92), .A2 (\Input1_1_Positive[63] ), .B1 (n_0_94), .B2 (\Input1_1_Negative[63] ));
OAI22_X1 i_0_373 (.ZN (n_0_349__0), .A1 (n_0_262), .A2 (hfn_ipo_n28), .B1 (n_0_274), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_372 (.ZN (n_0_274), .A1 (n_0_249), .A2 (hfn_ipo_n30), .B1 (n_0_273), .B2 (hfn_ipo_n26));
OAI22_X1 i_0_371 (.ZN (n_0_273), .A1 (n_0_272), .A2 (drc_ipo_n33), .B1 (n_0_224), .B2 (n_0_61));
AOI22_X1 i_0_370 (.ZN (n_0_272), .A1 (n_0_271), .A2 (n_0_109), .B1 (n_0_175), .B2 (n_0_16));
NAND2_X1 i_0_369 (.ZN (n_0_271), .A1 (n_0_269), .A2 (n_0_270));
AOI22_X1 i_0_368 (.ZN (n_0_270), .A1 (n_0_92), .A2 (\Input1_2_Positive[31] ), .B1 (n_0_94), .B2 (\Input1_2_Negative[31] ));
AOI22_X1 i_0_367 (.ZN (n_0_269), .A1 (n_0_89), .A2 (\Input1_1_Negative[63] ), .B1 (n_0_90), .B2 (\Input1_1_Positive[63] ));
OAI22_X1 i_0_366 (.ZN (n_0_348__0), .A1 (n_0_268), .A2 (hfn_ipo_n32), .B1 (n_0_256), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_365 (.ZN (n_0_268), .A1 (n_0_243), .A2 (hfn_ipo_n30), .B1 (n_0_267), .B2 (hfn_ipo_n26));
OAI22_X1 i_0_364 (.ZN (n_0_267), .A1 (n_0_266), .A2 (drc_ipo_n33), .B1 (n_0_218), .B2 (n_0_61));
AOI22_X1 i_0_363 (.ZN (n_0_266), .A1 (n_0_265), .A2 (n_0_109), .B1 (n_0_168), .B2 (n_0_16));
NAND2_X1 i_0_362 (.ZN (n_0_265), .A1 (n_0_263), .A2 (n_0_264));
AOI22_X1 i_0_361 (.ZN (n_0_264), .A1 (n_0_90), .A2 (\Input1_2_Positive[31] ), .B1 (\Input1_1_Positive[29] ), .B2 (n_0_92));
AOI22_X1 i_0_360 (.ZN (n_0_263), .A1 (n_0_89), .A2 (\Input1_2_Negative[31] ), .B1 (\Input1_1_Negative[29] ), .B2 (n_0_94));
OAI22_X1 i_0_359 (.ZN (n_0_347__0), .A1 (n_0_262), .A2 (hfn_ipo_n32), .B1 (n_0_250), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_358 (.ZN (n_0_262), .A1 (n_0_237), .A2 (hfn_ipo_n29), .B1 (n_0_261), .B2 (n_0_20));
OAI22_X1 i_0_357 (.ZN (n_0_261), .A1 (n_0_260), .A2 (drc_ipo_n33), .B1 (n_0_212), .B2 (n_0_17));
AOI22_X1 i_0_356 (.ZN (n_0_260), .A1 (n_0_161), .A2 (n_0_16), .B1 (n_0_259), .B2 (n_0_109));
NAND2_X1 i_0_355 (.ZN (n_0_259), .A1 (n_0_257), .A2 (n_0_258));
AOI22_X1 i_0_354 (.ZN (n_0_258), .A1 (n_0_89), .A2 (\Input1_1_Negative[29] ), .B1 (\Input1_2_Negative[29] ), .B2 (n_0_94));
AOI22_X1 i_0_353 (.ZN (n_0_257), .A1 (n_0_90), .A2 (\Input1_1_Positive[29] ), .B1 (\Input1_2_Positive[29] ), .B2 (n_0_92));
OAI22_X1 i_0_352 (.ZN (n_0_346__0), .A1 (n_0_256), .A2 (hfn_ipo_n32), .B1 (n_0_244), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_351 (.ZN (n_0_256), .A1 (n_0_255), .A2 (hfn_ipo_n26), .B1 (n_0_231), .B2 (hfn_ipo_n30));
OAI22_X1 i_0_350 (.ZN (n_0_255), .A1 (n_0_254), .A2 (drc_ipo_n33), .B1 (n_0_206), .B2 (n_0_17));
AOI22_X1 i_0_349 (.ZN (n_0_254), .A1 (n_0_253), .A2 (n_0_109), .B1 (n_0_155), .B2 (n_0_16));
NAND2_X1 i_0_348 (.ZN (n_0_253), .A1 (n_0_251), .A2 (n_0_252));
AOI22_X1 i_0_347 (.ZN (n_0_252), .A1 (n_0_89), .A2 (\Input1_2_Negative[29] ), .B1 (\Input1_1_Positive[27] ), .B2 (n_0_92));
AOI22_X1 i_0_346 (.ZN (n_0_251), .A1 (n_0_90), .A2 (\Input1_2_Positive[29] ), .B1 (n_0_94), .B2 (\Input1_1_Negative[27] ));
OAI22_X1 i_0_345 (.ZN (n_0_345__0), .A1 (n_0_238), .A2 (hfn_ipo_n28), .B1 (n_0_250), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_344 (.ZN (n_0_250), .A1 (n_0_249), .A2 (hfn_ipo_n26), .B1 (n_0_225), .B2 (hfn_ipo_n30));
OAI22_X1 i_0_343 (.ZN (n_0_249), .A1 (n_0_248), .A2 (drc_ipo_n33), .B1 (n_0_200), .B2 (n_0_61));
AOI22_X1 i_0_342 (.ZN (n_0_248), .A1 (n_0_148), .A2 (n_0_16), .B1 (n_0_247), .B2 (n_0_109));
NAND2_X1 i_0_341 (.ZN (n_0_247), .A1 (n_0_245), .A2 (n_0_246));
AOI22_X1 i_0_340 (.ZN (n_0_246), .A1 (n_0_90), .A2 (\Input1_1_Positive[27] ), .B1 (\Input1_2_Positive[27] ), .B2 (n_0_92));
AOI22_X1 i_0_339 (.ZN (n_0_245), .A1 (n_0_89), .A2 (\Input1_1_Negative[27] ), .B1 (\Input1_2_Negative[27] ), .B2 (n_0_94));
OAI22_X1 i_0_338 (.ZN (n_0_344__0), .A1 (n_0_244), .A2 (hfn_ipo_n32), .B1 (n_0_232), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_337 (.ZN (n_0_244), .A1 (n_0_243), .A2 (hfn_ipo_n26), .B1 (n_0_219), .B2 (hfn_ipo_n30));
OAI22_X1 i_0_336 (.ZN (n_0_243), .A1 (n_0_242), .A2 (drc_ipo_n33), .B1 (n_0_194), .B2 (n_0_61));
AOI22_X1 i_0_335 (.ZN (n_0_242), .A1 (n_0_142), .A2 (n_0_16), .B1 (n_0_241), .B2 (n_0_109));
NAND2_X1 i_0_334 (.ZN (n_0_241), .A1 (n_0_239), .A2 (n_0_240));
AOI22_X1 i_0_333 (.ZN (n_0_240), .A1 (n_0_90), .A2 (\Input1_2_Positive[27] ), .B1 (\Input1_1_Positive[25] ), .B2 (n_0_92));
AOI22_X1 i_0_332 (.ZN (n_0_239), .A1 (n_0_89), .A2 (\Input1_2_Negative[27] ), .B1 (\Input1_1_Negative[25] ), .B2 (n_0_94));
OAI22_X1 i_0_331 (.ZN (n_0_343__0), .A1 (n_0_238), .A2 (hfn_ipo_n32), .B1 (n_0_226), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_330 (.ZN (n_0_238), .A1 (n_0_237), .A2 (n_0_20), .B1 (n_0_213), .B2 (hfn_ipo_n29));
OAI22_X1 i_0_329 (.ZN (n_0_237), .A1 (n_0_188), .A2 (n_0_61), .B1 (drc_ipo_n33), .B2 (n_0_236));
AOI22_X1 i_0_328 (.ZN (n_0_236), .A1 (n_0_235), .A2 (n_0_109), .B1 (n_0_136), .B2 (n_0_16));
NAND2_X2 i_0_327 (.ZN (n_0_235), .A1 (n_0_233), .A2 (n_0_234));
AOI22_X1 i_0_326 (.ZN (n_0_234), .A1 (n_0_89), .A2 (\Input1_1_Negative[25] ), .B1 (\Input1_2_Negative[25] ), .B2 (n_0_94));
AOI22_X1 i_0_325 (.ZN (n_0_233), .A1 (n_0_90), .A2 (\Input1_1_Positive[25] ), .B1 (n_0_92), .B2 (\Input1_2_Positive[25] ));
OAI22_X1 i_0_324 (.ZN (n_0_342__0), .A1 (n_0_232), .A2 (hfn_ipo_n32), .B1 (n_0_220), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_323 (.ZN (n_0_232), .A1 (n_0_231), .A2 (hfn_ipo_n26), .B1 (n_0_207), .B2 (hfn_ipo_n30));
OAI22_X1 i_0_322 (.ZN (n_0_231), .A1 (n_0_230), .A2 (drc_ipo_n33), .B1 (n_0_182), .B2 (n_0_17));
AOI22_X1 i_0_321 (.ZN (n_0_230), .A1 (n_0_229), .A2 (n_0_109), .B1 (n_0_129), .B2 (n_0_16));
NAND2_X1 i_0_320 (.ZN (n_0_229), .A1 (n_0_227), .A2 (n_0_228));
AOI22_X1 i_0_319 (.ZN (n_0_228), .A1 (n_0_89), .A2 (\Input1_2_Negative[25] ), .B1 (\Input1_1_Negative[23] ), .B2 (n_0_94));
AOI22_X1 i_0_318 (.ZN (n_0_227), .A1 (n_0_90), .A2 (\Input1_2_Positive[25] ), .B1 (n_0_92), .B2 (\Input1_1_Positive[23] ));
OAI22_X1 i_0_317 (.ZN (n_0_341__0), .A1 (n_0_214), .A2 (hfn_ipo_n28), .B1 (n_0_226), .B2 (hfn_ipo_n32));
AOI22_X1 i_0_316 (.ZN (n_0_226), .A1 (n_0_201), .A2 (hfn_ipo_n30), .B1 (n_0_225), .B2 (hfn_ipo_n26));
OAI22_X1 i_0_315 (.ZN (n_0_225), .A1 (n_0_224), .A2 (n_0_59), .B1 (n_0_131), .B2 (n_0_176));
OAI22_X1 i_0_314 (.ZN (n_0_224), .A1 (n_0_125), .A2 (n_0_28), .B1 (n_0_223), .B2 (\shiftingAmount[4] ));
NAND2_X1 i_0_313 (.ZN (n_0_223), .A1 (n_0_221), .A2 (n_0_222));
AOI22_X1 i_0_312 (.ZN (n_0_222), .A1 (n_0_90), .A2 (\Input1_1_Positive[23] ), .B1 (\Input1_2_Negative[23] ), .B2 (n_0_94));
AOI22_X1 i_0_311 (.ZN (n_0_221), .A1 (n_0_89), .A2 (\Input1_1_Negative[23] ), .B1 (\Input1_2_Positive[23] ), .B2 (n_0_92));
OAI22_X1 i_0_310 (.ZN (n_0_340__0), .A1 (n_0_220), .A2 (hfn_ipo_n32), .B1 (n_0_208), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_309 (.ZN (n_0_220), .A1 (n_0_195), .A2 (hfn_ipo_n30), .B1 (n_0_219), .B2 (hfn_ipo_n26));
OAI22_X1 i_0_308 (.ZN (n_0_219), .A1 (n_0_218), .A2 (n_0_59), .B1 (n_0_131), .B2 (n_0_169));
OAI22_X1 i_0_307 (.ZN (n_0_218), .A1 (n_0_119), .A2 (n_0_28), .B1 (n_0_217), .B2 (\shiftingAmount[4] ));
NAND2_X1 i_0_306 (.ZN (n_0_217), .A1 (n_0_215), .A2 (n_0_216));
AOI22_X1 i_0_305 (.ZN (n_0_216), .A1 (n_0_90), .A2 (\Input1_2_Positive[23] ), .B1 (\Input1_1_Negative[21] ), .B2 (n_0_94));
AOI22_X1 i_0_304 (.ZN (n_0_215), .A1 (n_0_89), .A2 (\Input1_2_Negative[23] ), .B1 (\Input1_1_Positive[21] ), .B2 (n_0_92));
OAI22_X1 i_0_303 (.ZN (n_0_339__0), .A1 (n_0_214), .A2 (hfn_ipo_n32), .B1 (hfn_ipo_n28), .B2 (n_0_202));
AOI22_X1 i_0_302 (.ZN (n_0_214), .A1 (n_0_189), .A2 (hfn_ipo_n29), .B1 (n_0_213), .B2 (n_0_20));
OAI22_X1 i_0_301 (.ZN (n_0_213), .A1 (n_0_212), .A2 (drc_ipo_n33), .B1 (n_0_131), .B2 (n_0_162));
AOI22_X1 i_0_300 (.ZN (n_0_212), .A1 (n_0_115), .A2 (n_0_16), .B1 (n_0_211), .B2 (n_0_109));
NAND2_X1 i_0_299 (.ZN (n_0_211), .A1 (n_0_209), .A2 (n_0_210));
AOI22_X1 i_0_298 (.ZN (n_0_210), .A1 (n_0_90), .A2 (\Input1_1_Positive[21] ), .B1 (\Input1_2_Positive[21] ), .B2 (n_0_92));
AOI22_X1 i_0_297 (.ZN (n_0_209), .A1 (n_0_89), .A2 (\Input1_1_Negative[21] ), .B1 (\Input1_2_Negative[21] ), .B2 (n_0_94));
OAI22_X1 i_0_296 (.ZN (n_0_338__0), .A1 (n_0_208), .A2 (hfn_ipo_n32), .B1 (n_0_196), .B2 (hfn_ipo_n28));
AOI22_X1 i_0_295 (.ZN (n_0_208), .A1 (n_0_207), .A2 (hfn_ipo_n26), .B1 (n_0_183), .B2 (hfn_ipo_n30));
OAI22_X1 i_0_294 (.ZN (n_0_207), .A1 (n_0_206), .A2 (drc_ipo_n33), .B1 (n_0_131), .B2 (n_0_156));
AOI22_X1 i_0_293 (.ZN (n_0_206), .A1 (n_0_205), .A2 (n_0_109), .B1 (n_0_105), .B2 (n_0_16));
NAND2_X1 i_0_292 (.ZN (n_0_205), .A1 (n_0_203), .A2 (n_0_204));
AOI22_X1 i_0_291 (.ZN (n_0_204), .A1 (n_0_90), .A2 (\Input1_2_Positive[21] ), .B1 (\Input1_1_Positive[19] ), .B2 (n_0_92));
AOI22_X1 i_0_290 (.ZN (n_0_203), .A1 (n_0_89), .A2 (\Input1_2_Negative[21] ), .B1 (\Input1_1_Negative[19] ), .B2 (n_0_94));
OAI22_X1 i_0_289 (.ZN (n_0_337__0), .A1 (n_0_190), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n31), .B2 (n_0_202));
AOI22_X1 i_0_288 (.ZN (n_0_202), .A1 (n_0_201), .A2 (n_0_20), .B1 (hfn_ipo_n29), .B2 (n_0_177));
OAI22_X1 i_0_287 (.ZN (n_0_201), .A1 (n_0_200), .A2 (n_0_59), .B1 (n_0_131), .B2 (n_0_149));
OAI22_X1 i_0_286 (.ZN (n_0_200), .A1 (n_0_101), .A2 (n_0_28), .B1 (n_0_199), .B2 (\shiftingAmount[4] ));
NAND2_X1 i_0_285 (.ZN (n_0_199), .A1 (n_0_197), .A2 (n_0_198));
AOI22_X1 i_0_284 (.ZN (n_0_198), .A1 (n_0_90), .A2 (\Input1_1_Positive[19] ), .B1 (\Input1_2_Negative[19] ), .B2 (n_0_94));
AOI22_X1 i_0_283 (.ZN (n_0_197), .A1 (n_0_89), .A2 (\Input1_1_Negative[19] ), .B1 (\Input1_2_Positive[19] ), .B2 (n_0_92));
OAI22_X1 i_0_282 (.ZN (n_0_336__0), .A1 (n_0_196), .A2 (hfn_ipo_n31), .B1 (n_0_184), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_281 (.ZN (n_0_196), .A1 (n_0_195), .A2 (n_0_20), .B1 (hfn_ipo_n29), .B2 (n_0_170));
OAI22_X1 i_0_280 (.ZN (n_0_195), .A1 (n_0_194), .A2 (n_0_59), .B1 (n_0_131), .B2 (n_0_143));
OAI22_X1 i_0_279 (.ZN (n_0_194), .A1 (n_0_96), .A2 (n_0_28), .B1 (n_0_193), .B2 (\shiftingAmount[4] ));
NAND2_X1 i_0_278 (.ZN (n_0_193), .A1 (n_0_191), .A2 (n_0_192));
AOI22_X1 i_0_277 (.ZN (n_0_192), .A1 (n_0_90), .A2 (\Input1_2_Positive[19] ), .B1 (\Input1_1_Positive[17] ), .B2 (n_0_92));
AOI22_X1 i_0_276 (.ZN (n_0_191), .A1 (n_0_89), .A2 (\Input1_2_Negative[19] ), .B1 (\Input1_1_Negative[17] ), .B2 (n_0_94));
OAI22_X1 i_0_275 (.ZN (n_0_335__0), .A1 (n_0_190), .A2 (hfn_ipo_n31), .B1 (hfn_ipo_n27), .B2 (n_0_178));
AOI22_X1 i_0_274 (.ZN (n_0_190), .A1 (n_0_189), .A2 (n_0_20), .B1 (hfn_ipo_n29), .B2 (n_0_164));
OAI22_X1 i_0_273 (.ZN (n_0_189), .A1 (n_0_188), .A2 (n_0_59), .B1 (n_0_131), .B2 (n_0_137));
OAI22_X1 i_0_272 (.ZN (n_0_188), .A1 (n_0_112), .A2 (n_0_28), .B1 (n_0_187), .B2 (\shiftingAmount[4] ));
NAND2_X1 i_0_271 (.ZN (n_0_187), .A1 (n_0_185), .A2 (n_0_186));
AOI22_X1 i_0_270 (.ZN (n_0_186), .A1 (n_0_90), .A2 (\Input1_1_Positive[17] ), .B1 (\Input1_2_Positive[17] ), .B2 (n_0_92));
AOI22_X1 i_0_269 (.ZN (n_0_185), .A1 (n_0_89), .A2 (\Input1_1_Negative[17] ), .B1 (\Input1_2_Negative[17] ), .B2 (n_0_94));
OAI22_X1 i_0_268 (.ZN (n_0_334__0), .A1 (n_0_184), .A2 (hfn_ipo_n31), .B1 (n_0_171), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_267 (.ZN (n_0_184), .A1 (n_0_183), .A2 (n_0_20), .B1 (hfn_ipo_n29), .B2 (n_0_157));
OAI22_X1 i_0_266 (.ZN (n_0_183), .A1 (n_0_182), .A2 (drc_ipo_n33), .B1 (n_0_131), .B2 (n_0_130));
AOI22_X1 i_0_265 (.ZN (n_0_182), .A1 (n_0_181), .A2 (n_0_109), .B1 (n_0_16), .B2 (n_0_108));
NAND2_X1 i_0_264 (.ZN (n_0_181), .A1 (n_0_179), .A2 (n_0_180));
AOI22_X1 i_0_263 (.ZN (n_0_180), .A1 (n_0_90), .A2 (\Input1_2_Positive[17] ), .B1 (\Input1_1_Positive[15] ), .B2 (n_0_92));
AOI22_X1 i_0_262 (.ZN (n_0_179), .A1 (n_0_89), .A2 (\Input1_2_Negative[17] ), .B1 (\Input1_1_Negative[15] ), .B2 (n_0_94));
OAI22_X1 i_0_261 (.ZN (n_0_333__0), .A1 (n_0_165), .A2 (hfn_ipo_n27), .B1 (n_0_178), .B2 (hfn_ipo_n31));
AOI22_X1 i_0_260 (.ZN (n_0_178), .A1 (n_0_177), .A2 (n_0_20), .B1 (n_0_150), .B2 (hfn_ipo_n29));
OAI22_X1 i_0_259 (.ZN (n_0_177), .A1 (n_0_172), .A2 (n_0_131), .B1 (n_0_176), .B2 (n_0_106));
INV_X1 i_0_258 (.ZN (n_0_176), .A (n_0_175));
NAND2_X1 i_0_257 (.ZN (n_0_175), .A1 (n_0_173), .A2 (n_0_174));
AOI22_X1 i_0_256 (.ZN (n_0_174), .A1 (n_0_90), .A2 (\Input1_1_Positive[15] ), .B1 (\Input1_2_Positive[15] ), .B2 (n_0_92));
AOI22_X1 i_0_255 (.ZN (n_0_173), .A1 (n_0_89), .A2 (\Input1_1_Negative[15] ), .B1 (\Input1_2_Negative[15] ), .B2 (n_0_94));
INV_X1 i_0_254 (.ZN (n_0_172), .A (n_0_125));
OAI22_X1 i_0_253 (.ZN (n_0_332__0), .A1 (n_0_171), .A2 (hfn_ipo_n31), .B1 (n_0_158), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_252 (.ZN (n_0_171), .A1 (n_0_144), .A2 (hfn_ipo_n29), .B1 (n_0_170), .B2 (n_0_20));
OAI22_X1 i_0_251 (.ZN (n_0_170), .A1 (n_0_120), .A2 (n_0_131), .B1 (n_0_169), .B2 (n_0_106));
INV_X1 i_0_250 (.ZN (n_0_169), .A (n_0_168));
NAND2_X1 i_0_249 (.ZN (n_0_168), .A1 (n_0_166), .A2 (n_0_167));
AOI22_X1 i_0_248 (.ZN (n_0_167), .A1 (n_0_90), .A2 (\Input1_2_Positive[15] ), .B1 (\Input1_1_Positive[13] ), .B2 (n_0_92));
AOI22_X1 i_0_247 (.ZN (n_0_166), .A1 (n_0_89), .A2 (\Input1_2_Negative[15] ), .B1 (\Input1_1_Negative[13] ), .B2 (n_0_94));
OAI22_X1 i_0_246 (.ZN (n_0_331__0), .A1 (n_0_165), .A2 (hfn_ipo_n31), .B1 (n_0_151), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_245 (.ZN (n_0_165), .A1 (n_0_138), .A2 (hfn_ipo_n29), .B1 (n_0_164), .B2 (n_0_20));
OAI22_X1 i_0_244 (.ZN (n_0_164), .A1 (n_0_162), .A2 (n_0_106), .B1 (n_0_163), .B2 (n_0_131));
INV_X1 i_0_243 (.ZN (n_0_163), .A (n_0_115));
INV_X1 i_0_242 (.ZN (n_0_162), .A (n_0_161));
NAND2_X1 i_0_241 (.ZN (n_0_161), .A1 (n_0_159), .A2 (n_0_160));
AOI22_X1 i_0_240 (.ZN (n_0_160), .A1 (n_0_89), .A2 (\Input1_1_Negative[13] ), .B1 (\Input1_2_Negative[13] ), .B2 (n_0_94));
AOI22_X1 i_0_239 (.ZN (n_0_159), .A1 (n_0_90), .A2 (\Input1_1_Positive[13] ), .B1 (n_0_92), .B2 (\Input1_2_Positive[13] ));
OAI22_X1 i_0_238 (.ZN (n_0_330__0), .A1 (n_0_158), .A2 (hfn_ipo_n31), .B1 (n_0_145), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_237 (.ZN (n_0_158), .A1 (n_0_157), .A2 (n_0_20), .B1 (n_0_132), .B2 (hfn_ipo_n29));
OAI22_X1 i_0_236 (.ZN (n_0_157), .A1 (n_0_152), .A2 (n_0_131), .B1 (n_0_156), .B2 (n_0_106));
INV_X1 i_0_235 (.ZN (n_0_156), .A (n_0_155));
NAND2_X1 i_0_234 (.ZN (n_0_155), .A1 (n_0_153), .A2 (n_0_154));
AOI22_X1 i_0_233 (.ZN (n_0_154), .A1 (n_0_90), .A2 (\Input1_2_Positive[13] ), .B1 (\Input1_1_Negative[11] ), .B2 (n_0_94));
AOI22_X1 i_0_232 (.ZN (n_0_153), .A1 (n_0_89), .A2 (\Input1_2_Negative[13] ), .B1 (\Input1_1_Positive[11] ), .B2 (n_0_92));
INV_X1 i_0_231 (.ZN (n_0_152), .A (n_0_105));
OAI22_X1 i_0_230 (.ZN (n_0_329__0), .A1 (n_0_139), .A2 (hfn_ipo_n27), .B1 (n_0_151), .B2 (hfn_ipo_n31));
AOI22_X1 i_0_229 (.ZN (n_0_151), .A1 (n_0_150), .A2 (n_0_20), .B1 (n_0_125), .B2 (n_0_110));
OAI22_X1 i_0_228 (.ZN (n_0_150), .A1 (n_0_149), .A2 (n_0_106), .B1 (n_0_102), .B2 (n_0_131));
INV_X1 i_0_227 (.ZN (n_0_149), .A (n_0_148));
NAND2_X1 i_0_226 (.ZN (n_0_148), .A1 (n_0_146), .A2 (n_0_147));
AOI22_X1 i_0_225 (.ZN (n_0_147), .A1 (n_0_90), .A2 (\Input1_1_Positive[11] ), .B1 (\Input1_2_Negative[11] ), .B2 (n_0_94));
AOI22_X1 i_0_224 (.ZN (n_0_146), .A1 (n_0_89), .A2 (\Input1_1_Negative[11] ), .B1 (n_0_92), .B2 (\Input1_2_Positive[11] ));
OAI22_X1 i_0_223 (.ZN (n_0_328__0), .A1 (n_0_145), .A2 (hfn_ipo_n31), .B1 (n_0_133), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_222 (.ZN (n_0_145), .A1 (n_0_144), .A2 (n_0_20), .B1 (n_0_121), .B2 (hfn_ipo_n29));
OAI22_X1 i_0_221 (.ZN (n_0_144), .A1 (n_0_97), .A2 (n_0_131), .B1 (n_0_143), .B2 (n_0_106));
INV_X1 i_0_220 (.ZN (n_0_143), .A (n_0_142));
NAND2_X1 i_0_219 (.ZN (n_0_142), .A1 (n_0_140), .A2 (n_0_141));
AOI22_X1 i_0_218 (.ZN (n_0_141), .A1 (n_0_90), .A2 (\Input1_2_Positive[11] ), .B1 (\Input1_1_Negative[9] ), .B2 (n_0_94));
AOI22_X1 i_0_217 (.ZN (n_0_140), .A1 (n_0_89), .A2 (\Input1_2_Negative[11] ), .B1 (\Input1_1_Positive[9] ), .B2 (n_0_92));
OAI22_X1 i_0_216 (.ZN (n_0_327__0), .A1 (n_0_139), .A2 (hfn_ipo_n31), .B1 (hfn_ipo_n27), .B2 (n_0_126));
AOI22_X1 i_0_215 (.ZN (n_0_139), .A1 (n_0_138), .A2 (n_0_20), .B1 (n_0_110), .B2 (n_0_115));
OAI22_X1 i_0_214 (.ZN (n_0_138), .A1 (n_0_91), .A2 (n_0_131), .B1 (n_0_137), .B2 (n_0_106));
INV_X1 i_0_213 (.ZN (n_0_137), .A (n_0_136));
NAND2_X1 i_0_212 (.ZN (n_0_136), .A1 (n_0_134), .A2 (n_0_135));
AOI22_X1 i_0_211 (.ZN (n_0_135), .A1 (n_0_89), .A2 (\Input1_1_Negative[9] ), .B1 (\Input1_2_Negative[9] ), .B2 (n_0_94));
AOI22_X1 i_0_210 (.ZN (n_0_134), .A1 (n_0_90), .A2 (\Input1_1_Positive[9] ), .B1 (\Input1_2_Positive[9] ), .B2 (n_0_92));
OAI22_X1 i_0_209 (.ZN (n_0_326__0), .A1 (n_0_133), .A2 (hfn_ipo_n31), .B1 (n_0_122), .B2 (hfn_ipo_n27));
AOI22_X1 i_0_208 (.ZN (n_0_133), .A1 (n_0_132), .A2 (n_0_20), .B1 (n_0_105), .B2 (n_0_110));
OAI22_X1 i_0_207 (.ZN (n_0_132), .A1 (n_0_130), .A2 (n_0_106), .B1 (n_0_131), .B2 (n_0_70));
INV_X1 i_0_206 (.ZN (n_0_131), .A (n_0_62));
INV_X1 i_0_205 (.ZN (n_0_130), .A (n_0_129));
NAND2_X1 i_0_204 (.ZN (n_0_129), .A1 (n_0_127), .A2 (n_0_128));
AOI22_X1 i_0_203 (.ZN (n_0_128), .A1 (n_0_89), .A2 (\Input1_2_Negative[9] ), .B1 (\Input1_1_Negative[7] ), .B2 (n_0_94));
AOI22_X1 i_0_202 (.ZN (n_0_127), .A1 (n_0_90), .A2 (\Input1_2_Positive[9] ), .B1 (\Input1_1_Positive[7] ), .B2 (n_0_92));
OAI22_X1 i_0_201 (.ZN (n_0_325__0), .A1 (n_0_116), .A2 (hfn_ipo_n27), .B1 (hfn_ipo_n31), .B2 (n_0_126));
AOI22_X1 i_0_200 (.ZN (n_0_126), .A1 (n_0_125), .A2 (n_0_107), .B1 (n_0_101), .B2 (n_0_110));
NAND2_X1 i_0_199 (.ZN (n_0_125), .A1 (n_0_123), .A2 (n_0_124));
AOI22_X1 i_0_198 (.ZN (n_0_124), .A1 (n_0_89), .A2 (\Input1_1_Negative[7] ), .B1 (\Input1_2_Negative[7] ), .B2 (n_0_94));
AOI22_X1 i_0_197 (.ZN (n_0_123), .A1 (n_0_90), .A2 (\Input1_1_Positive[7] ), .B1 (\Input1_2_Positive[7] ), .B2 (n_0_92));
OAI22_X1 i_0_196 (.ZN (n_0_324__0), .A1 (n_0_122), .A2 (hfn_ipo_n31), .B1 (hfn_ipo_n27), .B2 (n_0_111));
AOI22_X1 i_0_195 (.ZN (n_0_122), .A1 (n_0_121), .A2 (n_0_20), .B1 (n_0_96), .B2 (n_0_110));
NOR2_X1 i_0_194 (.ZN (n_0_121), .A1 (n_0_120), .A2 (n_0_106));
INV_X1 i_0_193 (.ZN (n_0_120), .A (n_0_119));
NAND2_X1 i_0_192 (.ZN (n_0_119), .A1 (n_0_117), .A2 (n_0_118));
AOI22_X1 i_0_191 (.ZN (n_0_118), .A1 (n_0_90), .A2 (\Input1_2_Positive[7] ), .B1 (\Input1_1_Negative[5] ), .B2 (n_0_94));
AOI22_X1 i_0_190 (.ZN (n_0_117), .A1 (n_0_89), .A2 (\Input1_2_Negative[7] ), .B1 (\Input1_1_Positive[5] ), .B2 (n_0_92));
OAI22_X1 i_0_189 (.ZN (n_0_323__0), .A1 (n_0_116), .A2 (hfn_ipo_n31), .B1 (n_0_102), .B2 (n_0_98));
AOI22_X1 i_0_188 (.ZN (n_0_116), .A1 (n_0_112), .A2 (n_0_110), .B1 (n_0_107), .B2 (n_0_115));
NAND2_X1 i_0_187 (.ZN (n_0_115), .A1 (n_0_113), .A2 (n_0_114));
AOI22_X1 i_0_186 (.ZN (n_0_114), .A1 (n_0_90), .A2 (\Input1_1_Positive[5] ), .B1 (\Input1_2_Negative[5] ), .B2 (n_0_94));
AOI22_X1 i_0_185 (.ZN (n_0_113), .A1 (n_0_89), .A2 (\Input1_1_Negative[5] ), .B1 (\Input1_2_Positive[5] ), .B2 (n_0_92));
INV_X1 i_0_184 (.ZN (n_0_112), .A (n_0_91));
OAI22_X1 i_0_183 (.ZN (n_0_322__0), .A1 (n_0_111), .A2 (hfn_ipo_n31), .B1 (n_0_97), .B2 (n_0_98));
AOI22_X1 i_0_182 (.ZN (n_0_111), .A1 (n_0_105), .A2 (n_0_107), .B1 (n_0_108), .B2 (n_0_110));
AND2_X1 i_0_181 (.ZN (n_0_110), .A1 (n_0_30), .A2 (n_0_109));
NOR2_X2 i_0_180 (.ZN (n_0_109), .A1 (\shiftingAmount[4] ), .A2 (drc_ipo_n34));
INV_X1 i_0_179 (.ZN (n_0_108), .A (n_0_70));
NOR2_X1 i_0_178 (.ZN (n_0_107), .A1 (n_0_106), .A2 (hfn_ipo_n29));
INV_X1 i_0_177 (.ZN (n_0_106), .A (n_0_60));
NAND2_X1 i_0_176 (.ZN (n_0_105), .A1 (n_0_103), .A2 (n_0_104));
AOI22_X1 i_0_175 (.ZN (n_0_104), .A1 (n_0_89), .A2 (\Input1_2_Negative[5] ), .B1 (\Input1_1_Negative[3] ), .B2 (n_0_94));
AOI22_X1 i_0_174 (.ZN (n_0_103), .A1 (n_0_90), .A2 (\Input1_2_Positive[5] ), .B1 (\Input1_1_Positive[3] ), .B2 (n_0_92));
OAI22_X1 i_0_173 (.ZN (n_0_321__0), .A1 (n_0_91), .A2 (n_0_98), .B1 (n_0_71), .B2 (n_0_102));
INV_X1 i_0_172 (.ZN (n_0_102), .A (n_0_101));
NAND2_X1 i_0_171 (.ZN (n_0_101), .A1 (n_0_99), .A2 (n_0_100));
AOI22_X1 i_0_170 (.ZN (n_0_100), .A1 (n_0_89), .A2 (\Input1_1_Negative[3] ), .B1 (\Input1_2_Negative[3] ), .B2 (n_0_94));
AOI22_X1 i_0_169 (.ZN (n_0_99), .A1 (n_0_90), .A2 (\Input1_1_Positive[3] ), .B1 (\Input1_2_Positive[3] ), .B2 (n_0_92));
OAI22_X1 i_0_168 (.ZN (n_0_320__0), .A1 (n_0_97), .A2 (n_0_71), .B1 (n_0_70), .B2 (n_0_98));
NAND2_X1 i_0_167 (.ZN (n_0_98), .A1 (n_0_60), .A2 (n_0_22));
INV_X4 i_0_166 (.ZN (n_0_97), .A (n_0_96));
NAND2_X2 i_0_165 (.ZN (n_0_96), .A1 (n_0_93), .A2 (n_0_95));
AOI22_X1 i_0_164 (.ZN (n_0_95), .A1 (n_0_89), .A2 (\Input1_2_Negative[3] ), .B1 (\Input1_1_Negative[1] ), .B2 (n_0_94));
INV_X2 i_0_163 (.ZN (n_0_94), .A (n_0_86));
AOI22_X1 i_0_162 (.ZN (n_0_93), .A1 (n_0_90), .A2 (\Input1_2_Positive[3] ), .B1 (\Input1_1_Positive[1] ), .B2 (n_0_92));
INV_X2 i_0_161 (.ZN (n_0_92), .A (n_0_87));
NOR2_X2 i_0_160 (.ZN (n_0_318__0), .A1 (n_0_91), .A2 (n_0_71));
AOI221_X2 i_0_159 (.ZN (n_0_91), .A (n_0_88), .B1 (n_0_89), .B2 (\Input1_1_Negative[1] )
    , .C1 (\Input1_1_Positive[1] ), .C2 (n_0_90));
NOR2_X4 i_0_158 (.ZN (n_0_90), .A1 (n_0_68), .A2 (n_0_85));
NOR2_X4 i_0_157 (.ZN (n_0_89), .A1 (n_0_68), .A2 (n_0_84));
AOI21_X1 i_0_156 (.ZN (n_0_88), .A (n_0_69), .B1 (n_0_86), .B2 (n_0_87));
NAND3_X1 i_0_155 (.ZN (n_0_87), .A1 (n_0_44), .A2 (n_0_66), .A3 (n_0_84));
NAND3_X1 i_0_154 (.ZN (n_0_86), .A1 (n_0_67), .A2 (n_0_65), .A3 (n_0_85));
INV_X1 i_0_153 (.ZN (n_0_85), .A (n_0_84));
AOI211_X2 i_0_152 (.ZN (n_0_84), .A (n_0_72), .B (n_0_75), .C1 (n_0_83), .C2 (n_0_8));
OAI22_X1 i_0_151 (.ZN (n_0_83), .A1 (n_0_51), .A2 (hfn_ipo_n31), .B1 (n_0_82), .B2 (hfn_ipo_n27));
AOI222_X1 i_0_150 (.ZN (n_0_82), .A1 (n_0_77), .A2 (\shiftingAmount[4] ), .B1 (n_0_80)
    , .B2 (n_0_9), .C1 (n_0_81), .C2 (n_0_34));
AOI22_X1 i_0_149 (.ZN (n_0_81), .A1 (n_0_55), .A2 (n_0_28), .B1 (n_0_13), .B2 (\shiftingAmount[4] ));
OAI22_X1 i_0_148 (.ZN (n_0_80), .A1 (n_0_78), .A2 (n_0_20), .B1 (n_0_79), .B2 (hfn_ipo_n29));
INV_X1 i_0_147 (.ZN (n_0_79), .A (\newB[4] ));
INV_X1 i_0_146 (.ZN (n_0_78), .A (\newB[8] ));
OAI22_X1 i_0_145 (.ZN (n_0_77), .A1 (n_0_31), .A2 (n_0_76), .B1 (n_0_29), .B2 (n_0_54));
INV_X1 i_0_144 (.ZN (n_0_76), .A (\newB[28] ));
OAI211_X1 i_0_143 (.ZN (n_0_75), .A (n_0_14), .B (n_0_73), .C1 (n_0_23), .C2 (n_0_74));
NAND2_X1 i_0_142 (.ZN (n_0_74), .A1 (n_0_58), .A2 (\newB[20] ));
NAND3_X1 i_0_141 (.ZN (n_0_73), .A1 (n_0_62), .A2 (\newB[12] ), .A3 (n_0_22));
NOR3_X1 i_0_140 (.ZN (n_0_72), .A1 (n_0_45), .A2 (n_0_12), .A3 (n_0_15));
NOR2_X1 i_0_139 (.ZN (n_0_316__0), .A1 (n_0_70), .A2 (n_0_71));
NAND2_X1 i_0_138 (.ZN (n_0_71), .A1 (n_0_60), .A2 (n_0_11));
OR2_X1 i_0_137 (.ZN (n_0_70), .A1 (n_0_68), .A2 (n_0_69));
INV_X1 i_0_136 (.ZN (n_0_69), .A (\Input1_2_Positive[1] ));
OAI22_X2 i_0_135 (.ZN (n_0_68), .A1 (n_0_44), .A2 (n_0_66), .B1 (n_0_67), .B2 (n_0_65));
INV_X1 i_0_134 (.ZN (n_0_67), .A (n_0_44));
INV_X1 i_0_133 (.ZN (n_0_66), .A (n_0_65));
AOI221_X2 i_0_132 (.ZN (n_0_65), .A (n_0_46), .B1 (n_0_8), .B2 (n_0_53), .C1 (n_0_64), .C2 (hfn_ipo_n27));
OAI22_X1 i_0_131 (.ZN (n_0_64), .A1 (n_0_57), .A2 (n_0_15), .B1 (n_0_20), .B2 (n_0_63));
AOI22_X1 i_0_130 (.ZN (n_0_63), .A1 (\newB[4] ), .A2 (n_0_60), .B1 (n_0_62), .B2 (\newB[12] ));
NOR2_X1 i_0_129 (.ZN (n_0_62), .A1 (n_0_61), .A2 (\shiftingAmount[4] ));
NAND2_X1 i_0_128 (.ZN (n_0_61), .A1 (n_0_8), .A2 (drc_ipo_n33));
NOR2_X1 i_0_127 (.ZN (n_0_60), .A1 (n_0_59), .A2 (\shiftingAmount[4] ));
INV_X1 i_0_126 (.ZN (n_0_59), .A (n_0_58));
NOR2_X1 i_0_125 (.ZN (n_0_58), .A1 (drc_ipo_n33), .A2 (drc_ipo_n34));
AOI221_X1 i_0_124 (.ZN (n_0_57), .A (n_0_56), .B1 (\newB[20] ), .B2 (n_0_30), .C1 (\newB[28] ), .C2 (n_0_34));
AOI221_X1 i_0_123 (.ZN (n_0_56), .A (hfn_ipo_n29), .B1 (n_0_54), .B2 (drc_ipo_n33)
    , .C1 (n_0_55), .C2 (n_0_17));
INV_X1 i_0_122 (.ZN (n_0_55), .A (\newB[16] ));
INV_X1 i_0_121 (.ZN (n_0_54), .A (\newB[24] ));
OAI22_X1 i_0_120 (.ZN (n_0_53), .A1 (n_0_51), .A2 (hfn_ipo_n27), .B1 (n_0_12), .B2 (n_0_52));
NAND2_X1 i_0_119 (.ZN (n_0_52), .A1 (n_0_25), .A2 (\newB[8] ));
INV_X1 i_0_118 (.ZN (n_0_51), .A (n_0_50));
OAI222_X1 i_0_117 (.ZN (n_0_50), .A1 (\shiftingAmount[4] ), .A2 (n_0_47), .B1 (n_0_48)
    , .B2 (n_0_28), .C1 (n_0_49), .C2 (hfn_ipo_n29));
AOI22_X1 i_0_116 (.ZN (n_0_49), .A1 (n_0_25), .A2 (\newB[10] ), .B1 (n_0_9), .B2 (\newB[2] ));
AOI22_X1 i_0_115 (.ZN (n_0_48), .A1 (n_0_34), .A2 (\newB[30] ), .B1 (n_0_30), .B2 (\newB[22] ));
AOI22_X1 i_0_114 (.ZN (n_0_47), .A1 (n_0_34), .A2 (\newB[14] ), .B1 (n_0_30), .B2 (\newB[6] ));
OAI33_X1 i_0_113 (.ZN (n_0_46), .A1 (n_0_10), .A2 (n_0_13), .A3 (hfn_ipo_n29), .B1 (n_0_45)
    , .B2 (n_0_15), .B3 (n_0_21));
AOI22_X1 i_0_112 (.ZN (n_0_45), .A1 (n_0_17), .A2 (\newB[18] ), .B1 (\newB[26] ), .B2 (drc_ipo_n33));
OAI211_X2 i_0_111 (.ZN (n_0_44), .A (n_0_14), .B (n_0_18), .C1 (n_0_43), .C2 (drc_ipo_n34));
AOI211_X1 i_0_110 (.ZN (n_0_43), .A (n_0_27), .B (n_0_40), .C1 (hfn_ipo_n31), .C2 (n_0_42));
NOR2_X1 i_0_109 (.ZN (n_0_42), .A1 (n_0_41), .A2 (n_0_28));
AOI22_X1 i_0_108 (.ZN (n_0_41), .A1 (n_0_34), .A2 (\newB[31] ), .B1 (n_0_30), .B2 (\newB[23] ));
OAI33_X1 i_0_107 (.ZN (n_0_40), .A1 (n_0_33), .A2 (n_0_35), .A3 (hfn_ipo_n31), .B1 (n_0_37)
    , .B2 (n_0_39), .B3 (n_0_20));
AOI221_X1 i_0_106 (.ZN (n_0_39), .A (hfn_ipo_n27), .B1 (n_0_9), .B2 (\newB[7] ), .C1 (n_0_25), .C2 (\newB[15] ));
INV_X1 i_0_105 (.ZN (n_0_38), .A (hfn_ipo_n32));
AOI211_X1 i_0_104 (.ZN (n_0_37), .A (hfn_ipo_n31), .B (n_0_36), .C1 (\newB[5] ), .C2 (n_0_9));
AND3_X1 i_0_103 (.ZN (n_0_36), .A1 (\newB[29] ), .A2 (\shiftingAmount[4] ), .A3 (drc_ipo_n33));
AOI221_X1 i_0_102 (.ZN (n_0_35), .A (\shiftingAmount[4] ), .B1 (n_0_32), .B2 (\newB[9] )
    , .C1 (\newB[13] ), .C2 (n_0_34));
NOR2_X1 i_0_101 (.ZN (n_0_34), .A1 (n_0_17), .A2 (n_0_20));
AOI221_X1 i_0_100 (.ZN (n_0_33), .A (n_0_28), .B1 (n_0_30), .B2 (\newB[21] ), .C1 (\newB[25] ), .C2 (n_0_32));
INV_X1 i_0_99 (.ZN (n_0_32), .A (n_0_31));
NAND2_X1 i_0_98 (.ZN (n_0_31), .A1 (n_0_20), .A2 (drc_ipo_n33));
INV_X1 i_0_97 (.ZN (n_0_30), .A (n_0_29));
NAND2_X1 i_0_96 (.ZN (n_0_29), .A1 (n_0_17), .A2 (hfn_ipo_n29));
INV_X1 i_0_95 (.ZN (n_0_28), .A (\shiftingAmount[4] ));
OAI221_X1 i_0_94 (.ZN (n_0_27), .A (n_0_19), .B1 (n_0_23), .B2 (n_0_24), .C1 (n_0_26), .C2 (n_0_21));
AOI22_X1 i_0_93 (.ZN (n_0_26), .A1 (n_0_25), .A2 (\newB[11] ), .B1 (n_0_9), .B2 (\newB[3] ));
NOR2_X1 i_0_92 (.ZN (n_0_25), .A1 (n_0_17), .A2 (\shiftingAmount[4] ));
OAI22_X1 i_0_91 (.ZN (n_0_24), .A1 (n_0_17), .A2 (\newB[27] ), .B1 (\newB[19] ), .B2 (drc_ipo_n33));
NAND2_X1 i_0_90 (.ZN (n_0_23), .A1 (n_0_22), .A2 (\shiftingAmount[4] ));
INV_X1 i_0_89 (.ZN (n_0_22), .A (n_0_21));
NAND2_X1 i_0_88 (.ZN (n_0_21), .A1 (n_0_20), .A2 (hfn_ipo_n31));
INV_X4 i_0_87 (.ZN (n_0_20), .A (hfn_ipo_n29));
NAND3_X1 i_0_86 (.ZN (n_0_19), .A1 (n_0_9), .A2 (n_0_11), .A3 (\newB[1] ));
NAND4_X1 i_0_85 (.ZN (n_0_18), .A1 (n_0_16), .A2 (n_0_11), .A3 (\newB[17] ), .A4 (n_0_17));
INV_X4 i_0_84 (.ZN (n_0_17), .A (drc_ipo_n33));
INV_X2 i_0_83 (.ZN (n_0_16), .A (n_0_15));
NAND2_X1 i_0_82 (.ZN (n_0_15), .A1 (n_0_8), .A2 (\shiftingAmount[4] ));
OR3_X1 i_0_81 (.ZN (n_0_14), .A1 (n_0_10), .A2 (n_0_12), .A3 (n_0_13));
INV_X1 i_0_80 (.ZN (n_0_13), .A (\newB[34] ));
NOR3_X1 i_0_79 (.ZN (n_168), .A1 (n_0_10), .A2 (start), .A3 (n_0_12));
INV_X1 i_0_78 (.ZN (n_0_12), .A (n_0_11));
NOR2_X1 i_0_77 (.ZN (n_0_11), .A1 (hfn_ipo_n29), .A2 (hfn_ipo_n31));
NAND2_X1 i_0_76 (.ZN (n_0_10), .A1 (n_0_9), .A2 (drc_ipo_n34));
NOR2_X2 i_0_75 (.ZN (n_0_9), .A1 (\shiftingAmount[4] ), .A2 (drc_ipo_n33));
AOI221_X1 i_0_74 (.ZN (n_167), .A (CLOCK_slh_n239), .B1 (n_0_2), .B2 (drc_ipo_n34)
    , .C1 (n_0_7), .C2 (n_0_8));
INV_X4 i_0_73 (.ZN (n_0_8), .A (drc_ipo_n34));
INV_X1 i_0_72 (.ZN (n_0_7), .A (n_0_2));
AND2_X1 i_0_71 (.ZN (n_166), .A1 (hfn_ipo_n24), .A2 (n_0_5));
AND2_X1 i_0_70 (.ZN (n_165), .A1 (hfn_ipo_n24), .A2 (n_0_4));
AND2_X1 i_0_69 (.ZN (n_164), .A1 (hfn_ipo_n23), .A2 (n_0_3));
NOR2_X1 i_0_68 (.ZN (n_163), .A1 (CLOCK_slh_n239), .A2 (hfn_ipo_n31));
AND2_X1 i_0_67 (.ZN (n_162), .A1 (hfn_ipo_n24), .A2 (n_95));
AND2_X1 i_0_66 (.ZN (n_161), .A1 (hfn_ipo_n24), .A2 (n_94));
AND2_X1 i_0_65 (.ZN (n_160), .A1 (hfn_ipo_n24), .A2 (n_93));
AND2_X1 i_0_64 (.ZN (n_159), .A1 (hfn_ipo_n24), .A2 (n_92));
AND2_X1 i_0_63 (.ZN (n_158), .A1 (hfn_ipo_n24), .A2 (n_91));
AND2_X1 i_0_62 (.ZN (n_157), .A1 (hfn_ipo_n24), .A2 (n_90));
AND2_X1 i_0_61 (.ZN (n_156), .A1 (hfn_ipo_n24), .A2 (n_89));
AND2_X1 i_0_60 (.ZN (n_155), .A1 (hfn_ipo_n24), .A2 (n_88));
AND2_X1 i_0_59 (.ZN (n_154), .A1 (hfn_ipo_n24), .A2 (n_87));
AND2_X1 i_0_58 (.ZN (n_153), .A1 (hfn_ipo_n24), .A2 (n_86));
AND2_X1 i_0_57 (.ZN (n_152), .A1 (hfn_ipo_n24), .A2 (n_85));
AND2_X1 i_0_56 (.ZN (n_151), .A1 (hfn_ipo_n24), .A2 (n_84));
AND2_X1 i_0_55 (.ZN (n_150), .A1 (hfn_ipo_n24), .A2 (n_83));
AND2_X1 i_0_54 (.ZN (n_149), .A1 (hfn_ipo_n24), .A2 (n_82));
AND2_X1 i_0_53 (.ZN (n_148), .A1 (hfn_ipo_n24), .A2 (n_81));
AND2_X1 i_0_52 (.ZN (n_144), .A1 (hfn_ipo_n24), .A2 (n_80));
AND2_X1 i_0_51 (.ZN (n_143), .A1 (hfn_ipo_n23), .A2 (n_79));
AND2_X1 i_0_50 (.ZN (n_142), .A1 (hfn_ipo_n23), .A2 (n_78));
AND2_X1 i_0_49 (.ZN (n_141), .A1 (hfn_ipo_n23), .A2 (n_77));
AND2_X1 i_0_48 (.ZN (n_140), .A1 (hfn_ipo_n23), .A2 (n_76));
AND2_X1 i_0_47 (.ZN (n_139), .A1 (hfn_ipo_n23), .A2 (n_75));
AND2_X1 i_0_46 (.ZN (n_138), .A1 (hfn_ipo_n23), .A2 (n_74));
AND2_X1 i_0_45 (.ZN (n_137), .A1 (hfn_ipo_n23), .A2 (n_73));
AND2_X1 i_0_44 (.ZN (n_136), .A1 (hfn_ipo_n23), .A2 (n_72));
AND2_X1 i_0_43 (.ZN (n_135), .A1 (hfn_ipo_n23), .A2 (n_71));
AND2_X1 i_0_42 (.ZN (n_134), .A1 (hfn_ipo_n23), .A2 (n_70));
AND2_X1 i_0_41 (.ZN (n_133), .A1 (hfn_ipo_n23), .A2 (n_69));
AND2_X1 i_0_40 (.ZN (n_132), .A1 (hfn_ipo_n23), .A2 (n_68));
AND2_X1 i_0_39 (.ZN (n_131), .A1 (hfn_ipo_n23), .A2 (n_67));
AND2_X1 i_0_38 (.ZN (n_130), .A1 (hfn_ipo_n24), .A2 (n_66));
AND2_X1 i_0_37 (.ZN (n_129), .A1 (hfn_ipo_n24), .A2 (n_65));
AND2_X1 i_0_36 (.ZN (n_128), .A1 (hfn_ipo_n24), .A2 (n_64));
AND2_X1 i_0_35 (.ZN (n_127), .A1 (hfn_ipo_n24), .A2 (n_32));
AND2_X1 i_0_34 (.ZN (n_126), .A1 (hfn_ipo_n24), .A2 (n_31));
AND2_X1 i_0_33 (.ZN (n_125), .A1 (hfn_ipo_n24), .A2 (n_30));
AND2_X1 i_0_32 (.ZN (n_124), .A1 (hfn_ipo_n24), .A2 (n_29));
AND2_X1 i_0_31 (.ZN (n_123), .A1 (hfn_ipo_n24), .A2 (n_28));
AND2_X1 i_0_30 (.ZN (n_122), .A1 (hfn_ipo_n24), .A2 (n_27));
AND2_X1 i_0_29 (.ZN (n_121), .A1 (hfn_ipo_n24), .A2 (n_26));
AND2_X1 i_0_28 (.ZN (n_120), .A1 (hfn_ipo_n24), .A2 (n_25));
AND2_X1 i_0_27 (.ZN (n_119), .A1 (hfn_ipo_n24), .A2 (n_24));
AND2_X1 i_0_26 (.ZN (n_118), .A1 (hfn_ipo_n24), .A2 (n_23));
AND2_X1 i_0_25 (.ZN (n_117), .A1 (hfn_ipo_n24), .A2 (n_22));
AND2_X1 i_0_24 (.ZN (n_116), .A1 (hfn_ipo_n24), .A2 (n_21));
AND2_X1 i_0_23 (.ZN (n_115), .A1 (hfn_ipo_n23), .A2 (n_20));
AND2_X1 i_0_22 (.ZN (n_114), .A1 (hfn_ipo_n23), .A2 (n_19));
AND2_X1 i_0_21 (.ZN (n_113), .A1 (hfn_ipo_n23), .A2 (n_18));
AND2_X1 i_0_20 (.ZN (n_112), .A1 (hfn_ipo_n23), .A2 (n_17));
AND2_X1 i_0_19 (.ZN (n_111), .A1 (hfn_ipo_n23), .A2 (n_16));
AND2_X1 i_0_18 (.ZN (n_110), .A1 (hfn_ipo_n23), .A2 (n_15));
AND2_X1 i_0_17 (.ZN (n_109), .A1 (hfn_ipo_n23), .A2 (n_14));
AND2_X1 i_0_16 (.ZN (n_108), .A1 (hfn_ipo_n23), .A2 (n_13));
AND2_X1 i_0_15 (.ZN (n_107), .A1 (hfn_ipo_n23), .A2 (n_12));
AND2_X1 i_0_14 (.ZN (n_106), .A1 (hfn_ipo_n23), .A2 (n_11));
AND2_X1 i_0_13 (.ZN (n_105), .A1 (hfn_ipo_n23), .A2 (n_10));
AND2_X1 i_0_12 (.ZN (n_104), .A1 (hfn_ipo_n23), .A2 (n_9));
AND2_X1 i_0_11 (.ZN (n_103), .A1 (hfn_ipo_n23), .A2 (n_8));
AND2_X1 i_0_10 (.ZN (n_102), .A1 (hfn_ipo_n23), .A2 (n_7));
AND2_X1 i_0_9 (.ZN (n_101), .A1 (hfn_ipo_n23), .A2 (n_6));
AND2_X1 i_0_8 (.ZN (n_100), .A1 (hfn_ipo_n23), .A2 (n_5));
AND2_X1 i_0_7 (.ZN (n_99), .A1 (hfn_ipo_n23), .A2 (n_4));
AND2_X1 i_0_6 (.ZN (n_98), .A1 (hfn_ipo_n23), .A2 (n_3));
AND2_X1 i_0_5 (.ZN (n_97), .A1 (hfn_ipo_n23), .A2 (n_2));
AND2_X1 i_0_4 (.ZN (n_96), .A1 (hfn_ipo_n23), .A2 (n_1));
INV_X1 i_0_3 (.ZN (n_0_6), .A (CLOCK_slh_n239));
HA_X1 i_0_2 (.CO (n_0_2), .S (n_0_5), .A (\shiftingAmount[4] ), .B (n_0_1));
HA_X1 i_0_1 (.CO (n_0_1), .S (n_0_4), .A (drc_ipo_n33), .B (n_0_0));
HA_X1 i_0_0 (.CO (n_0_0), .S (n_0_3), .A (hfn_ipo_n29), .B (hfn_ipo_n31));
datapath__0_12 i_12 (.p_1 ({n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, 
    n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, 
    n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_32, n_31, n_30, 
    n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
    n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, 
    n_2, n_1}), .p_0 ({n_0_381, n_0_380, n_0_379, n_0_378, n_0_377, n_0_376, n_0_375, 
    n_0_374, n_0_373, n_0_372, n_0_371__0, n_0_370__0, n_0_369__0, n_0_368__0, n_0_367__0, 
    n_0_366__0, n_0_365__0, n_0_364__0, n_0_363__0, n_0_362__0, n_0_361__0, n_0_360__0, 
    n_0_359__0, n_0_358__0, n_0_357__0, n_0_356__0, n_0_355__0, n_0_354__0, n_0_353__0, 
    n_0_352__0, n_0_351__0, n_0_350__0, n_0_349__0, n_0_348__0, n_0_347__0, n_0_346__0, 
    n_0_345__0, n_0_344__0, n_0_343__0, n_0_342__0, n_0_341__0, n_0_340__0, n_0_339__0, 
    n_0_338__0, n_0_337__0, n_0_336__0, n_0_335__0, n_0_334__0, n_0_333__0, n_0_332__0, 
    n_0_331__0, n_0_330__0, n_0_329__0, n_0_328__0, n_0_327__0, n_0_326__0, n_0_325__0, 
    n_0_324__0, n_0_323__0, n_0_322__0, n_0_321__0, n_0_320__0, n_0_318__0, n_0_316__0})
    , .tempResult ({\tempResult[63] , \tempResult[62] , \tempResult[61] , \tempResult[60] , 
    \tempResult[59] , \tempResult[58] , \tempResult[57] , \tempResult[56] , \tempResult[55] , 
    \tempResult[54] , \tempResult[53] , \tempResult[52] , \tempResult[51] , \tempResult[50] , 
    \tempResult[49] , \tempResult[48] , \tempResult[47] , \tempResult[46] , \tempResult[45] , 
    \tempResult[44] , \tempResult[43] , \tempResult[42] , \tempResult[41] , \tempResult[40] , 
    \tempResult[39] , \tempResult[38] , \tempResult[37] , \tempResult[36] , \tempResult[35] , 
    \tempResult[34] , \tempResult[33] , \tempResult[32] , \tempResult[31] , \tempResult[30] , 
    \tempResult[29] , \tempResult[28] , \tempResult[27] , \tempResult[26] , \tempResult[25] , 
    \tempResult[24] , \tempResult[23] , \tempResult[22] , \tempResult[21] , \tempResult[20] , 
    \tempResult[19] , \tempResult[18] , \tempResult[17] , \tempResult[16] , \tempResult[15] , 
    \tempResult[14] , \tempResult[13] , \tempResult[12] , \tempResult[11] , \tempResult[10] , 
    \tempResult[9] , \tempResult[8] , \tempResult[7] , \tempResult[6] , \tempResult[5] , 
    \tempResult[4] , \tempResult[3] , \tempResult[2] , \tempResult[1] , \tempResult[0] }));
datapath__0_0 i_2 (.p_0 ({n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
    n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
    n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, uc_0, uc_1}), .p_1 ({in1[31], 
    in1[30], in1[29], in1[28], in1[27], in1[26], in1[25], in1[24], in1[23], in1[22], 
    in1[21], in1[20], in1[19], in1[18], in1[17], in1[16], in1[15], in1[14], in1[13], 
    in1[12], in1[11], in1[10], in1[9], in1[8], in1[7], in1[6], in1[5], in1[4], in1[3], 
    in1[2], in1[1], in1[0], 1'b0 }));
DFF_X1 \result_reg[0]  (.Q (result[0]), .CK (CTS_n_tid0_142), .D (\tempResult[0] ));
DFF_X1 \result_reg[1]  (.Q (result[1]), .CK (CTS_n_tid0_142), .D (\tempResult[1] ));
DFF_X1 \result_reg[2]  (.Q (result[2]), .CK (CTS_n_tid0_142), .D (\tempResult[2] ));
DFF_X1 \result_reg[3]  (.Q (result[3]), .CK (CTS_n_tid0_142), .D (\tempResult[3] ));
DFF_X1 \result_reg[4]  (.Q (result[4]), .CK (CTS_n_tid0_142), .D (\tempResult[4] ));
DFF_X1 \result_reg[5]  (.Q (result[5]), .CK (CTS_n_tid0_142), .D (\tempResult[5] ));
DFF_X1 \result_reg[6]  (.Q (result[6]), .CK (CTS_n_tid0_142), .D (\tempResult[6] ));
DFF_X1 \result_reg[7]  (.Q (result[7]), .CK (CTS_n_tid0_142), .D (\tempResult[7] ));
DFF_X1 \result_reg[8]  (.Q (result[8]), .CK (CTS_n_tid0_142), .D (\tempResult[8] ));
DFF_X1 \result_reg[9]  (.Q (result[9]), .CK (CTS_n_tid0_142), .D (\tempResult[9] ));
DFF_X1 \result_reg[10]  (.Q (result[10]), .CK (CTS_n_tid0_142), .D (\tempResult[10] ));
DFF_X1 \result_reg[11]  (.Q (result[11]), .CK (CTS_n_tid0_142), .D (\tempResult[11] ));
DFF_X1 \result_reg[12]  (.Q (result[12]), .CK (CTS_n_tid0_142), .D (\tempResult[12] ));
DFF_X1 \result_reg[13]  (.Q (result[13]), .CK (CTS_n_tid0_142), .D (\tempResult[13] ));
DFF_X1 \result_reg[14]  (.Q (result[14]), .CK (CTS_n_tid0_142), .D (\tempResult[14] ));
DFF_X1 \result_reg[15]  (.Q (result[15]), .CK (CTS_n_tid0_142), .D (\tempResult[15] ));
DFF_X1 \result_reg[16]  (.Q (result[16]), .CK (CTS_n_tid0_142), .D (\tempResult[16] ));
DFF_X1 \result_reg[17]  (.Q (result[17]), .CK (CTS_n_tid0_142), .D (\tempResult[17] ));
DFF_X1 \result_reg[18]  (.Q (result[18]), .CK (CTS_n_tid0_142), .D (\tempResult[18] ));
DFF_X1 \result_reg[19]  (.Q (result[19]), .CK (CTS_n_tid0_142), .D (\tempResult[19] ));
DFF_X1 \result_reg[20]  (.Q (result[20]), .CK (CTS_n_tid0_142), .D (\tempResult[20] ));
DFF_X1 \result_reg[21]  (.Q (result[21]), .CK (CTS_n_tid0_142), .D (\tempResult[21] ));
DFF_X1 \result_reg[22]  (.Q (result[22]), .CK (CTS_n_tid0_142), .D (\tempResult[22] ));
DFF_X1 \result_reg[23]  (.Q (result[23]), .CK (CTS_n_tid0_142), .D (\tempResult[23] ));
DFF_X1 \result_reg[24]  (.Q (result[24]), .CK (CTS_n_tid0_142), .D (\tempResult[24] ));
DFF_X1 \result_reg[25]  (.Q (result[25]), .CK (CTS_n_tid0_142), .D (\tempResult[25] ));
DFF_X1 \result_reg[26]  (.Q (result[26]), .CK (CTS_n_tid0_142), .D (\tempResult[26] ));
DFF_X1 \result_reg[27]  (.Q (result[27]), .CK (CTS_n_tid0_142), .D (\tempResult[27] ));
DFF_X1 \result_reg[28]  (.Q (result[28]), .CK (CTS_n_tid0_142), .D (\tempResult[28] ));
DFF_X1 \result_reg[29]  (.Q (result[29]), .CK (CTS_n_tid0_142), .D (\tempResult[29] ));
DFF_X1 \result_reg[30]  (.Q (result[30]), .CK (CTS_n_tid0_142), .D (\tempResult[30] ));
DFF_X1 \result_reg[31]  (.Q (result[31]), .CK (CTS_n_tid0_142), .D (\tempResult[31] ));
DFF_X1 \result_reg[32]  (.Q (result[32]), .CK (CTS_n_tid0_142), .D (\tempResult[32] ));
DFF_X1 \result_reg[33]  (.Q (result[33]), .CK (CTS_n_tid0_142), .D (\tempResult[33] ));
DFF_X1 \result_reg[34]  (.Q (result[34]), .CK (CTS_n_tid0_142), .D (\tempResult[34] ));
DFF_X1 \result_reg[35]  (.Q (result[35]), .CK (CTS_n_tid0_142), .D (\tempResult[35] ));
DFF_X1 \result_reg[36]  (.Q (result[36]), .CK (CTS_n_tid0_142), .D (\tempResult[36] ));
DFF_X1 \result_reg[37]  (.Q (result[37]), .CK (CTS_n_tid0_142), .D (\tempResult[37] ));
DFF_X1 \result_reg[38]  (.Q (result[38]), .CK (CTS_n_tid0_142), .D (\tempResult[38] ));
DFF_X1 \result_reg[39]  (.Q (result[39]), .CK (CTS_n_tid0_142), .D (\tempResult[39] ));
DFF_X1 \result_reg[40]  (.Q (result[40]), .CK (CTS_n_tid0_142), .D (\tempResult[40] ));
DFF_X1 \result_reg[41]  (.Q (result[41]), .CK (CTS_n_tid0_142), .D (\tempResult[41] ));
DFF_X1 \result_reg[42]  (.Q (result[42]), .CK (CTS_n_tid0_142), .D (\tempResult[42] ));
DFF_X1 \result_reg[43]  (.Q (result[43]), .CK (CTS_n_tid0_142), .D (\tempResult[43] ));
DFF_X1 \result_reg[44]  (.Q (result[44]), .CK (CTS_n_tid0_142), .D (\tempResult[44] ));
DFF_X1 \result_reg[45]  (.Q (result[45]), .CK (CTS_n_tid0_142), .D (\tempResult[45] ));
DFF_X1 \result_reg[46]  (.Q (result[46]), .CK (CTS_n_tid0_142), .D (\tempResult[46] ));
DFF_X1 \result_reg[47]  (.Q (result[47]), .CK (CTS_n_tid0_142), .D (\tempResult[47] ));
DFF_X1 \result_reg[48]  (.Q (result[48]), .CK (CTS_n_tid0_142), .D (\tempResult[48] ));
DFF_X1 \result_reg[49]  (.Q (result[49]), .CK (CTS_n_tid0_142), .D (\tempResult[49] ));
DFF_X1 \result_reg[50]  (.Q (result[50]), .CK (CTS_n_tid0_142), .D (\tempResult[50] ));
DFF_X1 \result_reg[51]  (.Q (result[51]), .CK (CTS_n_tid0_142), .D (\tempResult[51] ));
DFF_X1 \result_reg[52]  (.Q (result[52]), .CK (CTS_n_tid0_142), .D (\tempResult[52] ));
DFF_X1 \result_reg[53]  (.Q (result[53]), .CK (CTS_n_tid0_142), .D (\tempResult[53] ));
DFF_X1 \result_reg[54]  (.Q (result[54]), .CK (CTS_n_tid0_142), .D (\tempResult[54] ));
DFF_X1 \result_reg[55]  (.Q (result[55]), .CK (CTS_n_tid0_142), .D (\tempResult[55] ));
DFF_X1 \result_reg[56]  (.Q (result[56]), .CK (CTS_n_tid0_142), .D (\tempResult[56] ));
DFF_X1 \result_reg[57]  (.Q (result[57]), .CK (CTS_n_tid0_142), .D (\tempResult[57] ));
DFF_X1 \result_reg[58]  (.Q (result[58]), .CK (CTS_n_tid0_142), .D (\tempResult[58] ));
DFF_X1 \result_reg[59]  (.Q (result[59]), .CK (CTS_n_tid0_142), .D (\tempResult[59] ));
DFF_X1 \result_reg[60]  (.Q (result[60]), .CK (CTS_n_tid0_142), .D (\tempResult[60] ));
DFF_X1 \result_reg[61]  (.Q (result[61]), .CK (CTS_n_tid0_142), .D (\tempResult[61] ));
DFF_X1 \result_reg[62]  (.Q (result[62]), .CK (CTS_n_tid0_142), .D (\tempResult[62] ));
DFF_X1 \result_reg[63]  (.Q (result[63]), .CK (CTS_n_tid0_142), .D (\tempResult[63] ));
CLKGATETST_X8 clk_gate_result_reg (.GCK (CTS_n_tid0_143), .CK (clk_CTS_1_PP_2), .E (n_168), .SE (1'b0 ));
BUF_X2 hfn_ipo_c23 (.Z (hfn_ipo_n23), .A (n_0_6));
CLKBUF_X3 hfn_ipo_c24 (.Z (hfn_ipo_n24), .A (n_0_6));
BUF_X2 hfn_ipo_c27 (.Z (hfn_ipo_n27), .A (n_0_38));
CLKBUF_X1 hfn_ipo_c28 (.Z (hfn_ipo_n28), .A (n_0_38));
BUF_X4 hfn_ipo_c31 (.Z (hfn_ipo_n31), .A (\shiftingAmount[1] ));
BUF_X4 hfn_ipo_c32 (.Z (hfn_ipo_n32), .A (\shiftingAmount[1] ));
CLKBUF_X1 hfn_ipo_c26 (.Z (hfn_ipo_n26), .A (n_0_20));
BUF_X4 hfn_ipo_c29 (.Z (hfn_ipo_n29), .A (\shiftingAmount[2] ));
CLKBUF_X1 hfn_ipo_c30 (.Z (hfn_ipo_n30), .A (\shiftingAmount[2] ));
BUF_X8 drc_ipo_c33 (.Z (drc_ipo_n33), .A (\shiftingAmount[3] ));
CLKBUF_X3 CTS_L4_c_tid0_41 (.Z (CTS_n_tid0_39), .A (CTS_n_tid0_105));
CLKBUF_X2 drc_ipo_c34 (.Z (drc_ipo_n34), .A (\shiftingAmount[5] ));
CLKBUF_X3 CTS_L4_c_tid0_42 (.Z (CTS_n_tid0_40), .A (CTS_n_tid0_105));
CLKBUF_X3 CTS_L3_c_tid1_43 (.Z (CTS_n_tid1_41), .A (CTS_n_tid1_133));
CLKBUF_X3 CTS_L3_c_tid1_44 (.Z (CTS_n_tid1_42), .A (CTS_n_tid1_133));
CLKBUF_X3 CTS_L3_c_tid0_111 (.Z (CTS_n_tid0_142), .A (CTS_n_tid0_143));
CLKBUF_X1 CLOCK_slh__c157 (.Z (CLOCK_slh_n239), .A (start));
CLKBUF_X2 CTS_L2_tid1__c2_tid1__c151 (.Z (n_tid1_233), .A (CTSclk_CTS_1_PP_2PP_0));

endmodule //Noaman_4_Booth

module Radix4 (clk, inputA, inputB, outResult, start);

output [63:0] outResult;
input clk;
input [31:0] inputA;
input [31:0] inputB;
input start;
wire CTS_n_tid1_3;
wire CLOCK_slh_n291;
wire CLOCK_slh_n286;
wire CLOCK_slh_n356;
wire CLOCK_slh_n246;
wire CLOCK_slh_n351;
wire CLOCK_slh_n346;
wire CLOCK_slh_n341;
wire CLOCK_slh_n256;
wire CLOCK_slh_n251;
wire CLOCK_slh_n261;
wire CLOCK_slh_n336;
wire CLOCK_slh_n331;
wire CLOCK_slh_n326;
wire CLOCK_slh_n321;
wire CLOCK_slh_n316;
wire CLOCK_slh_n311;
wire CLOCK_slh_n281;
wire CLOCK_slh_n306;
wire CLOCK_slh_n271;
wire CLOCK_slh_n301;
wire CLOCK_slh_n296;
wire CLOCK_slh_n266;
wire CLOCK_slh_n366;
wire CLOCK_slh_n361;
wire CLOCK_slh_n171;
wire CLOCK_slh_n276;
wire CLOCK_slh_n51;
wire CLOCK_slh_n201;
wire CLOCK_slh_n166;
wire CLOCK_slh_n196;
wire CLOCK_slh_n66;
wire CLOCK_slh_n61;
wire CLOCK_slh_n241;
wire CLOCK_slh_n96;
wire CLOCK_slh_n156;
wire CLOCK_slh_n231;
wire CLOCK_slh_n191;
wire CLOCK_slh_n226;
wire CLOCK_slh_n221;
wire CLOCK_slh_n141;
wire CLOCK_slh_n181;
wire CLOCK_slh_n86;
wire CLOCK_slh_n151;
wire CLOCK_slh_n216;
wire CLOCK_slh_n76;
wire CLOCK_slh_n71;
wire CLOCK_slh_n56;
wire CLOCK_slh_n176;
wire CLOCK_slh_n211;
wire CLOCK_slh_n81;
wire CLOCK_slh_n146;
wire CLOCK_slh_n111;
wire CLOCK_slh_n126;
wire CLOCK_slh_n131;
wire CLOCK_slh_n161;
wire CLOCK_slh_n186;
wire CLOCK_slh_n106;
wire CLOCK_slh_n91;
wire CLOCK_slh_n121;
wire CLOCK_slh_n101;
wire CLOCK_slh_n116;
wire CLOCK_slh_n236;
wire CLOCK_slh_n136;
wire CLOCK_slh_n206;
wire \result[63] ;
wire \result[62] ;
wire \result[61] ;
wire \result[60] ;
wire \result[59] ;
wire \result[58] ;
wire \result[57] ;
wire \result[56] ;
wire \result[55] ;
wire \result[54] ;
wire \result[53] ;
wire \result[52] ;
wire \result[51] ;
wire \result[50] ;
wire \result[49] ;
wire \result[48] ;
wire \result[47] ;
wire \result[46] ;
wire \result[45] ;
wire \result[44] ;
wire \result[43] ;
wire \result[42] ;
wire \result[41] ;
wire \result[40] ;
wire \result[39] ;
wire \result[38] ;
wire \result[37] ;
wire \result[36] ;
wire \result[35] ;
wire \result[34] ;
wire \result[33] ;
wire \result[32] ;
wire \result[31] ;
wire \result[30] ;
wire \result[29] ;
wire \result[28] ;
wire \result[27] ;
wire \result[26] ;
wire \result[25] ;
wire \result[24] ;
wire \result[23] ;
wire \result[22] ;
wire \result[21] ;
wire \result[20] ;
wire \result[19] ;
wire \result[18] ;
wire \result[17] ;
wire \result[16] ;
wire \result[15] ;
wire \result[14] ;
wire \result[13] ;
wire \result[12] ;
wire \result[11] ;
wire \result[10] ;
wire \result[9] ;
wire \result[8] ;
wire \result[7] ;
wire \result[6] ;
wire \result[5] ;
wire \result[4] ;
wire \result[3] ;
wire \result[2] ;
wire \result[1] ;
wire \result[0] ;
wire \B[31] ;
wire \B[30] ;
wire \B[29] ;
wire \B[28] ;
wire \B[27] ;
wire \B[26] ;
wire \B[25] ;
wire \B[24] ;
wire \B[23] ;
wire \B[22] ;
wire \B[21] ;
wire \B[20] ;
wire \B[19] ;
wire \B[18] ;
wire \B[17] ;
wire \B[16] ;
wire \B[15] ;
wire \B[14] ;
wire \B[13] ;
wire \B[12] ;
wire \B[11] ;
wire \B[10] ;
wire \B[9] ;
wire \B[8] ;
wire \B[7] ;
wire \B[6] ;
wire \B[5] ;
wire \B[4] ;
wire \B[3] ;
wire \B[2] ;
wire \B[1] ;
wire \B[0] ;
wire \A[31] ;
wire \A[30] ;
wire \A[29] ;
wire \A[28] ;
wire \A[27] ;
wire \A[26] ;
wire \A[25] ;
wire \A[24] ;
wire \A[23] ;
wire \A[22] ;
wire \A[21] ;
wire \A[20] ;
wire \A[19] ;
wire \A[18] ;
wire \A[17] ;
wire \A[16] ;
wire \A[15] ;
wire \A[14] ;
wire \A[13] ;
wire \A[12] ;
wire \A[11] ;
wire \A[10] ;
wire \A[9] ;
wire \A[8] ;
wire \A[7] ;
wire \A[6] ;
wire \A[5] ;
wire \A[4] ;
wire \A[3] ;
wire \A[2] ;
wire \A[1] ;
wire \A[0] ;
wire CTS_n_tid1_4;
wire CTS_n_tid1_5;
wire n_tid1_46;
wire CLOCK_slh__n367;
wire CLOCK_slh__n368;
wire CLOCK_slh__n371;
wire CLOCK_slh__n372;
wire CLOCK_slh__n375;
wire CLOCK_slh__n376;
wire CLOCK_slh__n379;
wire CLOCK_slh__n380;
wire CLOCK_slh__n383;
wire CLOCK_slh__n384;
wire CLOCK_slh__n387;
wire CLOCK_slh__n388;
wire CLOCK_slh__n391;
wire CLOCK_slh__n392;
wire CLOCK_slh__n395;
wire CLOCK_slh__n396;
wire CLOCK_slh__n399;
wire CLOCK_slh__n400;
wire CLOCK_slh__n403;
wire CLOCK_slh__n404;
wire CLOCK_slh__n407;
wire CLOCK_slh__n408;
wire CLOCK_slh__n411;
wire CLOCK_slh__n412;
wire CLOCK_slh__n415;
wire CLOCK_slh__n416;
wire CLOCK_slh__n419;
wire CLOCK_slh__n420;
wire CLOCK_slh__n423;
wire CLOCK_slh__n424;
wire CLOCK_slh__n427;
wire CLOCK_slh__n428;
wire CLOCK_slh__n431;
wire CLOCK_slh__n432;
wire CLOCK_slh__n435;
wire CLOCK_slh__n436;
wire CLOCK_slh__n439;
wire CLOCK_slh__n440;
wire CLOCK_slh__n443;
wire CLOCK_slh__n444;
wire CLOCK_slh__n447;
wire CLOCK_slh__n448;
wire CLOCK_slh__n451;
wire CLOCK_slh__n452;
wire CLOCK_slh__n455;
wire CLOCK_slh__n456;
wire CLOCK_slh__n459;
wire CLOCK_slh__n460;
wire CLOCK_slh__n463;
wire CLOCK_slh__n464;
wire CLOCK_slh__n467;
wire CLOCK_slh__n468;
wire CLOCK_slh__n471;
wire CLOCK_slh__n472;
wire CLOCK_slh__n475;
wire CLOCK_slh__n476;
wire CLOCK_slh__n479;
wire CLOCK_slh__n480;
wire CLOCK_slh__n483;
wire CLOCK_slh__n484;
wire CLOCK_slh__n487;
wire CLOCK_slh__n488;
wire CLOCK_slh__n491;
wire CLOCK_slh__n492;
wire CLOCK_slh__n495;
wire CLOCK_slh__n496;
wire CLOCK_slh__n499;
wire CLOCK_slh__n500;
wire CLOCK_slh__n503;
wire CLOCK_slh__n504;
wire CLOCK_slh__n507;
wire CLOCK_slh__n508;
wire CLOCK_slh__n511;
wire CLOCK_slh__n512;
wire CLOCK_slh__n515;
wire CLOCK_slh__n516;
wire CLOCK_slh__n519;
wire CLOCK_slh__n520;
wire CLOCK_slh__n523;
wire CLOCK_slh__n524;
wire CLOCK_slh__n527;
wire CLOCK_slh__n528;
wire CLOCK_slh__n531;
wire CLOCK_slh__n532;
wire CLOCK_slh__n535;
wire CLOCK_slh__n536;
wire CLOCK_slh__n539;
wire CLOCK_slh__n540;
wire CLOCK_slh__n543;
wire CLOCK_slh__n544;
wire CLOCK_slh__n547;
wire CLOCK_slh__n548;
wire CLOCK_slh__n551;
wire CLOCK_slh__n552;
wire CLOCK_slh__n555;
wire CLOCK_slh__n556;
wire CLOCK_slh__n559;
wire CLOCK_slh__n560;
wire CLOCK_slh__n563;
wire CLOCK_slh__n564;
wire CLOCK_slh__n567;
wire CLOCK_slh__n568;
wire CLOCK_slh__n571;
wire CLOCK_slh__n572;
wire CLOCK_slh__n575;
wire CLOCK_slh__n576;
wire CLOCK_slh__n579;
wire CLOCK_slh__n580;
wire CLOCK_slh__n583;
wire CLOCK_slh__n584;
wire CLOCK_slh__n587;
wire CLOCK_slh__n588;
wire CLOCK_slh__n591;
wire CLOCK_slh__n592;
wire CLOCK_slh__n595;
wire CLOCK_slh__n596;
wire CLOCK_slh__n599;
wire CLOCK_slh__n600;
wire CLOCK_slh__n603;
wire CLOCK_slh__n604;
wire CLOCK_slh__n607;
wire CLOCK_slh__n608;
wire CLOCK_slh__n611;
wire CLOCK_slh__n612;
wire CLOCK_slh__n615;
wire CLOCK_slh__n616;
wire CLOCK_slh__n619;
wire CLOCK_slh__n620;


DFF_X1 \A_reg[0]  (.Q (\A[0] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n61));
DFF_X1 \A_reg[1]  (.Q (\A[1] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n66));
DFF_X1 \A_reg[2]  (.Q (\A[2] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n196));
DFF_X1 \A_reg[3]  (.Q (\A[3] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n166));
DFF_X1 \A_reg[4]  (.Q (\A[4] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n201));
DFF_X1 \A_reg[5]  (.Q (\A[5] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n51));
DFF_X1 \A_reg[6]  (.Q (\A[6] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n276));
DFF_X1 \A_reg[7]  (.Q (\A[7] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n171));
DFF_X1 \A_reg[8]  (.Q (\A[8] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n361));
DFF_X1 \A_reg[9]  (.Q (\A[9] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n366));
DFF_X1 \A_reg[10]  (.Q (\A[10] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n266));
DFF_X1 \A_reg[11]  (.Q (\A[11] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n296));
DFF_X1 \A_reg[12]  (.Q (\A[12] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n301));
DFF_X1 \A_reg[13]  (.Q (\A[13] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n271));
DFF_X1 \A_reg[14]  (.Q (\A[14] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n306));
DFF_X1 \A_reg[15]  (.Q (\A[15] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n281));
DFF_X1 \A_reg[16]  (.Q (\A[16] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n311));
DFF_X1 \A_reg[17]  (.Q (\A[17] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n316));
DFF_X1 \A_reg[18]  (.Q (\A[18] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n321));
DFF_X1 \A_reg[19]  (.Q (\A[19] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n326));
DFF_X1 \A_reg[20]  (.Q (\A[20] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n331));
DFF_X1 \A_reg[21]  (.Q (\A[21] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n336));
DFF_X1 \A_reg[22]  (.Q (\A[22] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n261));
DFF_X1 \A_reg[23]  (.Q (\A[23] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n251));
DFF_X1 \A_reg[24]  (.Q (\A[24] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n256));
DFF_X1 \A_reg[25]  (.Q (\A[25] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n341));
DFF_X1 \A_reg[26]  (.Q (\A[26] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n346));
DFF_X1 \A_reg[27]  (.Q (\A[27] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n351));
DFF_X1 \A_reg[28]  (.Q (\A[28] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n246));
DFF_X1 \A_reg[29]  (.Q (\A[29] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n356));
DFF_X1 \A_reg[30]  (.Q (\A[30] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n286));
DFF_X1 \A_reg[31]  (.Q (\A[31] ), .CK (CTS_n_tid1_5), .D (CLOCK_slh_n291));
DFF_X1 \B_reg[0]  (.Q (\B[0] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n206));
DFF_X1 \B_reg[1]  (.Q (\B[1] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n136));
DFF_X1 \B_reg[2]  (.Q (\B[2] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n236));
DFF_X1 \B_reg[3]  (.Q (\B[3] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n116));
DFF_X1 \B_reg[4]  (.Q (\B[4] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n101));
DFF_X1 \B_reg[5]  (.Q (\B[5] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n121));
DFF_X1 \B_reg[6]  (.Q (\B[6] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n91));
DFF_X1 \B_reg[7]  (.Q (\B[7] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n106));
DFF_X1 \B_reg[8]  (.Q (\B[8] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n186));
DFF_X1 \B_reg[9]  (.Q (\B[9] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n161));
DFF_X1 \B_reg[10]  (.Q (\B[10] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n131));
DFF_X1 \B_reg[11]  (.Q (\B[11] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n126));
DFF_X1 \B_reg[12]  (.Q (\B[12] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n111));
DFF_X1 \B_reg[13]  (.Q (\B[13] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n146));
DFF_X1 \B_reg[14]  (.Q (\B[14] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n81));
DFF_X1 \B_reg[15]  (.Q (\B[15] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n211));
DFF_X1 \B_reg[16]  (.Q (\B[16] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n176));
DFF_X1 \B_reg[17]  (.Q (\B[17] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n56));
DFF_X1 \B_reg[18]  (.Q (\B[18] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n71));
DFF_X1 \B_reg[19]  (.Q (\B[19] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n76));
DFF_X1 \B_reg[20]  (.Q (\B[20] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n216));
DFF_X1 \B_reg[21]  (.Q (\B[21] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n151));
DFF_X1 \B_reg[22]  (.Q (\B[22] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n86));
DFF_X1 \B_reg[23]  (.Q (\B[23] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n181));
DFF_X1 \B_reg[24]  (.Q (\B[24] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n141));
DFF_X1 \B_reg[25]  (.Q (\B[25] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n221));
DFF_X1 \B_reg[26]  (.Q (\B[26] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n226));
DFF_X1 \B_reg[27]  (.Q (\B[27] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n191));
DFF_X1 \B_reg[28]  (.Q (\B[28] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n231));
DFF_X1 \B_reg[29]  (.Q (\B[29] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n156));
DFF_X1 \B_reg[30]  (.Q (\B[30] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n96));
DFF_X1 \B_reg[31]  (.Q (\B[31] ), .CK (CTS_n_tid1_3), .D (CLOCK_slh_n241));
DFF_X1 \outResult_reg[0]  (.Q (outResult[0]), .CK (CTS_n_tid1_3), .D (\result[0] ));
DFF_X1 \outResult_reg[1]  (.Q (outResult[1]), .CK (CTS_n_tid1_3), .D (\result[1] ));
DFF_X1 \outResult_reg[2]  (.Q (outResult[2]), .CK (CTS_n_tid1_3), .D (\result[2] ));
DFF_X1 \outResult_reg[3]  (.Q (outResult[3]), .CK (CTS_n_tid1_3), .D (\result[3] ));
DFF_X1 \outResult_reg[4]  (.Q (outResult[4]), .CK (CTS_n_tid1_3), .D (\result[4] ));
DFF_X1 \outResult_reg[5]  (.Q (outResult[5]), .CK (CTS_n_tid1_3), .D (\result[5] ));
DFF_X1 \outResult_reg[6]  (.Q (outResult[6]), .CK (CTS_n_tid1_3), .D (\result[6] ));
DFF_X1 \outResult_reg[7]  (.Q (outResult[7]), .CK (CTS_n_tid1_3), .D (\result[7] ));
DFF_X1 \outResult_reg[8]  (.Q (outResult[8]), .CK (CTS_n_tid1_3), .D (\result[8] ));
DFF_X1 \outResult_reg[9]  (.Q (outResult[9]), .CK (CTS_n_tid1_3), .D (\result[9] ));
DFF_X1 \outResult_reg[10]  (.Q (outResult[10]), .CK (CTS_n_tid1_3), .D (\result[10] ));
DFF_X1 \outResult_reg[11]  (.Q (outResult[11]), .CK (CTS_n_tid1_3), .D (\result[11] ));
DFF_X1 \outResult_reg[12]  (.Q (outResult[12]), .CK (CTS_n_tid1_3), .D (\result[12] ));
DFF_X1 \outResult_reg[13]  (.Q (outResult[13]), .CK (CTS_n_tid1_3), .D (\result[13] ));
DFF_X1 \outResult_reg[14]  (.Q (outResult[14]), .CK (CTS_n_tid1_4), .D (\result[14] ));
DFF_X1 \outResult_reg[15]  (.Q (outResult[15]), .CK (CTS_n_tid1_4), .D (\result[15] ));
DFF_X1 \outResult_reg[16]  (.Q (outResult[16]), .CK (CTS_n_tid1_4), .D (\result[16] ));
DFF_X1 \outResult_reg[17]  (.Q (outResult[17]), .CK (CTS_n_tid1_4), .D (\result[17] ));
DFF_X1 \outResult_reg[18]  (.Q (outResult[18]), .CK (CTS_n_tid1_4), .D (\result[18] ));
DFF_X1 \outResult_reg[19]  (.Q (outResult[19]), .CK (CTS_n_tid1_4), .D (\result[19] ));
DFF_X1 \outResult_reg[20]  (.Q (outResult[20]), .CK (CTS_n_tid1_5), .D (\result[20] ));
DFF_X1 \outResult_reg[21]  (.Q (outResult[21]), .CK (CTS_n_tid1_5), .D (\result[21] ));
DFF_X1 \outResult_reg[22]  (.Q (outResult[22]), .CK (CTS_n_tid1_5), .D (\result[22] ));
DFF_X1 \outResult_reg[23]  (.Q (outResult[23]), .CK (CTS_n_tid1_5), .D (\result[23] ));
DFF_X1 \outResult_reg[24]  (.Q (outResult[24]), .CK (CTS_n_tid1_5), .D (\result[24] ));
DFF_X1 \outResult_reg[25]  (.Q (outResult[25]), .CK (CTS_n_tid1_5), .D (\result[25] ));
DFF_X1 \outResult_reg[26]  (.Q (outResult[26]), .CK (CTS_n_tid1_5), .D (\result[26] ));
DFF_X1 \outResult_reg[27]  (.Q (outResult[27]), .CK (CTS_n_tid1_5), .D (\result[27] ));
DFF_X1 \outResult_reg[28]  (.Q (outResult[28]), .CK (CTS_n_tid1_5), .D (\result[28] ));
DFF_X1 \outResult_reg[29]  (.Q (outResult[29]), .CK (CTS_n_tid1_5), .D (\result[29] ));
DFF_X1 \outResult_reg[30]  (.Q (outResult[30]), .CK (CTS_n_tid1_5), .D (\result[30] ));
DFF_X1 \outResult_reg[31]  (.Q (outResult[31]), .CK (CTS_n_tid1_5), .D (\result[31] ));
DFF_X1 \outResult_reg[32]  (.Q (outResult[32]), .CK (CTS_n_tid1_5), .D (\result[32] ));
DFF_X1 \outResult_reg[33]  (.Q (outResult[33]), .CK (CTS_n_tid1_5), .D (\result[33] ));
DFF_X1 \outResult_reg[34]  (.Q (outResult[34]), .CK (CTS_n_tid1_4), .D (\result[34] ));
DFF_X1 \outResult_reg[35]  (.Q (outResult[35]), .CK (CTS_n_tid1_4), .D (\result[35] ));
DFF_X1 \outResult_reg[36]  (.Q (outResult[36]), .CK (CTS_n_tid1_4), .D (\result[36] ));
DFF_X1 \outResult_reg[37]  (.Q (outResult[37]), .CK (CTS_n_tid1_4), .D (\result[37] ));
DFF_X1 \outResult_reg[38]  (.Q (outResult[38]), .CK (CTS_n_tid1_4), .D (\result[38] ));
DFF_X1 \outResult_reg[39]  (.Q (outResult[39]), .CK (CTS_n_tid1_4), .D (\result[39] ));
DFF_X1 \outResult_reg[40]  (.Q (outResult[40]), .CK (CTS_n_tid1_4), .D (\result[40] ));
DFF_X1 \outResult_reg[41]  (.Q (outResult[41]), .CK (CTS_n_tid1_4), .D (\result[41] ));
DFF_X1 \outResult_reg[42]  (.Q (outResult[42]), .CK (CTS_n_tid1_3), .D (\result[42] ));
DFF_X1 \outResult_reg[43]  (.Q (outResult[43]), .CK (CTS_n_tid1_4), .D (\result[43] ));
DFF_X1 \outResult_reg[44]  (.Q (outResult[44]), .CK (CTS_n_tid1_4), .D (\result[44] ));
DFF_X1 \outResult_reg[45]  (.Q (outResult[45]), .CK (CTS_n_tid1_4), .D (\result[45] ));
DFF_X1 \outResult_reg[46]  (.Q (outResult[46]), .CK (CTS_n_tid1_4), .D (\result[46] ));
DFF_X1 \outResult_reg[47]  (.Q (outResult[47]), .CK (CTS_n_tid1_4), .D (\result[47] ));
DFF_X1 \outResult_reg[48]  (.Q (outResult[48]), .CK (CTS_n_tid1_5), .D (\result[48] ));
DFF_X1 \outResult_reg[49]  (.Q (outResult[49]), .CK (CTS_n_tid1_5), .D (\result[49] ));
DFF_X1 \outResult_reg[50]  (.Q (outResult[50]), .CK (CTS_n_tid1_5), .D (\result[50] ));
DFF_X1 \outResult_reg[51]  (.Q (outResult[51]), .CK (CTS_n_tid1_5), .D (\result[51] ));
DFF_X1 \outResult_reg[52]  (.Q (outResult[52]), .CK (CTS_n_tid1_5), .D (\result[52] ));
DFF_X1 \outResult_reg[53]  (.Q (outResult[53]), .CK (CTS_n_tid1_5), .D (\result[53] ));
DFF_X1 \outResult_reg[54]  (.Q (outResult[54]), .CK (CTS_n_tid1_5), .D (\result[54] ));
DFF_X1 \outResult_reg[55]  (.Q (outResult[55]), .CK (CTS_n_tid1_5), .D (\result[55] ));
DFF_X1 \outResult_reg[56]  (.Q (outResult[56]), .CK (CTS_n_tid1_5), .D (\result[56] ));
DFF_X1 \outResult_reg[57]  (.Q (outResult[57]), .CK (CTS_n_tid1_5), .D (\result[57] ));
DFF_X1 \outResult_reg[58]  (.Q (outResult[58]), .CK (CTS_n_tid1_5), .D (\result[58] ));
DFF_X1 \outResult_reg[59]  (.Q (outResult[59]), .CK (CTS_n_tid1_5), .D (\result[59] ));
DFF_X1 \outResult_reg[60]  (.Q (outResult[60]), .CK (CTS_n_tid1_5), .D (\result[60] ));
DFF_X1 \outResult_reg[61]  (.Q (outResult[61]), .CK (CTS_n_tid1_5), .D (\result[61] ));
DFF_X1 \outResult_reg[62]  (.Q (outResult[62]), .CK (CTS_n_tid1_5), .D (\result[62] ));
DFF_X1 \outResult_reg[63]  (.Q (outResult[63]), .CK (CTS_n_tid1_5), .D (\result[63] ));
Noaman_4_Booth mult (.result ({\result[63] , \result[62] , \result[61] , \result[60] , 
    \result[59] , \result[58] , \result[57] , \result[56] , \result[55] , \result[54] , 
    \result[53] , \result[52] , \result[51] , \result[50] , \result[49] , \result[48] , 
    \result[47] , \result[46] , \result[45] , \result[44] , \result[43] , \result[42] , 
    \result[41] , \result[40] , \result[39] , \result[38] , \result[37] , \result[36] , 
    \result[35] , \result[34] , \result[33] , \result[32] , \result[31] , \result[30] , 
    \result[29] , \result[28] , \result[27] , \result[26] , \result[25] , \result[24] , 
    \result[23] , \result[22] , \result[21] , \result[20] , \result[19] , \result[18] , 
    \result[17] , \result[16] , \result[15] , \result[14] , \result[13] , \result[12] , 
    \result[11] , \result[10] , \result[9] , \result[8] , \result[7] , \result[6] , 
    \result[5] , \result[4] , \result[3] , \result[2] , \result[1] , \result[0] })
    , .in1 ({\A[31] , \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , 
    \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] , \A[15] , 
    \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] , 
    \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] }), .in2 ({\B[31] , \B[30] , \B[29] , 
    \B[28] , \B[27] , \B[26] , \B[25] , \B[24] , \B[23] , \B[22] , \B[21] , \B[20] , 
    \B[19] , \B[18] , \B[17] , \B[16] , \B[15] , \B[14] , \B[13] , \B[12] , \B[11] , 
    \B[10] , \B[9] , \B[8] , \B[7] , \B[6] , \B[5] , \B[4] , \B[3] , \B[2] , \B[1] , 
    \B[0] }), .start (start), .clk_CTS_1_PP_2 (n_tid1_46), .CTSclk_CTS_1_PP_2PP_0 (n_tid1_46));
CLKBUF_X2 CTS_L2_c_tid1_2 (.Z (CTS_n_tid1_3), .A (n_tid1_46));
CLKBUF_X1 CTS_L2_c_tid1_3 (.Z (CTS_n_tid1_4), .A (n_tid1_46));
CLKBUF_X2 CTS_L2_c_tid1_4 (.Z (CTS_n_tid1_5), .A (n_tid1_46));
CLKBUF_X1 CLOCK_slh__c19 (.Z (CLOCK_slh__n487), .A (inputA[5]));
CLKBUF_X1 CLOCK_slh__c21 (.Z (CLOCK_slh__n371), .A (inputB[17]));
CLKBUF_X3 CTS_L1_tid1__c1_tid1__c15 (.Z (n_tid1_46), .A (clk));
CLKBUF_X1 CLOCK_slh__c23 (.Z (CLOCK_slh__n419), .A (inputA[0]));
CLKBUF_X1 CLOCK_slh__c25 (.Z (CLOCK_slh__n463), .A (inputA[1]));
CLKBUF_X1 CLOCK_slh__c27 (.Z (CLOCK_slh__n375), .A (inputB[18]));
CLKBUF_X1 CLOCK_slh__c29 (.Z (CLOCK_slh__n395), .A (inputB[19]));
CLKBUF_X1 CLOCK_slh__c31 (.Z (CLOCK_slh__n423), .A (inputB[14]));
CLKBUF_X1 CLOCK_slh__c33 (.Z (CLOCK_slh__n379), .A (inputB[22]));
CLKBUF_X1 CLOCK_slh__c35 (.Z (CLOCK_slh__n383), .A (inputB[6]));
CLKBUF_X1 CLOCK_slh__c37 (.Z (CLOCK_slh__n367), .A (inputB[30]));
CLKBUF_X1 CLOCK_slh__c39 (.Z (CLOCK_slh__n387), .A (inputB[4]));
CLKBUF_X1 CLOCK_slh__c41 (.Z (CLOCK_slh__n399), .A (inputB[7]));
CLKBUF_X1 CLOCK_slh__c43 (.Z (CLOCK_slh__n435), .A (inputB[12]));
CLKBUF_X1 CLOCK_slh__c45 (.Z (CLOCK_slh__n439), .A (inputB[3]));
CLKBUF_X1 CLOCK_slh__c47 (.Z (CLOCK_slh__n443), .A (inputB[5]));
CLKBUF_X1 CLOCK_slh__c49 (.Z (CLOCK_slh__n403), .A (inputB[11]));
CLKBUF_X1 CLOCK_slh__c51 (.Z (CLOCK_slh__n431), .A (inputB[10]));
CLKBUF_X1 CLOCK_slh__c53 (.Z (CLOCK_slh__n427), .A (inputB[1]));
CLKBUF_X1 CLOCK_slh__c55 (.Z (CLOCK_slh__n391), .A (inputB[24]));
CLKBUF_X1 CLOCK_slh__c57 (.Z (CLOCK_slh__n447), .A (inputB[13]));
CLKBUF_X1 CLOCK_slh__c59 (.Z (CLOCK_slh__n411), .A (inputB[21]));
CLKBUF_X1 CLOCK_slh__c61 (.Z (CLOCK_slh__n407), .A (inputB[29]));
CLKBUF_X1 CLOCK_slh__c63 (.Z (CLOCK_slh__n415), .A (inputB[9]));
CLKBUF_X1 CLOCK_slh__c65 (.Z (CLOCK_slh__n507), .A (inputA[3]));
CLKBUF_X1 CLOCK_slh__c67 (.Z (CLOCK_slh__n475), .A (inputA[7]));
CLKBUF_X1 CLOCK_slh__c69 (.Z (CLOCK_slh__n495), .A (inputB[16]));
CLKBUF_X1 CLOCK_slh__c71 (.Z (CLOCK_slh__n479), .A (inputB[23]));
CLKBUF_X1 CLOCK_slh__c73 (.Z (CLOCK_slh__n483), .A (inputB[8]));
CLKBUF_X1 CLOCK_slh__c75 (.Z (CLOCK_slh__n467), .A (inputB[27]));
CLKBUF_X1 CLOCK_slh__c77 (.Z (CLOCK_slh__n499), .A (inputA[2]));
CLKBUF_X1 CLOCK_slh__c79 (.Z (CLOCK_slh__n511), .A (inputA[4]));
CLKBUF_X1 CLOCK_slh__c81 (.Z (CLOCK_slh__n519), .A (inputB[0]));
CLKBUF_X1 CLOCK_slh__c83 (.Z (CLOCK_slh__n471), .A (inputB[15]));
CLKBUF_X1 CLOCK_slh__c85 (.Z (CLOCK_slh__n455), .A (inputB[20]));
CLKBUF_X1 CLOCK_slh__c87 (.Z (CLOCK_slh__n515), .A (inputB[25]));
CLKBUF_X1 CLOCK_slh__c89 (.Z (CLOCK_slh__n459), .A (inputB[26]));
CLKBUF_X1 CLOCK_slh__c91 (.Z (CLOCK_slh__n451), .A (inputB[28]));
CLKBUF_X1 CLOCK_slh__c93 (.Z (CLOCK_slh__n491), .A (inputB[2]));
CLKBUF_X1 CLOCK_slh__c95 (.Z (CLOCK_slh__n503), .A (inputB[31]));
CLKBUF_X1 CLOCK_slh__c97 (.Z (CLOCK_slh__n591), .A (inputA[28]));
CLKBUF_X1 CLOCK_slh__c99 (.Z (CLOCK_slh__n575), .A (inputA[23]));
CLKBUF_X1 CLOCK_slh__c101 (.Z (CLOCK_slh__n571), .A (inputA[24]));
CLKBUF_X1 CLOCK_slh__c103 (.Z (CLOCK_slh__n583), .A (inputA[22]));
CLKBUF_X1 CLOCK_slh__c105 (.Z (CLOCK_slh__n567), .A (inputA[10]));
CLKBUF_X1 CLOCK_slh__c107 (.Z (CLOCK_slh__n563), .A (inputA[13]));
CLKBUF_X1 CLOCK_slh__c109 (.Z (CLOCK_slh__n607), .A (inputA[6]));
CLKBUF_X1 CLOCK_slh__c111 (.Z (CLOCK_slh__n587), .A (inputA[15]));
CLKBUF_X1 CLOCK_slh__c113 (.Z (CLOCK_slh__n551), .A (inputA[30]));
CLKBUF_X1 CLOCK_slh__c115 (.Z (CLOCK_slh__n555), .A (inputA[31]));
CLKBUF_X1 CLOCK_slh__c117 (.Z (CLOCK_slh__n599), .A (inputA[11]));
CLKBUF_X1 CLOCK_slh__c119 (.Z (CLOCK_slh__n543), .A (inputA[12]));
CLKBUF_X1 CLOCK_slh__c121 (.Z (CLOCK_slh__n595), .A (inputA[14]));
CLKBUF_X1 CLOCK_slh__c123 (.Z (CLOCK_slh__n547), .A (inputA[16]));
CLKBUF_X1 CLOCK_slh__c125 (.Z (CLOCK_slh__n603), .A (inputA[17]));
CLKBUF_X1 CLOCK_slh__c127 (.Z (CLOCK_slh__n535), .A (inputA[18]));
CLKBUF_X1 CLOCK_slh__c129 (.Z (CLOCK_slh__n611), .A (inputA[19]));
CLKBUF_X1 CLOCK_slh__c131 (.Z (CLOCK_slh__n531), .A (inputA[20]));
CLKBUF_X1 CLOCK_slh__c133 (.Z (CLOCK_slh__n579), .A (inputA[21]));
CLKBUF_X1 CLOCK_slh__c135 (.Z (CLOCK_slh__n523), .A (inputA[25]));
CLKBUF_X1 CLOCK_slh__c137 (.Z (CLOCK_slh__n527), .A (inputA[26]));
CLKBUF_X1 CLOCK_slh__c139 (.Z (CLOCK_slh__n539), .A (inputA[27]));
CLKBUF_X1 CLOCK_slh__c141 (.Z (CLOCK_slh__n559), .A (inputA[29]));
CLKBUF_X1 CLOCK_slh__c143 (.Z (CLOCK_slh__n619), .A (inputA[8]));
CLKBUF_X1 CLOCK_slh__c145 (.Z (CLOCK_slh__n615), .A (inputA[9]));
CLKBUF_X1 CLOCK_slh__c147 (.Z (CLOCK_slh__n368), .A (CLOCK_slh__n367));
CLKBUF_X1 CLOCK_slh__c148 (.Z (CLOCK_slh_n96), .A (CLOCK_slh__n368));
CLKBUF_X1 CLOCK_slh__c151 (.Z (CLOCK_slh__n372), .A (CLOCK_slh__n371));
CLKBUF_X1 CLOCK_slh__c152 (.Z (CLOCK_slh_n56), .A (CLOCK_slh__n372));
CLKBUF_X1 CLOCK_slh__c155 (.Z (CLOCK_slh__n376), .A (CLOCK_slh__n375));
CLKBUF_X1 CLOCK_slh__c156 (.Z (CLOCK_slh_n71), .A (CLOCK_slh__n376));
CLKBUF_X1 CLOCK_slh__c159 (.Z (CLOCK_slh__n380), .A (CLOCK_slh__n379));
CLKBUF_X1 CLOCK_slh__c160 (.Z (CLOCK_slh_n86), .A (CLOCK_slh__n380));
CLKBUF_X1 CLOCK_slh__c163 (.Z (CLOCK_slh__n384), .A (CLOCK_slh__n383));
CLKBUF_X1 CLOCK_slh__c164 (.Z (CLOCK_slh_n91), .A (CLOCK_slh__n384));
CLKBUF_X1 CLOCK_slh__c167 (.Z (CLOCK_slh__n388), .A (CLOCK_slh__n387));
CLKBUF_X1 CLOCK_slh__c168 (.Z (CLOCK_slh_n101), .A (CLOCK_slh__n388));
CLKBUF_X1 CLOCK_slh__c171 (.Z (CLOCK_slh__n392), .A (CLOCK_slh__n391));
CLKBUF_X1 CLOCK_slh__c172 (.Z (CLOCK_slh_n141), .A (CLOCK_slh__n392));
CLKBUF_X1 CLOCK_slh__c175 (.Z (CLOCK_slh__n396), .A (CLOCK_slh__n395));
CLKBUF_X1 CLOCK_slh__c176 (.Z (CLOCK_slh_n76), .A (CLOCK_slh__n396));
CLKBUF_X1 CLOCK_slh__c179 (.Z (CLOCK_slh__n400), .A (CLOCK_slh__n399));
CLKBUF_X1 CLOCK_slh__c180 (.Z (CLOCK_slh_n106), .A (CLOCK_slh__n400));
CLKBUF_X1 CLOCK_slh__c183 (.Z (CLOCK_slh__n404), .A (CLOCK_slh__n403));
CLKBUF_X1 CLOCK_slh__c184 (.Z (CLOCK_slh_n126), .A (CLOCK_slh__n404));
CLKBUF_X1 CLOCK_slh__c187 (.Z (CLOCK_slh__n408), .A (CLOCK_slh__n407));
CLKBUF_X1 CLOCK_slh__c188 (.Z (CLOCK_slh_n156), .A (CLOCK_slh__n408));
CLKBUF_X1 CLOCK_slh__c191 (.Z (CLOCK_slh__n412), .A (CLOCK_slh__n411));
CLKBUF_X1 CLOCK_slh__c192 (.Z (CLOCK_slh_n151), .A (CLOCK_slh__n412));
CLKBUF_X1 CLOCK_slh__c195 (.Z (CLOCK_slh__n416), .A (CLOCK_slh__n415));
CLKBUF_X1 CLOCK_slh__c196 (.Z (CLOCK_slh_n161), .A (CLOCK_slh__n416));
CLKBUF_X1 CLOCK_slh__c199 (.Z (CLOCK_slh__n420), .A (CLOCK_slh__n419));
CLKBUF_X1 CLOCK_slh__c200 (.Z (CLOCK_slh_n61), .A (CLOCK_slh__n420));
CLKBUF_X1 CLOCK_slh__c203 (.Z (CLOCK_slh__n424), .A (CLOCK_slh__n423));
CLKBUF_X1 CLOCK_slh__c204 (.Z (CLOCK_slh_n81), .A (CLOCK_slh__n424));
CLKBUF_X1 CLOCK_slh__c207 (.Z (CLOCK_slh__n428), .A (CLOCK_slh__n427));
CLKBUF_X1 CLOCK_slh__c208 (.Z (CLOCK_slh_n136), .A (CLOCK_slh__n428));
CLKBUF_X1 CLOCK_slh__c211 (.Z (CLOCK_slh__n432), .A (CLOCK_slh__n431));
CLKBUF_X1 CLOCK_slh__c212 (.Z (CLOCK_slh_n131), .A (CLOCK_slh__n432));
CLKBUF_X1 CLOCK_slh__c215 (.Z (CLOCK_slh__n436), .A (CLOCK_slh__n435));
CLKBUF_X1 CLOCK_slh__c216 (.Z (CLOCK_slh_n111), .A (CLOCK_slh__n436));
CLKBUF_X1 CLOCK_slh__c219 (.Z (CLOCK_slh__n440), .A (CLOCK_slh__n439));
CLKBUF_X1 CLOCK_slh__c220 (.Z (CLOCK_slh_n116), .A (CLOCK_slh__n440));
CLKBUF_X1 CLOCK_slh__c223 (.Z (CLOCK_slh__n444), .A (CLOCK_slh__n443));
CLKBUF_X1 CLOCK_slh__c224 (.Z (CLOCK_slh_n121), .A (CLOCK_slh__n444));
CLKBUF_X1 CLOCK_slh__c227 (.Z (CLOCK_slh__n448), .A (CLOCK_slh__n447));
CLKBUF_X1 CLOCK_slh__c228 (.Z (CLOCK_slh_n146), .A (CLOCK_slh__n448));
CLKBUF_X1 CLOCK_slh__c231 (.Z (CLOCK_slh__n452), .A (CLOCK_slh__n451));
CLKBUF_X1 CLOCK_slh__c232 (.Z (CLOCK_slh_n231), .A (CLOCK_slh__n452));
CLKBUF_X1 CLOCK_slh__c235 (.Z (CLOCK_slh__n456), .A (CLOCK_slh__n455));
CLKBUF_X1 CLOCK_slh__c236 (.Z (CLOCK_slh_n216), .A (CLOCK_slh__n456));
CLKBUF_X1 CLOCK_slh__c239 (.Z (CLOCK_slh__n460), .A (CLOCK_slh__n459));
CLKBUF_X1 CLOCK_slh__c240 (.Z (CLOCK_slh_n226), .A (CLOCK_slh__n460));
CLKBUF_X1 CLOCK_slh__c243 (.Z (CLOCK_slh__n464), .A (CLOCK_slh__n463));
CLKBUF_X1 CLOCK_slh__c244 (.Z (CLOCK_slh_n66), .A (CLOCK_slh__n464));
CLKBUF_X1 CLOCK_slh__c247 (.Z (CLOCK_slh__n468), .A (CLOCK_slh__n467));
CLKBUF_X1 CLOCK_slh__c248 (.Z (CLOCK_slh_n191), .A (CLOCK_slh__n468));
CLKBUF_X1 CLOCK_slh__c251 (.Z (CLOCK_slh__n472), .A (CLOCK_slh__n471));
CLKBUF_X1 CLOCK_slh__c252 (.Z (CLOCK_slh_n211), .A (CLOCK_slh__n472));
CLKBUF_X1 CLOCK_slh__c255 (.Z (CLOCK_slh__n476), .A (CLOCK_slh__n475));
CLKBUF_X1 CLOCK_slh__c256 (.Z (CLOCK_slh_n171), .A (CLOCK_slh__n476));
CLKBUF_X1 CLOCK_slh__c259 (.Z (CLOCK_slh__n480), .A (CLOCK_slh__n479));
CLKBUF_X1 CLOCK_slh__c260 (.Z (CLOCK_slh_n181), .A (CLOCK_slh__n480));
CLKBUF_X1 CLOCK_slh__c263 (.Z (CLOCK_slh__n484), .A (CLOCK_slh__n483));
CLKBUF_X1 CLOCK_slh__c264 (.Z (CLOCK_slh_n186), .A (CLOCK_slh__n484));
CLKBUF_X1 CLOCK_slh__c267 (.Z (CLOCK_slh__n488), .A (CLOCK_slh__n487));
CLKBUF_X1 CLOCK_slh__c268 (.Z (CLOCK_slh_n51), .A (CLOCK_slh__n488));
CLKBUF_X1 CLOCK_slh__c271 (.Z (CLOCK_slh__n492), .A (CLOCK_slh__n491));
CLKBUF_X1 CLOCK_slh__c272 (.Z (CLOCK_slh_n236), .A (CLOCK_slh__n492));
CLKBUF_X1 CLOCK_slh__c275 (.Z (CLOCK_slh__n496), .A (CLOCK_slh__n495));
CLKBUF_X1 CLOCK_slh__c276 (.Z (CLOCK_slh_n176), .A (CLOCK_slh__n496));
CLKBUF_X1 CLOCK_slh__c279 (.Z (CLOCK_slh__n500), .A (CLOCK_slh__n499));
CLKBUF_X1 CLOCK_slh__c280 (.Z (CLOCK_slh_n196), .A (CLOCK_slh__n500));
CLKBUF_X1 CLOCK_slh__c283 (.Z (CLOCK_slh__n504), .A (CLOCK_slh__n503));
CLKBUF_X1 CLOCK_slh__c284 (.Z (CLOCK_slh_n241), .A (CLOCK_slh__n504));
CLKBUF_X1 CLOCK_slh__c287 (.Z (CLOCK_slh__n508), .A (CLOCK_slh__n507));
CLKBUF_X1 CLOCK_slh__c288 (.Z (CLOCK_slh_n166), .A (CLOCK_slh__n508));
CLKBUF_X1 CLOCK_slh__c291 (.Z (CLOCK_slh__n512), .A (CLOCK_slh__n511));
CLKBUF_X1 CLOCK_slh__c292 (.Z (CLOCK_slh_n201), .A (CLOCK_slh__n512));
CLKBUF_X1 CLOCK_slh__c295 (.Z (CLOCK_slh__n516), .A (CLOCK_slh__n515));
CLKBUF_X1 CLOCK_slh__c296 (.Z (CLOCK_slh_n221), .A (CLOCK_slh__n516));
CLKBUF_X1 CLOCK_slh__c299 (.Z (CLOCK_slh__n520), .A (CLOCK_slh__n519));
CLKBUF_X1 CLOCK_slh__c300 (.Z (CLOCK_slh_n206), .A (CLOCK_slh__n520));
CLKBUF_X1 CLOCK_slh__c303 (.Z (CLOCK_slh__n524), .A (CLOCK_slh__n523));
CLKBUF_X1 CLOCK_slh__c304 (.Z (CLOCK_slh_n341), .A (CLOCK_slh__n524));
CLKBUF_X1 CLOCK_slh__c307 (.Z (CLOCK_slh__n528), .A (CLOCK_slh__n527));
CLKBUF_X1 CLOCK_slh__c308 (.Z (CLOCK_slh_n346), .A (CLOCK_slh__n528));
CLKBUF_X1 CLOCK_slh__c311 (.Z (CLOCK_slh__n532), .A (CLOCK_slh__n531));
CLKBUF_X1 CLOCK_slh__c312 (.Z (CLOCK_slh_n331), .A (CLOCK_slh__n532));
CLKBUF_X1 CLOCK_slh__c315 (.Z (CLOCK_slh__n536), .A (CLOCK_slh__n535));
CLKBUF_X1 CLOCK_slh__c316 (.Z (CLOCK_slh_n321), .A (CLOCK_slh__n536));
CLKBUF_X1 CLOCK_slh__c319 (.Z (CLOCK_slh__n540), .A (CLOCK_slh__n539));
CLKBUF_X1 CLOCK_slh__c320 (.Z (CLOCK_slh_n351), .A (CLOCK_slh__n540));
CLKBUF_X1 CLOCK_slh__c323 (.Z (CLOCK_slh__n544), .A (CLOCK_slh__n543));
CLKBUF_X1 CLOCK_slh__c324 (.Z (CLOCK_slh_n301), .A (CLOCK_slh__n544));
CLKBUF_X1 CLOCK_slh__c327 (.Z (CLOCK_slh__n548), .A (CLOCK_slh__n547));
CLKBUF_X1 CLOCK_slh__c328 (.Z (CLOCK_slh_n311), .A (CLOCK_slh__n548));
CLKBUF_X1 CLOCK_slh__c331 (.Z (CLOCK_slh__n552), .A (CLOCK_slh__n551));
CLKBUF_X1 CLOCK_slh__c332 (.Z (CLOCK_slh_n286), .A (CLOCK_slh__n552));
CLKBUF_X1 CLOCK_slh__c335 (.Z (CLOCK_slh__n556), .A (CLOCK_slh__n555));
CLKBUF_X1 CLOCK_slh__c336 (.Z (CLOCK_slh_n291), .A (CLOCK_slh__n556));
CLKBUF_X1 CLOCK_slh__c339 (.Z (CLOCK_slh__n560), .A (CLOCK_slh__n559));
CLKBUF_X1 CLOCK_slh__c340 (.Z (CLOCK_slh_n356), .A (CLOCK_slh__n560));
CLKBUF_X1 CLOCK_slh__c343 (.Z (CLOCK_slh__n564), .A (CLOCK_slh__n563));
CLKBUF_X1 CLOCK_slh__c344 (.Z (CLOCK_slh_n271), .A (CLOCK_slh__n564));
CLKBUF_X1 CLOCK_slh__c347 (.Z (CLOCK_slh__n568), .A (CLOCK_slh__n567));
CLKBUF_X1 CLOCK_slh__c348 (.Z (CLOCK_slh_n266), .A (CLOCK_slh__n568));
CLKBUF_X1 CLOCK_slh__c351 (.Z (CLOCK_slh__n572), .A (CLOCK_slh__n571));
CLKBUF_X1 CLOCK_slh__c352 (.Z (CLOCK_slh_n256), .A (CLOCK_slh__n572));
CLKBUF_X1 CLOCK_slh__c355 (.Z (CLOCK_slh__n576), .A (CLOCK_slh__n575));
CLKBUF_X1 CLOCK_slh__c356 (.Z (CLOCK_slh_n251), .A (CLOCK_slh__n576));
CLKBUF_X1 CLOCK_slh__c359 (.Z (CLOCK_slh__n580), .A (CLOCK_slh__n579));
CLKBUF_X1 CLOCK_slh__c360 (.Z (CLOCK_slh_n336), .A (CLOCK_slh__n580));
CLKBUF_X1 CLOCK_slh__c363 (.Z (CLOCK_slh__n584), .A (CLOCK_slh__n583));
CLKBUF_X1 CLOCK_slh__c364 (.Z (CLOCK_slh_n261), .A (CLOCK_slh__n584));
CLKBUF_X1 CLOCK_slh__c367 (.Z (CLOCK_slh__n588), .A (CLOCK_slh__n587));
CLKBUF_X1 CLOCK_slh__c368 (.Z (CLOCK_slh_n281), .A (CLOCK_slh__n588));
CLKBUF_X1 CLOCK_slh__c371 (.Z (CLOCK_slh__n592), .A (CLOCK_slh__n591));
CLKBUF_X1 CLOCK_slh__c372 (.Z (CLOCK_slh_n246), .A (CLOCK_slh__n592));
CLKBUF_X1 CLOCK_slh__c375 (.Z (CLOCK_slh__n596), .A (CLOCK_slh__n595));
CLKBUF_X1 CLOCK_slh__c376 (.Z (CLOCK_slh_n306), .A (CLOCK_slh__n596));
CLKBUF_X1 CLOCK_slh__c379 (.Z (CLOCK_slh__n600), .A (CLOCK_slh__n599));
CLKBUF_X1 CLOCK_slh__c380 (.Z (CLOCK_slh_n296), .A (CLOCK_slh__n600));
CLKBUF_X1 CLOCK_slh__c383 (.Z (CLOCK_slh__n604), .A (CLOCK_slh__n603));
CLKBUF_X1 CLOCK_slh__c384 (.Z (CLOCK_slh_n316), .A (CLOCK_slh__n604));
CLKBUF_X1 CLOCK_slh__c387 (.Z (CLOCK_slh__n608), .A (CLOCK_slh__n607));
CLKBUF_X1 CLOCK_slh__c388 (.Z (CLOCK_slh_n276), .A (CLOCK_slh__n608));
CLKBUF_X1 CLOCK_slh__c391 (.Z (CLOCK_slh__n612), .A (CLOCK_slh__n611));
CLKBUF_X1 CLOCK_slh__c392 (.Z (CLOCK_slh_n326), .A (CLOCK_slh__n612));
CLKBUF_X1 CLOCK_slh__c395 (.Z (CLOCK_slh__n616), .A (CLOCK_slh__n615));
CLKBUF_X1 CLOCK_slh__c396 (.Z (CLOCK_slh_n366), .A (CLOCK_slh__n616));
CLKBUF_X1 CLOCK_slh__c399 (.Z (CLOCK_slh__n620), .A (CLOCK_slh__n619));
CLKBUF_X1 CLOCK_slh__c400 (.Z (CLOCK_slh_n361), .A (CLOCK_slh__n620));

endmodule //Radix4


