
// 	Wed Jan  4 04:22:53 2023
//	vlsi
//	localhost.localdomain

module buffer__parameterized0 (clk_CTS_1_PP_0, clk, rst, en, D, Q);

output [0:0] Q;
input [0:0] D;
input clk;
input en;
input rst;
input clk_CTS_1_PP_0;
wire n_0_0;
wire n_0_1;
wire n_0;


INV_X1 i_0_2 (.ZN (n_0_1), .A (D[0]));
NOR2_X1 i_0_1 (.ZN (n_0_0), .A1 (Q[0]), .A2 (en));
AOI211_X1 i_0_0 (.ZN (n_0), .A (rst), .B (n_0_0), .C1 (n_0_1), .C2 (en));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (clk_CTS_1_PP_0), .D (n_0));

endmodule //buffer__parameterized0

module buffer__parameterized0__0_52 (clk_CTS_1_PP_0, clk_CTS_1_PP_8, clk, rst, en, 
    D, Q);

output [0:0] Q;
output clk_CTS_1_PP_0;
input [0:0] D;
input clk;
input en;
input rst;
input clk_CTS_1_PP_8;
wire n_0_0;
wire n_0_1;
wire n_0;


INV_X1 i_0_2 (.ZN (n_0_1), .A (D[0]));
NOR2_X1 i_0_1 (.ZN (n_0_0), .A1 (Q[0]), .A2 (en));
AOI211_X1 i_0_0 (.ZN (n_0), .A (rst), .B (n_0_0), .C1 (n_0_1), .C2 (en));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (clk_CTS_1_PP_0), .D (n_0));
CLKBUF_X3 CTS_L1_c_tid1_2 (.Z (clk_CTS_1_PP_0), .A (clk_CTS_1_PP_8));

endmodule //buffer__parameterized0__0_52

module buffer (clk_CTS_1_PP_3, clk, rst, en, D, Q);

output [31:0] Q;
input [31:0] D;
input clk;
input en;
input rst;
input clk_CTS_1_PP_3;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_tid1_46;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (D[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (D[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (D[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (D[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (D[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (D[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (D[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (D[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (D[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (D[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (D[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (D[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (D[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (D[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (D[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (D[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (D[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (D[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (D[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (D[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (D[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (D[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (D[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (D[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (D[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (D[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (D[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (D[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (D[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (D[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (D[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (D[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (rst));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (rst));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (n_0), .D (n_2));
DFF_X1 \Q_reg[1]  (.Q (Q[1]), .CK (n_0), .D (n_3));
DFF_X1 \Q_reg[2]  (.Q (Q[2]), .CK (n_0), .D (n_4));
DFF_X1 \Q_reg[3]  (.Q (Q[3]), .CK (n_0), .D (n_5));
DFF_X1 \Q_reg[4]  (.Q (Q[4]), .CK (n_0), .D (n_6));
DFF_X1 \Q_reg[5]  (.Q (Q[5]), .CK (n_0), .D (n_7));
DFF_X1 \Q_reg[6]  (.Q (Q[6]), .CK (n_0), .D (n_8));
DFF_X1 \Q_reg[7]  (.Q (Q[7]), .CK (n_0), .D (n_9));
DFF_X1 \Q_reg[8]  (.Q (Q[8]), .CK (n_0), .D (n_10));
DFF_X1 \Q_reg[9]  (.Q (Q[9]), .CK (n_0), .D (n_11));
DFF_X1 \Q_reg[10]  (.Q (Q[10]), .CK (n_0), .D (n_12));
DFF_X1 \Q_reg[11]  (.Q (Q[11]), .CK (n_0), .D (n_13));
DFF_X1 \Q_reg[12]  (.Q (Q[12]), .CK (n_0), .D (n_14));
DFF_X1 \Q_reg[13]  (.Q (Q[13]), .CK (n_0), .D (n_15));
DFF_X1 \Q_reg[14]  (.Q (Q[14]), .CK (n_0), .D (n_16));
DFF_X1 \Q_reg[15]  (.Q (Q[15]), .CK (n_0), .D (n_17));
DFF_X1 \Q_reg[16]  (.Q (Q[16]), .CK (n_0), .D (n_18));
DFF_X1 \Q_reg[17]  (.Q (Q[17]), .CK (n_0), .D (n_19));
DFF_X1 \Q_reg[18]  (.Q (Q[18]), .CK (n_0), .D (n_20));
DFF_X1 \Q_reg[19]  (.Q (Q[19]), .CK (n_0), .D (n_21));
DFF_X1 \Q_reg[20]  (.Q (Q[20]), .CK (n_0), .D (n_22));
DFF_X1 \Q_reg[21]  (.Q (Q[21]), .CK (n_0), .D (n_23));
DFF_X1 \Q_reg[22]  (.Q (Q[22]), .CK (n_0), .D (n_24));
DFF_X1 \Q_reg[23]  (.Q (Q[23]), .CK (n_0), .D (n_25));
DFF_X1 \Q_reg[24]  (.Q (Q[24]), .CK (n_0), .D (n_26));
DFF_X1 \Q_reg[25]  (.Q (Q[25]), .CK (n_0), .D (n_27));
DFF_X1 \Q_reg[26]  (.Q (Q[26]), .CK (n_0), .D (n_28));
DFF_X1 \Q_reg[27]  (.Q (Q[27]), .CK (n_0), .D (n_29));
DFF_X1 \Q_reg[28]  (.Q (Q[28]), .CK (n_0), .D (n_30));
DFF_X1 \Q_reg[29]  (.Q (Q[29]), .CK (n_0), .D (n_31));
DFF_X1 \Q_reg[30]  (.Q (Q[30]), .CK (n_0), .D (n_32));
DFF_X1 \Q_reg[31]  (.Q (Q[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_Q_reg (.GCK (n_0), .CK (n_tid1_46), .E (n_1), .SE (1'b0 ));
CLKBUF_X1 CTS_L1_tid1__c1_tid1__c7 (.Z (n_tid1_46), .A (clk_CTS_1_PP_3));

endmodule //buffer

module datapath__0_43 (mant_A, p_0);

output [31:0] p_0;
input [23:0] mant_A;
wire n_21;
wire n_0;
wire n_20;
wire n_19;
wire n_18;
wire n_1;
wire n_17;
wire n_16;
wire n_2;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_3;
wire n_6;
wire n_4;
wire n_5;
wire n_23;
wire n_22;


INV_X1 i_47 (.ZN (n_23), .A (mant_A[15]));
INV_X1 i_46 (.ZN (n_22), .A (mant_A[11]));
OR3_X1 i_45 (.ZN (n_21), .A1 (mant_A[2]), .A2 (mant_A[1]), .A3 (mant_A[0]));
OR2_X1 i_44 (.ZN (n_20), .A1 (n_21), .A2 (mant_A[3]));
OR2_X1 i_43 (.ZN (n_19), .A1 (n_20), .A2 (mant_A[4]));
OR3_X1 i_42 (.ZN (n_18), .A1 (n_19), .A2 (mant_A[5]), .A3 (mant_A[6]));
OR2_X1 i_41 (.ZN (n_17), .A1 (n_18), .A2 (mant_A[7]));
OR3_X1 i_40 (.ZN (n_16), .A1 (n_17), .A2 (mant_A[8]), .A3 (mant_A[9]));
NOR2_X1 i_39 (.ZN (n_15), .A1 (n_16), .A2 (mant_A[10]));
NAND2_X1 i_38 (.ZN (n_14), .A1 (n_15), .A2 (n_22));
OR2_X1 i_37 (.ZN (n_13), .A1 (n_14), .A2 (mant_A[12]));
NOR2_X1 i_36 (.ZN (n_12), .A1 (n_13), .A2 (mant_A[13]));
NOR3_X1 i_35 (.ZN (n_11), .A1 (n_13), .A2 (mant_A[13]), .A3 (mant_A[14]));
NAND2_X1 i_34 (.ZN (n_10), .A1 (n_11), .A2 (n_23));
OR2_X1 i_33 (.ZN (n_9), .A1 (n_10), .A2 (mant_A[16]));
OR2_X1 i_32 (.ZN (n_8), .A1 (n_9), .A2 (mant_A[17]));
OR3_X1 i_31 (.ZN (n_7), .A1 (n_8), .A2 (mant_A[18]), .A3 (mant_A[19]));
OR3_X1 i_30 (.ZN (n_6), .A1 (n_7), .A2 (mant_A[20]), .A3 (mant_A[21]));
OR3_X1 i_29 (.ZN (p_0[31]), .A1 (n_6), .A2 (mant_A[22]), .A3 (mant_A[23]));
OAI21_X1 i_28 (.ZN (n_5), .A (mant_A[23]), .B1 (n_6), .B2 (mant_A[22]));
AND2_X1 i_27 (.ZN (p_0[23]), .A1 (p_0[31]), .A2 (n_5));
XOR2_X1 i_26 (.Z (p_0[22]), .A (mant_A[22]), .B (n_6));
OAI21_X1 i_25 (.ZN (n_4), .A (mant_A[21]), .B1 (n_7), .B2 (mant_A[20]));
AND2_X1 i_24 (.ZN (p_0[21]), .A1 (n_6), .A2 (n_4));
XOR2_X1 i_23 (.Z (p_0[20]), .A (mant_A[20]), .B (n_7));
OAI21_X1 i_22 (.ZN (n_3), .A (mant_A[19]), .B1 (n_8), .B2 (mant_A[18]));
AND2_X1 i_21 (.ZN (p_0[19]), .A1 (n_7), .A2 (n_3));
XOR2_X1 i_20 (.Z (p_0[18]), .A (mant_A[18]), .B (n_8));
XOR2_X1 i_19 (.Z (p_0[17]), .A (mant_A[17]), .B (n_9));
XOR2_X1 i_18 (.Z (p_0[16]), .A (mant_A[16]), .B (n_10));
XNOR2_X1 i_17 (.ZN (p_0[15]), .A (mant_A[15]), .B (n_11));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (mant_A[14]), .B (n_12));
XOR2_X1 i_15 (.Z (p_0[13]), .A (mant_A[13]), .B (n_13));
XOR2_X1 i_14 (.Z (p_0[12]), .A (mant_A[12]), .B (n_14));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (mant_A[11]), .B (n_15));
XOR2_X1 i_12 (.Z (p_0[10]), .A (mant_A[10]), .B (n_16));
OAI21_X1 i_11 (.ZN (n_2), .A (mant_A[9]), .B1 (n_17), .B2 (mant_A[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_16), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (mant_A[8]), .B (n_17));
XOR2_X1 i_8 (.Z (p_0[7]), .A (mant_A[7]), .B (n_18));
OAI21_X1 i_7 (.ZN (n_1), .A (mant_A[6]), .B1 (n_19), .B2 (mant_A[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_18), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (mant_A[5]), .B (n_19));
XOR2_X1 i_4 (.Z (p_0[4]), .A (mant_A[4]), .B (n_20));
XOR2_X1 i_3 (.Z (p_0[3]), .A (mant_A[3]), .B (n_21));
OAI21_X1 i_2 (.ZN (n_0), .A (mant_A[2]), .B1 (mant_A[1]), .B2 (mant_A[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_21), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (mant_A[1]), .B (mant_A[0]));

endmodule //datapath__0_43

module datapath__0_38 (p_0, p_1);

output [10:0] p_1;
input [21:0] p_0;
wire drc_ipo_n10;
wire drc_ipo_n12;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire spc__n13;


HA_X1 i_4 (.CO (n_3), .S (spc__n13), .A (p_0[4]), .B (n_2));
HA_X1 i_3 (.CO (n_2), .S (p_1[3]), .A (p_0[3]), .B (n_1));
HA_X1 i_2 (.CO (n_1), .S (drc_ipo_n10), .A (p_0[2]), .B (n_0));
HA_X1 i_1 (.CO (n_0), .S (drc_ipo_n12), .A (p_0[1]), .B (p_0[11]));
INV_X1 i_0 (.ZN (p_1[0]), .A (p_0[11]));
CLKBUF_X1 drc_ipo_c5 (.Z (p_1[2]), .A (drc_ipo_n10));
CLKBUF_X1 drc_ipo_c6 (.Z (p_1[1]), .A (drc_ipo_n12));
CLKBUF_X1 spc__c7 (.Z (p_1[4]), .A (spc__n13));

endmodule //datapath__0_38

module datapath__0_25 (p_0, exp_Sum, p_1);

output p_0;
input [7:0] exp_Sum;
input [21:0] p_1;
wire n_6;
wire n_4;
wire n_18;
wire n_5;
wire n_7;
wire n_0;
wire n_8;
wire n_11;
wire n_1;
wire n_12;
wire n_15;
wire n_2;
wire n_16;
wire n_3;
wire n_17;
wire n_14;
wire n_13;
wire n_10;
wire n_9;


INV_X1 i_14 (.ZN (n_17), .A (exp_Sum[4]));
INV_X1 i_13 (.ZN (n_14), .A (exp_Sum[3]));
INV_X1 i_12 (.ZN (n_13), .A (exp_Sum[2]));
INV_X1 i_11 (.ZN (n_10), .A (exp_Sum[1]));
INV_X1 i_10 (.ZN (n_9), .A (exp_Sum[0]));
NOR3_X1 i_9 (.ZN (p_0), .A1 (exp_Sum[7]), .A2 (exp_Sum[6]), .A3 (n_3));
NAND2_X1 i_8 (.ZN (n_6), .A1 (n_9), .A2 (p_1[11]));
NAND2_X1 i_7 (.ZN (n_5), .A1 (n_10), .A2 (p_1[1]));
OAI21_X1 i_6 (.ZN (n_4), .A (n_5), .B1 (n_10), .B2 (p_1[1]));
NAND2_X1 i_5 (.ZN (n_8), .A1 (n_13), .A2 (p_1[2]));
OAI21_X1 i_4 (.ZN (n_7), .A (n_8), .B1 (n_13), .B2 (p_1[2]));
NAND2_X1 i_3 (.ZN (n_12), .A1 (n_14), .A2 (p_1[3]));
OAI21_X1 i_2 (.ZN (n_11), .A (n_12), .B1 (n_14), .B2 (p_1[3]));
NAND2_X1 i_1 (.ZN (n_16), .A1 (n_17), .A2 (p_1[4]));
OAI21_X1 i_0 (.ZN (n_15), .A (n_16), .B1 (n_17), .B2 (p_1[4]));
FA_X1 i_22 (.CO (n_3), .A (exp_Sum[5]), .B (n_16), .CI (n_2));
FA_X1 i_21 (.CO (n_2), .A (n_12), .B (n_15), .CI (n_1));
FA_X1 i_20 (.CO (n_1), .A (n_8), .B (n_11), .CI (n_0));
FA_X1 i_19 (.CO (n_0), .A (n_5), .B (n_7), .CI (n_18));
HA_X1 i_18 (.CO (n_18), .A (n_6), .B (n_4));

endmodule //datapath__0_25

module count_leading_zeros (valueIn, result);

output [4:0] result;
input [22:0] valueIn;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_22;
wire n_0_27;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_28;
wire n_0_29;


NOR4_X1 i_0_45 (.ZN (n_0_29), .A1 (valueIn[14]), .A2 (valueIn[13]), .A3 (valueIn[12]), .A4 (valueIn[11]));
OR2_X1 i_0_44 (.ZN (n_0_28), .A1 (valueIn[6]), .A2 (valueIn[5]));
NOR2_X1 i_0_43 (.ZN (n_0_26), .A1 (valueIn[10]), .A2 (valueIn[9]));
NOR2_X1 i_0_42 (.ZN (n_0_25), .A1 (valueIn[8]), .A2 (valueIn[7]));
NOR4_X1 i_0_41 (.ZN (n_0_24), .A1 (valueIn[18]), .A2 (valueIn[17]), .A3 (valueIn[16]), .A4 (valueIn[15]));
NOR4_X1 i_0_40 (.ZN (n_0_23), .A1 (valueIn[22]), .A2 (valueIn[21]), .A3 (valueIn[20]), .A4 (valueIn[19]));
INV_X1 i_0_39 (.ZN (n_0_21), .A (n_0_23));
NOR3_X1 i_0_38 (.ZN (n_0_20), .A1 (valueIn[3]), .A2 (n_0_28), .A3 (valueIn[4]));
NAND2_X1 i_0_37 (.ZN (n_0_19), .A1 (n_0_26), .A2 (n_0_25));
OAI21_X1 i_0_36 (.ZN (n_0_18), .A (n_0_29), .B1 (n_0_20), .B2 (n_0_19));
AOI21_X1 i_0_35 (.ZN (result[2]), .A (n_0_21), .B1 (n_0_24), .B2 (n_0_18));
INV_X1 i_0_34 (.ZN (n_0_40), .A (valueIn[21]));
INV_X1 i_0_33 (.ZN (n_0_39), .A (valueIn[20]));
INV_X1 i_0_32 (.ZN (n_0_38), .A (valueIn[17]));
INV_X1 i_0_31 (.ZN (n_0_37), .A (valueIn[16]));
INV_X1 i_0_30 (.ZN (n_0_36), .A (valueIn[13]));
INV_X1 i_0_29 (.ZN (n_0_35), .A (valueIn[12]));
INV_X1 i_0_28 (.ZN (n_0_34), .A (valueIn[9]));
INV_X1 i_0_27 (.ZN (n_0_33), .A (valueIn[8]));
INV_X1 i_0_26 (.ZN (n_0_32), .A (valueIn[5]));
INV_X1 i_0_25 (.ZN (n_0_31), .A (valueIn[4]));
INV_X1 i_0_24 (.ZN (n_0_30), .A (valueIn[1]));
NAND2_X1 i_0_23 (.ZN (n_0_27), .A1 (n_0_23), .A2 (n_0_24));
NAND3_X1 i_0_22 (.ZN (n_0_22), .A1 (n_0_29), .A2 (n_0_26), .A3 (n_0_25));
NOR2_X1 i_0_21 (.ZN (result[4]), .A1 (n_0_27), .A2 (n_0_22));
AND3_X1 i_0_20 (.ZN (result[3]), .A1 (n_0_22), .A2 (n_0_24), .A3 (n_0_23));
NOR2_X1 i_0_19 (.ZN (n_0_17), .A1 (valueIn[2]), .A2 (valueIn[1]));
NOR3_X1 i_0_18 (.ZN (n_0_16), .A1 (valueIn[4]), .A2 (valueIn[3]), .A3 (n_0_17));
OAI21_X1 i_0_17 (.ZN (n_0_15), .A (n_0_25), .B1 (n_0_16), .B2 (n_0_28));
AOI211_X1 i_0_16 (.ZN (n_0_14), .A (valueIn[12]), .B (valueIn[11]), .C1 (n_0_15), .C2 (n_0_26));
NOR3_X1 i_0_15 (.ZN (n_0_13), .A1 (valueIn[14]), .A2 (valueIn[13]), .A3 (n_0_14));
NOR3_X1 i_0_14 (.ZN (n_0_12), .A1 (valueIn[16]), .A2 (valueIn[15]), .A3 (n_0_13));
NOR3_X1 i_0_13 (.ZN (n_0_11), .A1 (valueIn[18]), .A2 (valueIn[17]), .A3 (n_0_12));
NOR3_X1 i_0_12 (.ZN (n_0_10), .A1 (valueIn[20]), .A2 (valueIn[19]), .A3 (n_0_11));
NOR3_X1 i_0_11 (.ZN (result[1]), .A1 (valueIn[22]), .A2 (valueIn[21]), .A3 (n_0_10));
AOI21_X1 i_0_10 (.ZN (n_0_9), .A (valueIn[2]), .B1 (n_0_30), .B2 (valueIn[0]));
OAI21_X1 i_0_9 (.ZN (n_0_8), .A (n_0_31), .B1 (valueIn[3]), .B2 (n_0_9));
AOI21_X1 i_0_8 (.ZN (n_0_7), .A (valueIn[6]), .B1 (n_0_32), .B2 (n_0_8));
OAI21_X1 i_0_7 (.ZN (n_0_6), .A (n_0_33), .B1 (valueIn[7]), .B2 (n_0_7));
AOI21_X1 i_0_6 (.ZN (n_0_5), .A (valueIn[10]), .B1 (n_0_34), .B2 (n_0_6));
OAI21_X1 i_0_5 (.ZN (n_0_4), .A (n_0_35), .B1 (valueIn[11]), .B2 (n_0_5));
AOI21_X1 i_0_4 (.ZN (n_0_3), .A (valueIn[14]), .B1 (n_0_36), .B2 (n_0_4));
OAI21_X1 i_0_3 (.ZN (n_0_2), .A (n_0_37), .B1 (valueIn[15]), .B2 (n_0_3));
AOI21_X1 i_0_2 (.ZN (n_0_1), .A (valueIn[18]), .B1 (n_0_38), .B2 (n_0_2));
OAI21_X1 i_0_1 (.ZN (n_0_0), .A (n_0_39), .B1 (valueIn[19]), .B2 (n_0_1));
AOI21_X1 i_0_0 (.ZN (result[0]), .A (valueIn[22]), .B1 (n_0_40), .B2 (n_0_0));

endmodule //count_leading_zeros

module CLA_4bit (a, b, cin, sum, cout);

output cout;
output [3:0] sum;
input [3:0] a;
input [3:0] b;
input cin;


XOR2_X1 i_0_0 (.Z (sum[0]), .A (a[3]), .B (cin));

endmodule //CLA_4bit

module CLA_4bit__0_114 (a, b, cin, sum, cout);

output cout;
output [3:0] sum;
input [3:0] a;
input [3:0] b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


XOR2_X1 i_0_14 (.Z (n_0_9), .A (b[0]), .B (a[0]));
AOI22_X1 i_0_13 (.ZN (n_0_8), .A1 (b[0]), .A2 (a[0]), .B1 (cin), .B2 (n_0_9));
INV_X1 i_0_12 (.ZN (n_0_7), .A (n_0_8));
XOR2_X1 i_0_11 (.Z (n_0_6), .A (b[1]), .B (a[1]));
AOI22_X1 i_0_10 (.ZN (n_0_5), .A1 (b[1]), .A2 (a[1]), .B1 (n_0_7), .B2 (n_0_6));
INV_X1 i_0_9 (.ZN (n_0_4), .A (n_0_5));
XOR2_X1 i_0_8 (.Z (n_0_3), .A (b[2]), .B (a[2]));
AOI22_X1 i_0_7 (.ZN (n_0_2), .A1 (b[2]), .A2 (a[2]), .B1 (n_0_4), .B2 (n_0_3));
NAND2_X1 i_0_6 (.ZN (n_0_1), .A1 (b[3]), .A2 (a[3]));
OAI21_X1 i_0_5 (.ZN (n_0_0), .A (n_0_1), .B1 (b[3]), .B2 (a[3]));
XOR2_X1 i_0_4 (.Z (sum[3]), .A (n_0_2), .B (n_0_0));
XNOR2_X1 i_0_3 (.ZN (sum[2]), .A (n_0_5), .B (n_0_3));
XNOR2_X1 i_0_2 (.ZN (sum[1]), .A (n_0_8), .B (n_0_6));
XOR2_X1 i_0_1 (.Z (sum[0]), .A (cin), .B (n_0_9));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_1), .B1 (n_0_2), .B2 (n_0_0));

endmodule //CLA_4bit__0_114

module CLA_4bit__0_106 (a, b, cin, sum, cout);

output cout;
output [3:0] sum;
input [3:0] a;
input [3:0] b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


XOR2_X1 i_0_14 (.Z (n_0_9), .A (b[0]), .B (a[0]));
AOI22_X1 i_0_13 (.ZN (n_0_8), .A1 (b[0]), .A2 (a[0]), .B1 (cin), .B2 (n_0_9));
INV_X1 i_0_12 (.ZN (n_0_7), .A (n_0_8));
XOR2_X1 i_0_11 (.Z (n_0_6), .A (b[1]), .B (a[1]));
AOI22_X1 i_0_10 (.ZN (n_0_5), .A1 (b[1]), .A2 (a[1]), .B1 (n_0_7), .B2 (n_0_6));
INV_X1 i_0_9 (.ZN (n_0_4), .A (n_0_5));
XOR2_X1 i_0_8 (.Z (n_0_3), .A (b[2]), .B (a[2]));
AOI22_X1 i_0_7 (.ZN (n_0_2), .A1 (b[2]), .A2 (a[2]), .B1 (n_0_4), .B2 (n_0_3));
NAND2_X1 i_0_6 (.ZN (n_0_1), .A1 (b[3]), .A2 (a[3]));
OAI21_X1 i_0_5 (.ZN (n_0_0), .A (n_0_1), .B1 (b[3]), .B2 (a[3]));
XOR2_X1 i_0_4 (.Z (sum[3]), .A (n_0_2), .B (n_0_0));
XNOR2_X1 i_0_3 (.ZN (sum[2]), .A (n_0_5), .B (n_0_3));
XNOR2_X1 i_0_2 (.ZN (sum[1]), .A (n_0_8), .B (n_0_6));
XOR2_X1 i_0_1 (.Z (sum[0]), .A (cin), .B (n_0_9));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_1), .B1 (n_0_2), .B2 (n_0_0));

endmodule //CLA_4bit__0_106

module CLA_4bit__0_98 (a, b, cin, sum, cout);

output cout;
output [3:0] sum;
input [3:0] a;
input [3:0] b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


XOR2_X1 i_0_14 (.Z (n_0_9), .A (b[0]), .B (a[0]));
AOI22_X1 i_0_13 (.ZN (n_0_8), .A1 (b[0]), .A2 (a[0]), .B1 (cin), .B2 (n_0_9));
INV_X1 i_0_12 (.ZN (n_0_7), .A (n_0_8));
XOR2_X1 i_0_11 (.Z (n_0_6), .A (b[1]), .B (a[1]));
AOI22_X1 i_0_10 (.ZN (n_0_5), .A1 (b[1]), .A2 (a[1]), .B1 (n_0_7), .B2 (n_0_6));
INV_X1 i_0_9 (.ZN (n_0_4), .A (n_0_5));
XOR2_X1 i_0_8 (.Z (n_0_3), .A (b[2]), .B (a[2]));
AOI22_X1 i_0_7 (.ZN (n_0_2), .A1 (b[2]), .A2 (a[2]), .B1 (n_0_4), .B2 (n_0_3));
NAND2_X1 i_0_6 (.ZN (n_0_1), .A1 (b[3]), .A2 (a[3]));
OAI21_X1 i_0_5 (.ZN (n_0_0), .A (n_0_1), .B1 (b[3]), .B2 (a[3]));
XOR2_X1 i_0_4 (.Z (sum[3]), .A (n_0_2), .B (n_0_0));
XNOR2_X1 i_0_3 (.ZN (sum[2]), .A (n_0_5), .B (n_0_3));
XNOR2_X1 i_0_2 (.ZN (sum[1]), .A (n_0_8), .B (n_0_6));
XOR2_X1 i_0_1 (.Z (sum[0]), .A (cin), .B (n_0_9));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_1), .B1 (n_0_2), .B2 (n_0_0));

endmodule //CLA_4bit__0_98

module CLA_4bit__0_90 (a, b, cin, sum, cout);

output cout;
output [3:0] sum;
input [3:0] a;
input [3:0] b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


XOR2_X1 i_0_14 (.Z (n_0_9), .A (b[0]), .B (a[0]));
AOI22_X1 i_0_13 (.ZN (n_0_8), .A1 (b[0]), .A2 (a[0]), .B1 (cin), .B2 (n_0_9));
INV_X1 i_0_12 (.ZN (n_0_7), .A (n_0_8));
XOR2_X1 i_0_11 (.Z (n_0_6), .A (b[1]), .B (a[1]));
AOI22_X1 i_0_10 (.ZN (n_0_5), .A1 (b[1]), .A2 (a[1]), .B1 (n_0_7), .B2 (n_0_6));
INV_X1 i_0_9 (.ZN (n_0_4), .A (n_0_5));
XOR2_X1 i_0_8 (.Z (n_0_3), .A (b[2]), .B (a[2]));
AOI22_X1 i_0_7 (.ZN (n_0_2), .A1 (b[2]), .A2 (a[2]), .B1 (n_0_4), .B2 (n_0_3));
NAND2_X1 i_0_6 (.ZN (n_0_1), .A1 (b[3]), .A2 (a[3]));
OAI21_X1 i_0_5 (.ZN (n_0_0), .A (n_0_1), .B1 (b[3]), .B2 (a[3]));
XOR2_X1 i_0_4 (.Z (sum[3]), .A (n_0_2), .B (n_0_0));
XNOR2_X1 i_0_3 (.ZN (sum[2]), .A (n_0_5), .B (n_0_3));
XNOR2_X1 i_0_2 (.ZN (sum[1]), .A (n_0_8), .B (n_0_6));
XOR2_X1 i_0_1 (.Z (sum[0]), .A (cin), .B (n_0_9));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_1), .B1 (n_0_2), .B2 (n_0_0));

endmodule //CLA_4bit__0_90

module CLA_4bit__0_82 (a, b, cin, sum, cout);

output cout;
output [3:0] sum;
input [3:0] a;
input [3:0] b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;


XOR2_X1 i_0_14 (.Z (n_0_9), .A (b[0]), .B (a[0]));
AOI22_X1 i_0_13 (.ZN (n_0_8), .A1 (b[0]), .A2 (a[0]), .B1 (cin), .B2 (n_0_9));
INV_X1 i_0_12 (.ZN (n_0_7), .A (n_0_8));
XOR2_X1 i_0_11 (.Z (n_0_6), .A (b[1]), .B (a[1]));
AOI22_X1 i_0_10 (.ZN (n_0_5), .A1 (b[1]), .A2 (a[1]), .B1 (n_0_7), .B2 (n_0_6));
INV_X1 i_0_9 (.ZN (n_0_4), .A (n_0_5));
XOR2_X1 i_0_8 (.Z (n_0_3), .A (b[2]), .B (a[2]));
AOI22_X1 i_0_7 (.ZN (n_0_2), .A1 (b[2]), .A2 (a[2]), .B1 (n_0_4), .B2 (n_0_3));
NAND2_X1 i_0_6 (.ZN (n_0_1), .A1 (b[3]), .A2 (a[3]));
OAI21_X1 i_0_5 (.ZN (n_0_0), .A (n_0_1), .B1 (b[3]), .B2 (a[3]));
XOR2_X1 i_0_4 (.Z (sum[3]), .A (n_0_2), .B (n_0_0));
XNOR2_X1 i_0_3 (.ZN (sum[2]), .A (n_0_5), .B (n_0_3));
XNOR2_X1 i_0_2 (.ZN (sum[1]), .A (n_0_8), .B (n_0_6));
XOR2_X1 i_0_1 (.Z (sum[0]), .A (cin), .B (n_0_9));
OAI21_X1 i_0_0 (.ZN (cout), .A (n_0_1), .B1 (n_0_2), .B2 (n_0_0));

endmodule //CLA_4bit__0_82

module CLA_4bit__0_66 (a, b, cin, sum, cout);

output cout;
output [3:0] sum;
input [3:0] a;
input [3:0] b;
input cin;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;


NOR2_X1 i_0_16 (.ZN (n_0_11), .A1 (b[3]), .A2 (a[3]));
NAND2_X1 i_0_15 (.ZN (n_0_10), .A1 (b[3]), .A2 (a[3]));
XOR2_X1 i_0_14 (.Z (n_0_9), .A (b[3]), .B (a[3]));
NOR2_X1 i_0_13 (.ZN (n_0_8), .A1 (b[1]), .A2 (a[1]));
NAND2_X1 i_0_12 (.ZN (n_0_7), .A1 (b[1]), .A2 (a[1]));
NAND2_X1 i_0_11 (.ZN (n_0_6), .A1 (b[0]), .A2 (a[0]));
OAI21_X1 i_0_10 (.ZN (n_0_5), .A (n_0_7), .B1 (n_0_8), .B2 (n_0_6));
AOI21_X1 i_0_9 (.ZN (n_0_4), .A (n_0_5), .B1 (a[2]), .B2 (b[2]));
INV_X1 i_0_8 (.ZN (n_0_3), .A (n_0_4));
OAI21_X1 i_0_7 (.ZN (n_0_2), .A (n_0_3), .B1 (a[2]), .B2 (b[2]));
XNOR2_X2 i_0_6 (.ZN (sum[3]), .A (n_0_9), .B (n_0_2));
XNOR2_X1 i_0_5 (.ZN (n_0_1), .A (b[2]), .B (a[2]));
XNOR2_X1 i_0_4 (.ZN (sum[2]), .A (n_0_5), .B (n_0_1));
XOR2_X1 i_0_3 (.Z (n_0_0), .A (b[1]), .B (a[1]));
XNOR2_X1 i_0_2 (.ZN (sum[1]), .A (n_0_6), .B (n_0_0));
XOR2_X1 i_0_1 (.Z (sum[0]), .A (b[0]), .B (a[0]));
AOI21_X1 i_0_0 (.ZN (cout), .A (n_0_11), .B1 (n_0_10), .B2 (n_0_2));

endmodule //CLA_4bit__0_66

module CLA (in1, in2, cin, sum, cout, of);

output cout;
output of;
output [31:0] sum;
input cin;
input [31:0] in1;
input [31:0] in2;
wire c;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;


CLA_4bit genblk1_24_cla (.sum ({uc_3, uc_4, uc_5, sum[24]}), .a ({in1[31], uc_0, 
    uc_1, uc_2}), .cin (n_4));
CLA_4bit__0_114 genblk1_20_cla (.cout (n_4), .sum ({sum[23], sum[22], sum[21], sum[20]})
    , .a ({in1[23], in1[22], in1[21], in1[20]}), .b ({in2[23], in2[22], in2[21], 
    in2[20]}), .cin (n_3));
CLA_4bit__0_106 genblk1_16_cla (.cout (n_3), .sum ({sum[19], sum[18], sum[17], sum[16]})
    , .a ({in1[19], in1[18], in1[17], in1[16]}), .b ({in2[19], in2[18], in2[17], 
    in2[16]}), .cin (n_2));
CLA_4bit__0_98 genblk1_12_cla (.cout (n_2), .sum ({sum[15], sum[14], sum[13], sum[12]})
    , .a ({in1[15], in1[14], in1[13], in1[12]}), .b ({in2[15], in2[14], in2[13], 
    in2[12]}), .cin (n_1));
CLA_4bit__0_90 genblk1_8_cla (.cout (n_1), .sum ({sum[11], sum[10], sum[9], sum[8]})
    , .a ({in1[11], in1[10], in1[9], in1[8]}), .b ({in2[11], in2[10], in2[9], in2[8]}), .cin (n_0));
CLA_4bit__0_82 genblk1_4_cla (.cout (n_0), .sum ({sum[7], sum[6], sum[5], sum[4]})
    , .a ({in1[7], in1[6], in1[5], in1[4]}), .b ({in2[7], in2[6], in2[5], in2[4]}), .cin (c));
CLA_4bit__0_66 cla1 (.cout (c), .sum ({sum[3], sum[2], sum[1], sum[0]}), .a ({in1[3], 
    in1[2], in1[1], in1[0]}), .b ({in2[3], in2[2], in2[1], in2[0]}));

endmodule //CLA

module fp_adder (A, B, Sum, overflow, underflow);

output [31:0] Sum;
output overflow;
output underflow;
input [31:0] A;
input [31:0] B;
wire \num_leading_zeros[4] ;
wire \num_leading_zeros[3] ;
wire \num_leading_zeros[2] ;
wire \num_leading_zeros[1] ;
wire \num_leading_zeros[0] ;
wire n_0_7;
wire n_0_0;
wire n_0_8;
wire n_0_1;
wire n_0_9;
wire n_0_2;
wire n_0_10;
wire n_0_3;
wire n_0_11;
wire n_0_4;
wire n_0_12;
wire n_0_5;
wire n_0_13;
wire n_0_6;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_97;
wire n_0_98;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_123;
wire n_0_124;
wire n_0_127;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_185;
wire n_0_186;
wire n_0_187;
wire n_0_188;
wire n_0_189;
wire n_0_190;
wire n_0_191;
wire \mant_A[31] ;
wire \mant_A[23] ;
wire \mant_A[22] ;
wire \mant_A[21] ;
wire \mant_A[20] ;
wire \mant_A[19] ;
wire \mant_A[18] ;
wire \mant_A[17] ;
wire \mant_A[16] ;
wire \mant_A[15] ;
wire \mant_A[14] ;
wire \mant_A[13] ;
wire \mant_A[12] ;
wire \mant_A[11] ;
wire \mant_A[10] ;
wire \mant_A[9] ;
wire \mant_A[8] ;
wire \mant_A[7] ;
wire \mant_A[6] ;
wire \mant_A[5] ;
wire \mant_A[4] ;
wire \mant_A[3] ;
wire \mant_A[2] ;
wire \mant_A[1] ;
wire drc_ipo_n4;
wire n_0_203;
wire n_0_204;
wire n_0_205;
wire n_0_206;
wire n_0_207;
wire n_0_208;
wire n_0_209;
wire n_0_210;
wire n_0_211;
wire n_0_212;
wire n_0_213;
wire n_0_214;
wire n_0_215;
wire n_0_216;
wire n_0_217;
wire n_0_218;
wire n_0_219;
wire n_0_220;
wire n_0_221;
wire n_0_222;
wire n_0_223;
wire n_0_224;
wire n_0_225;
wire n_0_226;
wire n_0_227;
wire n_0_228;
wire n_0_229;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_233;
wire n_0_234;
wire n_0_235;
wire n_0_236;
wire n_0_237;
wire n_0_238;
wire n_0_239;
wire n_0_240;
wire n_0_241;
wire n_0_242;
wire n_0_243;
wire n_0_244;
wire n_0_245;
wire n_0_246;
wire n_0_247;
wire n_0_248;
wire n_0_249;
wire n_0_250;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_257;
wire n_0_258;
wire n_0_259;
wire n_0_260;
wire n_0_261;
wire \exp_Sum[7] ;
wire \exp_Sum[6] ;
wire \exp_Sum[5] ;
wire \exp_Sum[4] ;
wire \exp_Sum[3] ;
wire \exp_Sum[2] ;
wire \exp_Sum[1] ;
wire \exp_Sum[0] ;
wire n_0_262;
wire n_0_263;
wire n_0_264;
wire n_0_265;
wire n_0_266;
wire n_0_267;
wire n_0_268;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_272;
wire n_0_273;
wire n_0_274;
wire n_0_275;
wire n_0_276;
wire n_0_277;
wire n_0_278;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_282;
wire n_0_283;
wire n_0_284;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_288;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_296;
wire n_0_297;
wire n_0_298;
wire n_0_299;
wire n_0_300;
wire n_0_301;
wire n_0_302;
wire n_0_303;
wire n_0_304;
wire n_0_305;
wire n_0_311;
wire n_0_317;
wire n_0_318;
wire n_0_320;
wire n_0_321;
wire n_0_322;
wire n_0_328;
wire n_0_329;
wire n_0_330;
wire n_0_331;
wire n_0_332;
wire n_0_334;
wire n_0_335;
wire n_0_336;
wire n_0_337;
wire n_0_338;
wire n_0_339;
wire n_0_340;
wire n_0_341;
wire n_0_342;
wire n_0_343;
wire n_0_344;
wire n_0_346;
wire n_0_347;
wire n_0_348;
wire n_0_349;
wire n_0_350;
wire n_0_351;
wire n_0_355;
wire n_0_356;
wire n_0_357;
wire n_0_358;
wire n_0_359;
wire n_0_360;
wire n_0_363;
wire n_0_364;
wire n_0_365;
wire n_0_367;
wire n_0_368;
wire n_0_370;
wire n_0_371;
wire n_0_372;
wire n_0_373;
wire n_0_376;
wire n_0_377;
wire n_0_378;
wire n_0_379;
wire n_0_380;
wire n_0_381;
wire n_0_382;
wire n_0_396;
wire n_0_397;
wire n_0_398;
wire n_0_399;
wire n_0_400;
wire n_0_401;
wire n_0_402;
wire n_0_403;
wire n_0_404;
wire n_0_405;
wire n_0_406;
wire n_0_407;
wire n_0_408;
wire n_0_409;
wire n_0_410;
wire n_0_411;
wire n_0_412;
wire n_0_413;
wire n_0_414;
wire n_0_415;
wire n_0_416;
wire n_0_417;
wire n_0_418;
wire n_0_419;
wire n_0_420;
wire n_0_426;
wire n_0_431;
wire n_0_432;
wire n_0_437;
wire n_0_438;
wire n_0_443;
wire n_0_444;
wire n_0_445;
wire n_0_446;
wire n_0_447;
wire n_0_448;
wire n_0_449;
wire n_0_451;
wire n_0_452;
wire n_0_453;
wire n_0_454;
wire n_0_455;
wire n_0_456;
wire n_0_457;
wire n_0_458;
wire n_0_459;
wire n_0_460;
wire n_0_461;
wire n_0_462;
wire n_0_463;
wire n_0_464;
wire n_0_465;
wire n_0_466;
wire n_0_467;
wire n_0_468;
wire n_0_469;
wire n_0_472;
wire n_0_473;
wire n_0_474;
wire n_0_475;
wire n_0_476;
wire n_0_477;
wire n_0_478;
wire n_0_479;
wire n_0_480;
wire n_0_481;
wire n_0_482;
wire n_0_483;
wire n_0_485;
wire n_0_486;
wire n_0_487;
wire n_0_488;
wire n_0_489;
wire n_0_490;
wire n_0_491;
wire n_0_494;
wire n_0_496;
wire n_0_497;
wire n_0_498;
wire n_0_499;
wire n_0_500;
wire n_0_501;
wire n_0_502;
wire n_0_504;
wire n_0_515;
wire n_0_95;
wire n_0_532;
wire n_0_563;
wire n_0_564;
wire n_0_578;
wire n_0_579;
wire n_0_580;
wire n_0_581;
wire n_0_582;
wire n_0_583;
wire n_0_584;
wire n_0_585;
wire n_0_586;
wire n_0_587;
wire n_0_588;
wire n_0_96;
wire n_0_603;
wire n_0_604;
wire n_0_605;
wire n_0_606;
wire n_0_607;
wire n_0_608;
wire n_0_609;
wire n_0_610;
wire n_0_611;
wire n_0_612;
wire n_0_613;
wire n_0_99;
wire n_0_94;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_125;
wire n_0_126;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_192;
wire n_0_193;
wire n_0_194;
wire n_0_195;
wire n_0_196;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_201;
wire n_0_202;
wire n_0_306;
wire n_0_307;
wire n_0_308;
wire n_0_309;
wire n_0_310;
wire n_0_312;
wire n_0_313;
wire n_0_314;
wire n_0_315;
wire n_0_316;
wire n_0_319;
wire n_0_323;
wire n_0_324;
wire n_0_325;
wire n_0_326;
wire n_0_327;
wire n_0_333;
wire n_0_345;
wire n_0_352;
wire n_0_353;
wire n_0_354;
wire n_0_361;
wire n_0_362;
wire n_0_366;
wire n_0_369;
wire n_0_374;
wire n_0_375;
wire n_0_383;
wire n_0_384;
wire n_0_385;
wire n_0_386;
wire n_0_387;
wire n_0_388;
wire n_0_389;
wire n_0_390;
wire n_0_391;
wire n_0_392;
wire n_0_393;
wire n_0_394;
wire n_0_395;
wire n_0_421;
wire n_0_422;
wire n_0_423;
wire n_0_424;
wire n_0_425;
wire n_0_427;
wire n_0_428;
wire n_0_429;
wire n_0_430;
wire n_0_433;
wire n_0_434;
wire n_0_435;
wire n_0_436;
wire n_0_439;
wire n_0_440;
wire n_0_441;
wire n_0_442;
wire n_0_450;
wire n_0_470;
wire n_0_471;
wire n_0_484;
wire n_0_492;
wire n_0_493;
wire n_0_495;
wire n_0_503;
wire n_0_505;
wire n_0_506;
wire n_0_507;
wire n_0_508;
wire n_0_509;
wire n_0_510;
wire n_0_511;
wire n_0_512;
wire n_0_513;
wire n_0_514;
wire n_0_517;
wire n_0_518;
wire n_0_519;
wire n_0_520;
wire n_0_521;
wire n_0_522;
wire n_0_523;
wire n_0_524;
wire n_0_525;
wire n_0_526;
wire n_0_527;
wire n_0_528;
wire n_0_529;
wire n_0_530;
wire n_0_531;
wire n_0_533;
wire n_0_534;
wire n_0_535;
wire n_0_536;
wire n_0_537;
wire n_0_538;
wire n_0_539;
wire n_0_540;
wire n_0_541;
wire n_0_542;
wire n_0_543;
wire n_0_544;
wire n_0_545;
wire n_0_546;
wire n_0_547;
wire n_0_548;
wire n_0_549;
wire n_0_550;
wire n_0_551;
wire n_0_552;
wire n_0_553;
wire n_0_554;
wire n_0_555;
wire n_0_556;
wire n_0_557;
wire n_0_558;
wire n_0_559;
wire n_0_560;
wire n_0_561;
wire n_0_562;
wire n_0_565;
wire n_0_566;
wire n_0_567;
wire n_0_568;
wire n_0_569;
wire n_0_570;
wire n_0_571;
wire n_0_572;
wire n_0_573;
wire n_0_574;
wire n_0_575;
wire n_0_576;
wire n_0_577;
wire n_0_589;
wire n_0_590;
wire n_0_591;
wire n_0_592;
wire n_0_593;
wire n_0_594;
wire n_0_595;
wire n_0_596;
wire n_0_597;
wire n_0_598;
wire n_0_599;
wire n_0_600;
wire n_0_601;
wire n_0_602;
wire n_0_614;
wire n_0_615;
wire n_0_616;
wire n_0_617;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire n_55;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire n_102;
wire n_98;
wire n_97;
wire n_96;
wire n_95;
wire n_94;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_101;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire n_0;
wire n_25;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_100;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_99;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_54;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire uc_35;


OAI21_X1 i_0_724 (.ZN (n_0_617), .A (n_0_527), .B1 (n_0_518), .B2 (n_0_505));
INV_X1 i_0_723 (.ZN (n_102), .A (n_0_617));
NAND2_X1 i_0_722 (.ZN (n_0_616), .A1 (n_0_537), .A2 (n_0_533));
NOR3_X1 i_0_721 (.ZN (n_0_615), .A1 (n_0_535), .A2 (A[28]), .A3 (n_0_544));
AOI21_X1 i_0_720 (.ZN (n_0_614), .A (n_0_530), .B1 (n_0_616), .B2 (n_0_615));
OAI21_X1 i_0_719 (.ZN (n_0_602), .A (n_0_517), .B1 (n_0_520), .B2 (n_0_614));
AND2_X1 i_0_718 (.ZN (n_0_601), .A1 (n_0_617), .A2 (n_0_602));
AND2_X1 i_0_717 (.ZN (n_0_600), .A1 (n_0_539), .A2 (n_0_601));
NAND2_X1 i_0_715 (.ZN (n_0_599), .A1 (n_0_510), .A2 (n_0_540));
OAI21_X2 i_0_713 (.ZN (n_0_598), .A (n_0_599), .B1 (n_0_540), .B2 (n_0_450));
INV_X1 i_0_710 (.ZN (n_0_597), .A (n_0_598));
NOR2_X1 i_0_709 (.ZN (n_0_596), .A1 (n_0_514), .A2 (n_0_95));
NAND2_X1 i_0_708 (.ZN (n_0_595), .A1 (n_0_513), .A2 (n_0_596));
OAI21_X1 i_0_707 (.ZN (n_0_594), .A (n_0_595), .B1 (n_0_513), .B2 (n_0_596));
INV_X1 i_0_706 (.ZN (n_0_593), .A (n_0_594));
OAI21_X1 i_0_705 (.ZN (n_0_592), .A (n_0_524), .B1 (n_0_526), .B2 (n_0_525));
XOR2_X1 i_0_704 (.Z (n_0_591), .A (n_0_523), .B (n_0_436));
INV_X1 i_0_703 (.ZN (n_0_590), .A (n_0_591));
NOR2_X1 i_0_702 (.ZN (n_0_589), .A1 (n_0_592), .A2 (n_0_591));
INV_X1 i_0_701 (.ZN (n_0_577), .A (n_0_589));
NOR2_X2 i_0_700 (.ZN (n_0_576), .A1 (n_0_593), .A2 (n_0_577));
NAND2_X1 i_0_699 (.ZN (n_0_575), .A1 (n_0_593), .A2 (n_0_589));
NAND2_X1 i_0_698 (.ZN (n_0_574), .A1 (n_0_592), .A2 (n_0_590));
INV_X1 i_0_697 (.ZN (n_0_573), .A (n_0_574));
NOR2_X1 i_0_696 (.ZN (n_0_572), .A1 (n_0_594), .A2 (n_0_574));
NOR2_X1 i_0_695 (.ZN (n_0_571), .A1 (n_0_593), .A2 (n_0_574));
NAND2_X1 i_0_694 (.ZN (n_0_570), .A1 (B[12]), .A2 (n_0_576));
OAI21_X1 i_0_693 (.ZN (n_0_569), .A (n_0_570), .B1 (n_0_314), .B2 (n_0_575));
AOI221_X1 i_0_686 (.ZN (n_0_568), .A (n_0_569), .B1 (B[16]), .B2 (n_0_572), .C1 (B[20]), .C2 (n_0_571));
AOI22_X1 i_0_684 (.ZN (n_0_567), .A1 (B[10]), .A2 (n_0_589), .B1 (B[18]), .B2 (n_0_573));
NOR2_X1 i_0_683 (.ZN (n_0_566), .A1 (n_0_592), .A2 (n_0_590));
AOI222_X1 i_0_682 (.ZN (n_0_565), .A1 (B[22]), .A2 (n_0_566), .B1 (B[6]), .B2 (n_0_589)
    , .C1 (B[14]), .C2 (n_0_573));
OAI22_X1 i_0_681 (.ZN (n_0_562), .A1 (n_0_594), .A2 (n_0_565), .B1 (n_0_593), .B2 (n_0_567));
INV_X1 i_0_680 (.ZN (n_0_561), .A (n_0_562));
OAI22_X1 i_0_679 (.ZN (n_0_560), .A1 (n_0_598), .A2 (n_0_561), .B1 (n_0_597), .B2 (n_0_568));
NAND2_X1 i_0_678 (.ZN (n_0_559), .A1 (n_0_540), .A2 (n_0_601));
INV_X1 i_0_677 (.ZN (n_0_558), .A (n_0_559));
AOI22_X1 i_0_676 (.ZN (n_0_557), .A1 (B[21]), .A2 (n_0_566), .B1 (B[13]), .B2 (n_0_573));
OAI21_X1 i_0_675 (.ZN (n_0_556), .A (n_0_557), .B1 (n_0_308), .B2 (n_0_577));
AOI222_X1 i_0_674 (.ZN (n_0_555), .A1 (B[9]), .A2 (n_0_576), .B1 (B[17]), .B2 (n_0_571)
    , .C1 (n_0_593), .C2 (n_0_556));
NAND2_X1 i_0_673 (.ZN (n_0_554), .A1 (B[15]), .A2 (n_0_590));
AOI22_X1 i_0_672 (.ZN (n_0_553), .A1 (n_0_592), .A2 (n_0_554), .B1 (n_0_312), .B2 (n_0_589));
AOI222_X1 i_0_671 (.ZN (n_0_552), .A1 (n_0_593), .A2 (n_0_553), .B1 (B[11]), .B2 (n_0_576)
    , .C1 (B[19]), .C2 (n_0_571));
OAI22_X1 i_0_670 (.ZN (n_0_551), .A1 (n_0_597), .A2 (n_0_552), .B1 (n_0_598), .B2 (n_0_555));
AOI222_X1 i_0_669 (.ZN (n_0_550), .A1 (n_0_600), .A2 (n_0_560), .B1 (B[5]), .B2 (n_102)
    , .C1 (n_0_558), .C2 (n_0_551));
INV_X1 i_0_668 (.ZN (n_101), .A (n_0_550));
INV_X1 i_0_667 (.ZN (n_0_549), .A (A[28]));
INV_X1 i_0_666 (.ZN (n_0_548), .A (A[25]));
INV_X1 i_0_665 (.ZN (n_0_547), .A (A[23]));
INV_X1 i_0_664 (.ZN (n_0_546), .A (B[30]));
INV_X1 i_0_663 (.ZN (n_0_545), .A (B[29]));
INV_X1 i_0_662 (.ZN (n_0_544), .A (B[28]));
INV_X1 i_0_661 (.ZN (n_0_543), .A (B[27]));
INV_X1 i_0_660 (.ZN (n_0_542), .A (B[26]));
NOR2_X1 i_0_659 (.ZN (n_0_541), .A1 (n_0_547), .A2 (B[23]));
AOI21_X1 i_0_658 (.ZN (n_0_540), .A (n_0_541), .B1 (n_0_547), .B2 (B[23]));
INV_X1 i_0_657 (.ZN (n_0_539), .A (n_0_540));
NOR2_X1 i_0_656 (.ZN (n_0_538), .A1 (A[30]), .A2 (B[30]));
AOI21_X1 i_0_655 (.ZN (n_0_537), .A (n_0_538), .B1 (A[30]), .B2 (B[30]));
INV_X1 i_0_654 (.ZN (n_0_536), .A (n_0_537));
AOI21_X1 i_0_653 (.ZN (n_0_535), .A (n_0_537), .B1 (A[29]), .B2 (n_0_545));
NOR2_X1 i_0_652 (.ZN (n_0_534), .A1 (A[29]), .A2 (n_0_545));
INV_X1 i_0_651 (.ZN (n_0_533), .A (n_0_534));
NAND2_X1 i_0_650 (.ZN (n_0_531), .A1 (n_0_535), .A2 (n_0_533));
NOR3_X1 i_0_649 (.ZN (n_0_530), .A1 (n_0_549), .A2 (B[28]), .A3 (n_0_531));
NOR2_X1 i_0_648 (.ZN (n_0_529), .A1 (A[30]), .A2 (n_0_546));
NOR2_X1 i_0_647 (.ZN (n_0_528), .A1 (n_0_535), .A2 (n_0_529));
NOR2_X1 i_0_646 (.ZN (n_0_527), .A1 (n_0_530), .A2 (n_0_528));
XOR2_X1 i_0_645 (.Z (n_0_526), .A (A[26]), .B (n_0_542));
OAI21_X1 i_0_644 (.ZN (n_0_525), .A (n_0_595), .B1 (A[25]), .B2 (n_0_99));
NAND2_X1 i_0_643 (.ZN (n_0_524), .A1 (n_0_526), .A2 (n_0_525));
OAI21_X1 i_0_642 (.ZN (n_0_523), .A (n_0_524), .B1 (A[26]), .B2 (n_0_542));
NAND2_X1 i_0_641 (.ZN (n_0_522), .A1 (A[27]), .A2 (n_0_543));
NOR2_X1 i_0_640 (.ZN (n_0_521), .A1 (A[27]), .A2 (n_0_543));
OAI21_X1 i_0_639 (.ZN (n_0_520), .A (n_0_522), .B1 (n_0_523), .B2 (n_0_521));
AOI211_X1 i_0_638 (.ZN (n_0_519), .A (n_0_529), .B (n_0_534), .C1 (n_0_549), .C2 (B[28]));
INV_X1 i_0_637 (.ZN (n_0_518), .A (n_0_519));
NAND3_X1 i_0_636 (.ZN (n_0_517), .A1 (n_0_527), .A2 (n_0_520), .A3 (n_0_519));
NAND2_X2 i_0_635 (.ZN (n_100), .A1 (n_0_527), .A2 (n_0_517));
NOR2_X1 i_0_633 (.ZN (n_0_514), .A1 (B[24]), .A2 (n_0_96));
OAI22_X1 i_0_632 (.ZN (n_0_513), .A1 (A[25]), .A2 (B[25]), .B1 (n_0_548), .B2 (n_0_99));
INV_X1 i_0_631 (.ZN (n_0_512), .A (n_0_513));
AOI21_X1 i_0_630 (.ZN (n_0_511), .A (n_0_514), .B1 (B[24]), .B2 (n_0_96));
INV_X1 i_0_629 (.ZN (n_0_510), .A (n_0_511));
AOI21_X1 i_0_628 (.ZN (n_0_509), .A (n_0_514), .B1 (n_0_541), .B2 (n_0_511));
OAI22_X1 i_0_627 (.ZN (n_0_508), .A1 (n_0_548), .A2 (B[25]), .B1 (n_0_512), .B2 (n_0_509));
AOI22_X1 i_0_626 (.ZN (n_0_507), .A1 (A[26]), .A2 (n_0_542), .B1 (n_0_526), .B2 (n_0_508));
AOI21_X1 i_0_625 (.ZN (n_0_506), .A (n_0_521), .B1 (n_0_522), .B2 (n_0_507));
INV_X1 i_0_624 (.ZN (n_0_505), .A (n_0_506));
AOI22_X1 i_0_623 (.ZN (n_0_503), .A1 (A[29]), .A2 (n_0_545), .B1 (n_0_536), .B2 (n_0_534));
OAI33_X1 i_0_622 (.ZN (n_0_495), .A1 (n_0_549), .A2 (B[28]), .A3 (n_0_503), .B1 (A[28])
    , .B2 (n_0_544), .B3 (n_0_531));
OAI221_X1 i_0_621 (.ZN (n_0_493), .A (n_0_396), .B1 (n_0_519), .B2 (n_0_506), .C1 (n_0_505), .C2 (n_0_495));
INV_X1 i_0_620 (.ZN (n_0_492), .A (n_0_493));
NOR2_X2 i_0_619 (.ZN (n_0_484), .A1 (n_0_539), .A2 (n_0_493));
INV_X1 i_0_618 (.ZN (n_0_471), .A (n_0_484));
XOR2_X1 i_0_617 (.Z (n_0_470), .A (n_0_541), .B (n_0_511));
INV_X1 i_0_616 (.ZN (n_0_450), .A (drc_ipo_n4));
XOR2_X1 i_0_615 (.Z (n_0_442), .A (n_0_512), .B (n_0_509));
INV_X1 i_0_614 (.ZN (n_0_441), .A (n_0_442));
XOR2_X1 i_0_613 (.Z (n_0_440), .A (n_0_526), .B (n_0_508));
INV_X1 i_0_612 (.ZN (n_0_439), .A (n_0_440));
OAI21_X1 i_0_611 (.ZN (n_0_436), .A (n_0_522), .B1 (A[27]), .B2 (n_0_543));
XOR2_X1 i_0_610 (.Z (n_0_435), .A (n_0_507), .B (n_0_436));
NAND2_X1 i_0_609 (.ZN (n_0_434), .A1 (n_0_439), .A2 (n_0_435));
INV_X1 i_0_608 (.ZN (n_0_433), .A (n_0_434));
NAND2_X1 i_0_607 (.ZN (n_0_430), .A1 (n_0_440), .A2 (n_0_435));
INV_X1 i_0_606 (.ZN (n_0_429), .A (n_0_430));
AOI22_X1 i_0_605 (.ZN (n_0_428), .A1 (A[11]), .A2 (n_0_429), .B1 (A[19]), .B2 (n_0_433));
INV_X1 i_0_604 (.ZN (n_0_427), .A (n_0_428));
NAND2_X1 i_0_602 (.ZN (n_0_425), .A1 (A[15]), .A2 (n_0_435));
AOI22_X1 i_0_601 (.ZN (n_0_424), .A1 (n_0_439), .A2 (n_0_425), .B1 (n_0_310), .B2 (n_0_429));
OAI22_X1 i_0_600 (.ZN (n_0_423), .A1 (n_0_441), .A2 (n_0_424), .B1 (n_0_442), .B2 (n_0_427));
NOR2_X2 i_0_599 (.ZN (n_0_422), .A1 (n_0_441), .A2 (n_0_430));
INV_X1 i_0_598 (.ZN (n_0_421), .A (n_0_422));
OAI22_X1 i_0_597 (.ZN (n_0_395), .A1 (A[21]), .A2 (n_0_442), .B1 (A[17]), .B2 (n_0_441));
NOR2_X1 i_0_596 (.ZN (n_0_394), .A1 (n_0_442), .A2 (n_0_430));
NOR2_X1 i_0_595 (.ZN (n_0_393), .A1 (n_0_434), .A2 (n_0_395));
AOI221_X1 i_0_594 (.ZN (n_0_392), .A (n_0_393), .B1 (A[9]), .B2 (n_0_422), .C1 (A[13]), .C2 (n_0_394));
OAI22_X1 i_0_593 (.ZN (n_0_391), .A1 (drc_ipo_n4), .A2 (n_0_392), .B1 (n_0_450), .B2 (n_0_423));
NOR2_X2 i_0_592 (.ZN (n_0_390), .A1 (n_0_540), .A2 (n_0_493));
NOR2_X1 i_0_591 (.ZN (n_0_389), .A1 (n_0_442), .A2 (n_0_434));
NOR2_X1 i_0_590 (.ZN (n_0_388), .A1 (n_0_441), .A2 (n_0_434));
AOI22_X1 i_0_589 (.ZN (n_0_387), .A1 (A[18]), .A2 (n_0_388), .B1 (A[14]), .B2 (n_0_394));
INV_X1 i_0_588 (.ZN (n_0_386), .A (n_0_387));
AOI221_X1 i_0_587 (.ZN (n_0_385), .A (n_0_386), .B1 (A[22]), .B2 (n_0_389), .C1 (A[10]), .C2 (n_0_422));
INV_X1 i_0_586 (.ZN (n_0_384), .A (n_0_385));
NAND2_X1 i_0_585 (.ZN (n_0_383), .A1 (A[12]), .A2 (n_0_394));
OAI21_X1 i_0_584 (.ZN (n_0_375), .A (n_0_383), .B1 (n_0_313), .B2 (n_0_421));
AOI221_X1 i_0_583 (.ZN (n_0_374), .A (n_0_375), .B1 (A[16]), .B2 (n_0_388), .C1 (A[20]), .C2 (n_0_389));
AOI22_X1 i_0_582 (.ZN (n_0_369), .A1 (drc_ipo_n4), .A2 (n_0_374), .B1 (n_0_450), .B2 (n_0_385));
AOI222_X1 i_0_581 (.ZN (n_0_366), .A1 (n_0_484), .A2 (n_0_391), .B1 (A[7]), .B2 (n_100)
    , .C1 (n_0_390), .C2 (n_0_369));
INV_X1 i_0_580 (.ZN (n_99), .A (n_0_366));
AOI221_X1 i_0_579 (.ZN (n_0_362), .A (n_0_354), .B1 (B[8]), .B2 (n_0_313), .C1 (B[9]), .C2 (n_0_361));
INV_X1 i_0_578 (.ZN (n_0_361), .A (A[9]));
AOI22_X1 i_0_577 (.ZN (n_0_354), .A1 (n_0_352), .A2 (n_0_353), .B1 (n_0_314), .B2 (A[8]));
NAND2_X1 i_0_576 (.ZN (n_0_353), .A1 (n_0_310), .A2 (B[7]));
OAI221_X1 i_0_575 (.ZN (n_0_352), .A (n_0_345), .B1 (n_0_309), .B2 (B[6]), .C1 (B[7]), .C2 (n_0_310));
OAI221_X1 i_0_574 (.ZN (n_0_345), .A (n_0_327), .B1 (A[6]), .B2 (n_0_333), .C1 (n_0_308), .C2 (A[5]));
INV_X1 i_0_573 (.ZN (n_0_333), .A (B[6]));
OAI221_X1 i_0_572 (.ZN (n_0_327), .A (n_0_326), .B1 (n_0_306), .B2 (B[4]), .C1 (B[5]), .C2 (n_0_307));
OAI221_X1 i_0_571 (.ZN (n_0_326), .A (n_0_325), .B1 (A[4]), .B2 (n_0_201), .C1 (n_0_202), .C2 (A[3]));
OAI221_X1 i_0_570 (.ZN (n_0_325), .A (n_0_319), .B1 (B[3]), .B2 (n_0_323), .C1 (n_0_324), .C2 (B[2]));
INV_X1 i_0_569 (.ZN (n_0_324), .A (A[2]));
INV_X1 i_0_568 (.ZN (n_0_323), .A (A[3]));
OAI221_X1 i_0_567 (.ZN (n_0_319), .A (n_0_316), .B1 (n_0_199), .B2 (A[2]), .C1 (n_0_200), .C2 (A[1]));
OAI22_X1 i_0_566 (.ZN (n_0_316), .A1 (n_0_315), .A2 (B[0]), .B1 (n_0_198), .B2 (B[1]));
INV_X1 i_0_565 (.ZN (n_0_315), .A (A[0]));
INV_X1 i_0_564 (.ZN (n_0_314), .A (B[8]));
INV_X1 i_0_563 (.ZN (n_0_313), .A (A[8]));
INV_X1 i_0_562 (.ZN (n_0_312), .A (B[7]));
INV_X1 i_0_561 (.ZN (n_0_310), .A (A[7]));
INV_X1 i_0_560 (.ZN (n_0_309), .A (A[6]));
INV_X1 i_0_559 (.ZN (n_0_308), .A (B[5]));
INV_X1 i_0_558 (.ZN (n_0_307), .A (A[5]));
INV_X1 i_0_557 (.ZN (n_0_306), .A (A[4]));
INV_X1 i_0_556 (.ZN (n_0_202), .A (B[3]));
INV_X1 i_0_555 (.ZN (n_0_201), .A (B[4]));
INV_X1 i_0_554 (.ZN (n_0_200), .A (B[1]));
INV_X1 i_0_553 (.ZN (n_0_199), .A (B[2]));
INV_X1 i_0_552 (.ZN (n_0_198), .A (A[1]));
AOI222_X1 i_0_551 (.ZN (n_0_197), .A1 (n_18), .A2 (n_0_114), .B1 (n_2), .B2 (n_0_122)
    , .C1 (n_10), .C2 (n_0_120));
AOI22_X1 i_0_550 (.ZN (n_0_196), .A1 (n_14), .A2 (n_0_114), .B1 (n_6), .B2 (n_0_120));
OAI22_X1 i_0_549 (.ZN (n_0_195), .A1 (n_28), .A2 (n_0_197), .B1 (n_0_126), .B2 (n_0_196));
AOI222_X1 i_0_548 (.ZN (n_0_194), .A1 (n_16), .A2 (n_0_114), .B1 (n_0), .B2 (n_0_122)
    , .C1 (n_8), .C2 (n_0_120));
AOI222_X1 i_0_547 (.ZN (n_0_193), .A1 (n_20), .A2 (n_0_113), .B1 (n_12), .B2 (n_0_119)
    , .C1 (n_4), .C2 (n_0_121));
OAI21_X1 i_0_546 (.ZN (n_0_192), .A (n_0_193), .B1 (n_0_126), .B2 (n_0_194));
INV_X1 i_0_545 (.ZN (n_0_132), .A (n_0_192));
NAND2_X1 i_0_544 (.ZN (n_0_131), .A1 (n_27), .A2 (n_0_195));
OAI21_X1 i_0_543 (.ZN (n_0_130), .A (n_0_131), .B1 (n_27), .B2 (n_0_132));
INV_X1 i_0_542 (.ZN (n_0_129), .A (n_30));
INV_X1 i_0_541 (.ZN (n_0_128), .A (n_29));
INV_X1 i_0_540 (.ZN (n_0_126), .A (n_28));
INV_X1 i_0_539 (.ZN (n_0_125), .A (n_27));
NOR2_X1 i_0_538 (.ZN (n_0_122), .A1 (n_0_129), .A2 (n_29));
NOR3_X1 i_0_537 (.ZN (n_0_121), .A1 (n_0_129), .A2 (n_29), .A3 (n_28));
NOR2_X1 i_0_536 (.ZN (n_0_120), .A1 (n_30), .A2 (n_0_128));
NOR3_X2 i_0_535 (.ZN (n_0_119), .A1 (n_30), .A2 (n_0_128), .A3 (n_28));
NOR2_X1 i_0_534 (.ZN (n_0_114), .A1 (n_30), .A2 (n_29));
NOR3_X4 i_0_533 (.ZN (n_0_113), .A1 (n_30), .A2 (n_29), .A3 (n_28));
AOI22_X1 i_0_532 (.ZN (n_0_112), .A1 (n_15), .A2 (n_0_114), .B1 (n_7), .B2 (n_0_120));
AOI222_X1 i_0_531 (.ZN (n_0_111), .A1 (n_19), .A2 (n_0_113), .B1 (n_11), .B2 (n_0_119)
    , .C1 (n_3), .C2 (n_0_121));
OAI21_X1 i_0_530 (.ZN (n_0_110), .A (n_0_111), .B1 (n_0_126), .B2 (n_0_112));
AOI22_X1 i_0_529 (.ZN (n_0_109), .A1 (n_13), .A2 (n_0_114), .B1 (n_5), .B2 (n_0_120));
AOI222_X1 i_0_528 (.ZN (n_0_102), .A1 (n_9), .A2 (n_0_120), .B1 (n_1), .B2 (n_0_122)
    , .C1 (n_17), .C2 (n_0_114));
AOI22_X1 i_0_527 (.ZN (n_0_101), .A1 (n_0_126), .A2 (n_0_102), .B1 (n_28), .B2 (n_0_109));
OAI22_X1 i_0_526 (.ZN (n_0_100), .A1 (n_27), .A2 (n_0_110), .B1 (n_0_125), .B2 (n_0_101));
INV_X1 i_0_525 (.ZN (n_0_94), .A (B[31]));
INV_X1 i_0_524 (.ZN (n_0_99), .A (B[25]));
INV_X1 i_0_523 (.ZN (n_0_613), .A (B[22]));
INV_X1 i_0_522 (.ZN (n_0_612), .A (B[20]));
INV_X1 i_0_521 (.ZN (n_0_611), .A (B[19]));
INV_X1 i_0_520 (.ZN (n_0_610), .A (B[18]));
INV_X1 i_0_716 (.ZN (n_0_609), .A (B[17]));
INV_X1 i_0_519 (.ZN (n_0_608), .A (B[16]));
INV_X1 i_0_714 (.ZN (n_0_607), .A (B[13]));
INV_X1 i_0_518 (.ZN (n_0_606), .A (B[12]));
INV_X1 i_0_712 (.ZN (n_0_605), .A (B[11]));
INV_X1 i_0_711 (.ZN (n_0_604), .A (B[10]));
INV_X1 i_0_517 (.ZN (n_0_603), .A (B[9]));
INV_X1 i_0_516 (.ZN (n_0_96), .A (A[24]));
INV_X1 i_0_515 (.ZN (n_0_588), .A (A[22]));
INV_X1 i_0_514 (.ZN (n_0_587), .A (A[21]));
INV_X1 i_0_513 (.ZN (n_0_586), .A (A[20]));
INV_X1 i_0_692 (.ZN (n_0_585), .A (A[19]));
INV_X1 i_0_691 (.ZN (n_0_584), .A (A[18]));
INV_X1 i_0_690 (.ZN (n_0_583), .A (A[17]));
INV_X1 i_0_689 (.ZN (n_0_582), .A (A[16]));
INV_X1 i_0_688 (.ZN (n_0_581), .A (A[15]));
INV_X1 i_0_687 (.ZN (n_0_580), .A (A[14]));
INV_X1 i_0_512 (.ZN (n_0_579), .A (A[13]));
INV_X1 i_0_685 (.ZN (n_0_578), .A (A[12]));
INV_X1 i_0_511 (.ZN (n_0_564), .A (n_53));
INV_X1 i_0_510 (.ZN (n_0_563), .A (n_0_6));
INV_X1 i_0_509 (.ZN (\exp_Sum[7] ), .A (n_0_538));
AOI21_X1 i_0_508 (.ZN (n_0_532), .A (B[22]), .B1 (n_0_617), .B2 (n_0_539));
AOI22_X1 i_0_507 (.ZN (n_0_95), .A1 (B[24]), .A2 (n_0_96), .B1 (B[23]), .B2 (n_0_547));
INV_X1 i_0_506 (.ZN (n_0_515), .A (n_0_575));
NAND3_X1 i_0_505 (.ZN (n_0_504), .A1 (n_0_602), .A2 (n_0_597), .A3 (n_0_515));
AOI21_X1 i_0_504 (.ZN (n_98), .A (n_0_532), .B1 (n_0_617), .B2 (n_0_504));
AOI211_X1 i_0_503 (.ZN (n_0_502), .A (drc_ipo_n4), .B (n_0_575), .C1 (n_0_613), .C2 (n_0_539));
AOI22_X1 i_0_502 (.ZN (n_0_501), .A1 (B[21]), .A2 (n_102), .B1 (n_0_601), .B2 (n_0_502));
INV_X1 i_0_501 (.ZN (n_97), .A (n_0_501));
NOR3_X1 i_0_603 (.ZN (n_0_500), .A1 (B[21]), .A2 (n_0_598), .A3 (n_0_540));
AOI22_X1 i_0_500 (.ZN (n_0_499), .A1 (B[22]), .A2 (n_0_598), .B1 (B[20]), .B2 (n_0_597));
INV_X1 i_0_499 (.ZN (n_0_498), .A (n_0_499));
AOI211_X1 i_0_498 (.ZN (n_0_497), .A (n_0_500), .B (n_0_575), .C1 (n_0_540), .C2 (n_0_499));
AOI22_X1 i_0_497 (.ZN (n_0_496), .A1 (B[20]), .A2 (n_102), .B1 (n_0_601), .B2 (n_0_497));
INV_X1 i_0_496 (.ZN (n_96), .A (n_0_496));
AND3_X1 i_0_495 (.ZN (n_0_494), .A1 (n_0_515), .A2 (n_0_498), .A3 (n_0_600));
NAND2_X1 i_0_494 (.ZN (n_0_491), .A1 (n_0_611), .A2 (n_0_593));
INV_X1 i_0_493 (.ZN (n_0_490), .A (n_0_491));
AOI21_X1 i_0_492 (.ZN (n_0_489), .A (n_0_597), .B1 (B[21]), .B2 (n_0_593));
AOI211_X1 i_0_491 (.ZN (n_0_488), .A (n_0_489), .B (n_0_577), .C1 (n_0_597), .C2 (n_0_490));
AOI221_X1 i_0_490 (.ZN (n_0_487), .A (n_0_494), .B1 (n_0_558), .B2 (n_0_488), .C1 (B[19]), .C2 (n_102));
INV_X1 i_0_489 (.ZN (n_95), .A (n_0_487));
OAI22_X1 i_0_488 (.ZN (n_0_486), .A1 (n_0_610), .A2 (n_0_598), .B1 (n_0_612), .B2 (n_0_597));
NAND2_X1 i_0_487 (.ZN (n_0_485), .A1 (n_0_515), .A2 (n_0_486));
NAND2_X1 i_0_486 (.ZN (n_0_483), .A1 (n_0_597), .A2 (n_0_576));
OAI21_X1 i_0_485 (.ZN (n_0_482), .A (n_0_485), .B1 (n_0_613), .B2 (n_0_483));
AOI222_X1 i_0_484 (.ZN (n_0_481), .A1 (n_0_558), .A2 (n_0_482), .B1 (B[18]), .B2 (n_102)
    , .C1 (n_0_600), .C2 (n_0_488));
INV_X1 i_0_483 (.ZN (n_94), .A (n_0_481));
AOI22_X1 i_0_482 (.ZN (n_0_480), .A1 (B[17]), .A2 (n_0_593), .B1 (B[21]), .B2 (n_0_594));
INV_X1 i_0_481 (.ZN (n_0_479), .A (n_0_480));
AOI221_X1 i_0_480 (.ZN (n_0_478), .A (n_0_577), .B1 (n_0_597), .B2 (n_0_480), .C1 (n_0_598), .C2 (n_0_490));
AOI222_X1 i_0_479 (.ZN (n_0_477), .A1 (n_0_558), .A2 (n_0_478), .B1 (B[17]), .B2 (n_102)
    , .C1 (n_0_600), .C2 (n_0_482));
INV_X1 i_0_478 (.ZN (n_93), .A (n_0_477));
AOI221_X1 i_0_477 (.ZN (n_0_476), .A (n_0_575), .B1 (n_0_608), .B2 (n_0_597), .C1 (n_0_610), .C2 (n_0_598));
AOI21_X1 i_0_476 (.ZN (n_0_475), .A (n_0_476), .B1 (n_0_498), .B2 (n_0_576));
INV_X1 i_0_475 (.ZN (n_0_474), .A (n_0_475));
AOI222_X1 i_0_474 (.ZN (n_0_473), .A1 (n_0_558), .A2 (n_0_474), .B1 (B[16]), .B2 (n_102)
    , .C1 (n_0_600), .C2 (n_0_478));
INV_X1 i_0_473 (.ZN (n_92), .A (n_0_473));
NAND2_X1 i_0_472 (.ZN (n_0_472), .A1 (n_0_598), .A2 (n_0_479));
AOI221_X1 i_0_471 (.ZN (n_0_469), .A (n_0_572), .B1 (B[19]), .B2 (n_0_576), .C1 (B[15]), .C2 (n_0_515));
OAI22_X1 i_0_470 (.ZN (n_0_468), .A1 (n_0_577), .A2 (n_0_472), .B1 (n_0_598), .B2 (n_0_469));
AOI222_X1 i_0_469 (.ZN (n_0_467), .A1 (n_0_600), .A2 (n_0_474), .B1 (B[15]), .B2 (n_102)
    , .C1 (n_0_558), .C2 (n_0_468));
INV_X1 i_0_468 (.ZN (n_91), .A (n_0_467));
AOI22_X1 i_0_467 (.ZN (n_0_466), .A1 (B[14]), .A2 (n_0_589), .B1 (B[22]), .B2 (n_0_573));
OR2_X1 i_0_466 (.ZN (n_0_465), .A1 (n_0_594), .A2 (n_0_466));
NOR3_X1 i_0_465 (.ZN (n_0_464), .A1 (n_0_608), .A2 (n_0_597), .A3 (n_0_575));
AOI21_X1 i_0_464 (.ZN (n_0_463), .A (n_0_464), .B1 (n_0_486), .B2 (n_0_576));
OAI21_X1 i_0_463 (.ZN (n_0_462), .A (n_0_463), .B1 (n_0_598), .B2 (n_0_465));
AOI222_X1 i_0_462 (.ZN (n_0_461), .A1 (B[14]), .A2 (n_102), .B1 (n_0_558), .B2 (n_0_462)
    , .C1 (n_0_600), .C2 (n_0_468));
INV_X1 i_0_460 (.ZN (n_90), .A (n_0_461));
AOI222_X1 i_0_459 (.ZN (n_0_460), .A1 (B[13]), .A2 (n_0_515), .B1 (B[21]), .B2 (n_0_572)
    , .C1 (B[17]), .C2 (n_0_576));
AOI22_X1 i_0_458 (.ZN (n_0_459), .A1 (n_0_597), .A2 (n_0_460), .B1 (n_0_598), .B2 (n_0_469));
AOI222_X1 i_0_457 (.ZN (n_0_458), .A1 (n_0_600), .A2 (n_0_462), .B1 (B[13]), .B2 (n_102)
    , .C1 (n_0_558), .C2 (n_0_459));
INV_X1 i_0_456 (.ZN (n_89), .A (n_0_458));
AOI222_X1 i_0_455 (.ZN (n_0_457), .A1 (B[16]), .A2 (n_0_576), .B1 (B[12]), .B2 (n_0_515)
    , .C1 (B[20]), .C2 (n_0_572));
AOI21_X1 i_0_454 (.ZN (n_0_456), .A (n_0_597), .B1 (B[18]), .B2 (n_0_576));
AOI22_X1 i_0_453 (.ZN (n_0_455), .A1 (n_0_597), .A2 (n_0_457), .B1 (n_0_465), .B2 (n_0_456));
AOI22_X1 i_0_452 (.ZN (n_0_454), .A1 (n_0_600), .A2 (n_0_459), .B1 (n_0_558), .B2 (n_0_455));
OAI21_X1 i_0_451 (.ZN (n_88), .A (n_0_454), .B1 (n_0_606), .B2 (n_0_617));
AOI222_X1 i_0_450 (.ZN (n_0_453), .A1 (B[11]), .A2 (n_0_515), .B1 (n_0_491), .B2 (n_0_573)
    , .C1 (B[15]), .C2 (n_0_576));
AOI22_X1 i_0_449 (.ZN (n_0_452), .A1 (n_0_597), .A2 (n_0_453), .B1 (n_0_598), .B2 (n_0_460));
AOI222_X1 i_0_448 (.ZN (n_0_451), .A1 (n_0_558), .A2 (n_0_452), .B1 (B[11]), .B2 (n_102)
    , .C1 (n_0_600), .C2 (n_0_455));
INV_X1 i_0_447 (.ZN (n_87), .A (n_0_451));
AOI22_X1 i_0_446 (.ZN (n_0_449), .A1 (n_0_594), .A2 (n_0_466), .B1 (n_0_593), .B2 (n_0_567));
INV_X1 i_0_445 (.ZN (n_0_448), .A (n_0_449));
AOI22_X1 i_0_444 (.ZN (n_0_447), .A1 (n_0_598), .A2 (n_0_457), .B1 (n_0_597), .B2 (n_0_448));
AOI222_X1 i_0_443 (.ZN (n_0_446), .A1 (B[10]), .A2 (n_102), .B1 (n_0_600), .B2 (n_0_452)
    , .C1 (n_0_558), .C2 (n_0_447));
INV_X1 i_0_442 (.ZN (n_86), .A (n_0_446));
AOI222_X1 i_0_441 (.ZN (n_0_445), .A1 (B[9]), .A2 (n_0_515), .B1 (n_0_479), .B2 (n_0_573)
    , .C1 (B[13]), .C2 (n_0_576));
AOI22_X1 i_0_440 (.ZN (n_0_444), .A1 (n_0_597), .A2 (n_0_445), .B1 (n_0_598), .B2 (n_0_453));
AOI22_X1 i_0_439 (.ZN (n_0_443), .A1 (n_0_558), .A2 (n_0_444), .B1 (n_0_600), .B2 (n_0_447));
OAI21_X1 i_0_438 (.ZN (n_85), .A (n_0_443), .B1 (n_0_603), .B2 (n_0_617));
AOI22_X1 i_0_437 (.ZN (n_0_438), .A1 (n_0_597), .A2 (n_0_568), .B1 (n_0_598), .B2 (n_0_448));
AOI222_X1 i_0_436 (.ZN (n_0_437), .A1 (n_0_558), .A2 (n_0_438), .B1 (B[8]), .B2 (n_102)
    , .C1 (n_0_600), .C2 (n_0_444));
INV_X1 i_0_435 (.ZN (n_84), .A (n_0_437));
AOI22_X1 i_0_434 (.ZN (n_0_432), .A1 (n_0_597), .A2 (n_0_552), .B1 (n_0_598), .B2 (n_0_445));
AOI222_X1 i_0_433 (.ZN (n_0_431), .A1 (n_0_558), .A2 (n_0_432), .B1 (B[7]), .B2 (n_102)
    , .C1 (n_0_600), .C2 (n_0_438));
INV_X1 i_0_432 (.ZN (n_83), .A (n_0_431));
AOI222_X1 i_0_431 (.ZN (n_0_426), .A1 (n_0_600), .A2 (n_0_432), .B1 (B[6]), .B2 (n_102)
    , .C1 (n_0_558), .C2 (n_0_560));
INV_X1 i_0_430 (.ZN (n_82), .A (n_0_426));
AOI22_X1 i_0_429 (.ZN (n_0_420), .A1 (B[12]), .A2 (n_0_573), .B1 (B[20]), .B2 (n_0_566));
OAI21_X1 i_0_428 (.ZN (n_0_419), .A (n_0_420), .B1 (n_0_201), .B2 (n_0_577));
AOI222_X1 i_0_427 (.ZN (n_0_418), .A1 (B[16]), .A2 (n_0_571), .B1 (B[8]), .B2 (n_0_576)
    , .C1 (n_0_593), .C2 (n_0_419));
AOI22_X1 i_0_426 (.ZN (n_0_417), .A1 (n_0_597), .A2 (n_0_418), .B1 (n_0_598), .B2 (n_0_561));
AOI222_X1 i_0_425 (.ZN (n_0_416), .A1 (n_0_558), .A2 (n_0_417), .B1 (B[4]), .B2 (n_102)
    , .C1 (n_0_600), .C2 (n_0_551));
INV_X1 i_0_424 (.ZN (n_81), .A (n_0_416));
NAND2_X1 i_0_423 (.ZN (n_0_415), .A1 (B[11]), .A2 (n_0_572));
NOR3_X1 i_0_422 (.ZN (n_0_414), .A1 (n_0_592), .A2 (n_0_590), .A3 (n_0_594));
OAI21_X1 i_0_421 (.ZN (n_0_413), .A (n_0_415), .B1 (n_0_202), .B2 (n_0_575));
AOI221_X1 i_0_420 (.ZN (n_0_412), .A (n_0_413), .B1 (n_0_594), .B2 (n_0_553), .C1 (B[19]), .C2 (n_0_414));
AOI22_X1 i_0_419 (.ZN (n_0_411), .A1 (n_0_597), .A2 (n_0_412), .B1 (n_0_598), .B2 (n_0_555));
AOI22_X1 i_0_418 (.ZN (n_0_410), .A1 (n_0_600), .A2 (n_0_417), .B1 (n_0_558), .B2 (n_0_411));
OAI21_X1 i_0_417 (.ZN (n_80), .A (n_0_410), .B1 (n_0_202), .B2 (n_0_617));
OAI22_X1 i_0_416 (.ZN (n_0_409), .A1 (n_0_593), .A2 (n_0_565), .B1 (n_0_199), .B2 (n_0_575));
AOI221_X1 i_0_415 (.ZN (n_0_408), .A (n_0_409), .B1 (B[10]), .B2 (n_0_572), .C1 (B[18]), .C2 (n_0_414));
AOI22_X1 i_0_414 (.ZN (n_0_407), .A1 (n_0_597), .A2 (n_0_408), .B1 (n_0_598), .B2 (n_0_418));
AOI222_X1 i_0_413 (.ZN (n_0_406), .A1 (B[2]), .A2 (n_102), .B1 (n_0_600), .B2 (n_0_411)
    , .C1 (n_0_558), .C2 (n_0_407));
INV_X1 i_0_412 (.ZN (n_79), .A (n_0_406));
AOI22_X1 i_0_411 (.ZN (n_0_405), .A1 (n_0_594), .A2 (n_0_556), .B1 (B[9]), .B2 (n_0_572));
INV_X1 i_0_410 (.ZN (n_0_404), .A (n_0_405));
AOI221_X1 i_0_409 (.ZN (n_0_403), .A (n_0_404), .B1 (B[17]), .B2 (n_0_414), .C1 (B[1]), .C2 (n_0_515));
AOI22_X1 i_0_408 (.ZN (n_0_402), .A1 (n_0_598), .A2 (n_0_412), .B1 (n_0_597), .B2 (n_0_403));
AOI22_X1 i_0_407 (.ZN (n_0_401), .A1 (n_0_558), .A2 (n_0_402), .B1 (n_0_600), .B2 (n_0_407));
OAI21_X1 i_0_406 (.ZN (n_78), .A (n_0_401), .B1 (n_0_200), .B2 (n_0_617));
AOI21_X1 i_0_405 (.ZN (n_0_400), .A (n_0_598), .B1 (B[16]), .B2 (n_0_414));
AOI222_X1 i_0_404 (.ZN (n_0_399), .A1 (B[8]), .A2 (n_0_572), .B1 (B[0]), .B2 (n_0_515)
    , .C1 (n_0_594), .C2 (n_0_419));
AOI221_X1 i_0_403 (.ZN (n_0_398), .A (n_0_559), .B1 (n_0_400), .B2 (n_0_399), .C1 (n_0_510), .C2 (n_0_408));
AOI221_X1 i_0_402 (.ZN (n_0_397), .A (n_0_398), .B1 (B[0]), .B2 (n_102), .C1 (n_0_600), .C2 (n_0_402));
INV_X1 i_0_401 (.ZN (n_77), .A (n_0_397));
INV_X1 i_0_400 (.ZN (n_0_396), .A (n_100));
AND2_X1 i_0_399 (.ZN (n_0_382), .A1 (n_0_422), .A2 (n_0_492));
AOI22_X1 i_0_398 (.ZN (n_0_381), .A1 (A[22]), .A2 (n_100), .B1 (drc_ipo_n4), .B2 (n_0_382));
INV_X1 i_0_461 (.ZN (n_76), .A (n_0_381));
AOI21_X1 i_0_397 (.ZN (n_0_380), .A (n_0_597), .B1 (n_0_588), .B2 (n_0_599));
AOI22_X1 i_0_396 (.ZN (n_0_379), .A1 (A[21]), .A2 (n_100), .B1 (n_0_382), .B2 (n_0_380));
INV_X1 i_0_395 (.ZN (n_75), .A (n_0_379));
AOI21_X1 i_0_394 (.ZN (n_0_378), .A (n_0_539), .B1 (A[22]), .B2 (n_0_450));
AOI21_X1 i_0_393 (.ZN (n_0_377), .A (n_0_378), .B1 (n_0_587), .B2 (drc_ipo_n4));
AOI22_X1 i_0_392 (.ZN (n_0_376), .A1 (A[20]), .A2 (n_100), .B1 (n_0_382), .B2 (n_0_377));
INV_X1 i_0_391 (.ZN (n_74), .A (n_0_376));
NAND2_X1 i_0_390 (.ZN (n_0_373), .A1 (n_0_450), .A2 (n_0_422));
NOR2_X1 i_0_389 (.ZN (n_0_372), .A1 (A[19]), .A2 (n_0_441));
OAI33_X1 i_0_388 (.ZN (n_0_371), .A1 (drc_ipo_n4), .A2 (n_0_421), .A3 (n_0_587), .B1 (n_0_430)
    , .B2 (n_0_372), .B3 (n_0_450));
OAI22_X1 i_0_387 (.ZN (n_0_370), .A1 (n_0_588), .A2 (drc_ipo_n4), .B1 (n_0_586), .B2 (n_0_450));
AND3_X1 i_0_386 (.ZN (n_0_368), .A1 (n_0_422), .A2 (n_0_370), .A3 (n_0_390));
AOI221_X1 i_0_385 (.ZN (n_0_367), .A (n_0_368), .B1 (n_0_484), .B2 (n_0_371), .C1 (A[19]), .C2 (n_100));
INV_X1 i_0_384 (.ZN (n_73), .A (n_0_367));
AOI22_X1 i_0_383 (.ZN (n_0_365), .A1 (A[18]), .A2 (n_0_422), .B1 (A[22]), .B2 (n_0_394));
OAI22_X1 i_0_382 (.ZN (n_0_364), .A1 (n_0_586), .A2 (n_0_373), .B1 (n_0_450), .B2 (n_0_365));
AOI222_X1 i_0_381 (.ZN (n_0_363), .A1 (A[18]), .A2 (n_100), .B1 (n_0_371), .B2 (n_0_390)
    , .C1 (n_0_484), .C2 (n_0_364));
INV_X1 i_0_380 (.ZN (n_72), .A (n_0_363));
AOI221_X1 i_0_379 (.ZN (n_0_360), .A (n_0_430), .B1 (drc_ipo_n4), .B2 (n_0_395), .C1 (n_0_450), .C2 (n_0_372));
AOI222_X1 i_0_378 (.ZN (n_0_359), .A1 (n_0_484), .A2 (n_0_360), .B1 (A[17]), .B2 (n_100)
    , .C1 (n_0_390), .C2 (n_0_364));
INV_X1 i_0_377 (.ZN (n_71), .A (n_0_359));
AOI22_X1 i_0_376 (.ZN (n_0_358), .A1 (A[16]), .A2 (n_0_422), .B1 (A[20]), .B2 (n_0_394));
AOI22_X1 i_0_375 (.ZN (n_0_357), .A1 (n_0_450), .A2 (n_0_365), .B1 (drc_ipo_n4), .B2 (n_0_358));
AOI222_X1 i_0_374 (.ZN (n_0_356), .A1 (n_0_390), .A2 (n_0_360), .B1 (A[16]), .B2 (n_100)
    , .C1 (n_0_484), .C2 (n_0_357));
INV_X1 i_0_373 (.ZN (n_70), .A (n_0_356));
NAND2_X1 i_0_372 (.ZN (n_0_355), .A1 (A[19]), .A2 (n_0_394));
AND2_X1 i_0_371 (.ZN (n_0_351), .A1 (n_0_434), .A2 (n_0_425));
OAI21_X1 i_0_370 (.ZN (n_0_350), .A (n_0_355), .B1 (n_0_441), .B2 (n_0_351));
NOR3_X1 i_0_369 (.ZN (n_0_349), .A1 (n_0_430), .A2 (n_0_395), .A3 (drc_ipo_n4));
AOI21_X1 i_0_368 (.ZN (n_0_348), .A (n_0_349), .B1 (drc_ipo_n4), .B2 (n_0_350));
INV_X1 i_0_367 (.ZN (n_0_347), .A (n_0_348));
AOI222_X1 i_0_366 (.ZN (n_0_346), .A1 (n_0_484), .A2 (n_0_347), .B1 (A[15]), .B2 (n_100)
    , .C1 (n_0_390), .C2 (n_0_357));
INV_X1 i_0_365 (.ZN (n_69), .A (n_0_346));
AOI222_X1 i_0_364 (.ZN (n_0_344), .A1 (A[22]), .A2 (n_0_388), .B1 (A[14]), .B2 (n_0_422)
    , .C1 (A[18]), .C2 (n_0_394));
AOI22_X1 i_0_363 (.ZN (n_0_343), .A1 (n_0_450), .A2 (n_0_358), .B1 (drc_ipo_n4), .B2 (n_0_344));
AOI222_X1 i_0_362 (.ZN (n_0_342), .A1 (A[14]), .A2 (n_100), .B1 (n_0_390), .B2 (n_0_347)
    , .C1 (n_0_484), .C2 (n_0_343));
INV_X1 i_0_361 (.ZN (n_68), .A (n_0_342));
AOI22_X1 i_0_360 (.ZN (n_0_341), .A1 (A[21]), .A2 (n_0_388), .B1 (A[17]), .B2 (n_0_394));
OAI21_X1 i_0_359 (.ZN (n_0_340), .A (n_0_341), .B1 (n_0_579), .B2 (n_0_421));
AOI22_X1 i_0_358 (.ZN (n_0_339), .A1 (n_0_450), .A2 (n_0_350), .B1 (drc_ipo_n4), .B2 (n_0_340));
INV_X1 i_0_357 (.ZN (n_0_338), .A (n_0_339));
AOI222_X1 i_0_356 (.ZN (n_0_337), .A1 (n_0_390), .A2 (n_0_343), .B1 (A[13]), .B2 (n_100)
    , .C1 (n_0_484), .C2 (n_0_338));
INV_X1 i_0_355 (.ZN (n_67), .A (n_0_337));
AOI222_X1 i_0_354 (.ZN (n_0_336), .A1 (A[16]), .A2 (n_0_394), .B1 (A[12]), .B2 (n_0_422)
    , .C1 (A[20]), .C2 (n_0_388));
AOI22_X1 i_0_353 (.ZN (n_0_335), .A1 (drc_ipo_n4), .A2 (n_0_336), .B1 (n_0_450), .B2 (n_0_344));
AOI222_X1 i_0_352 (.ZN (n_0_334), .A1 (n_0_390), .A2 (n_0_338), .B1 (A[12]), .B2 (n_100)
    , .C1 (n_0_484), .C2 (n_0_335));
INV_X1 i_0_351 (.ZN (n_66), .A (n_0_334));
AOI22_X1 i_0_350 (.ZN (n_0_332), .A1 (n_0_442), .A2 (n_0_428), .B1 (n_0_441), .B2 (n_0_351));
INV_X1 i_0_349 (.ZN (n_0_331), .A (n_0_332));
NAND2_X1 i_0_348 (.ZN (n_0_330), .A1 (n_0_450), .A2 (n_0_340));
OAI21_X1 i_0_347 (.ZN (n_0_329), .A (n_0_330), .B1 (n_0_450), .B2 (n_0_331));
AOI222_X1 i_0_346 (.ZN (n_0_328), .A1 (n_0_484), .A2 (n_0_329), .B1 (A[11]), .B2 (n_100)
    , .C1 (n_0_390), .C2 (n_0_335));
INV_X1 i_0_344 (.ZN (n_65), .A (n_0_328));
NOR2_X1 i_0_343 (.ZN (n_0_322), .A1 (n_0_450), .A2 (n_0_384));
AOI21_X1 i_0_342 (.ZN (n_0_321), .A (n_0_322), .B1 (n_0_450), .B2 (n_0_336));
AOI222_X1 i_0_341 (.ZN (n_0_320), .A1 (n_0_390), .A2 (n_0_329), .B1 (A[10]), .B2 (n_100)
    , .C1 (n_0_484), .C2 (n_0_321));
INV_X1 i_0_340 (.ZN (n_64), .A (n_0_320));
AOI22_X1 i_0_339 (.ZN (n_0_318), .A1 (drc_ipo_n4), .A2 (n_0_392), .B1 (n_0_450), .B2 (n_0_331));
AOI222_X1 i_0_338 (.ZN (n_0_317), .A1 (n_0_390), .A2 (n_0_321), .B1 (A[9]), .B2 (n_100)
    , .C1 (n_0_484), .C2 (n_0_318));
INV_X1 i_0_337 (.ZN (n_63), .A (n_0_317));
AOI222_X1 i_0_336 (.ZN (n_0_311), .A1 (n_0_390), .A2 (n_0_318), .B1 (A[8]), .B2 (n_100)
    , .C1 (n_0_484), .C2 (n_0_369));
INV_X1 i_0_335 (.ZN (n_62), .A (n_0_311));
NOR2_X1 i_0_334 (.ZN (n_0_305), .A1 (n_0_439), .A2 (n_0_435));
AOI22_X1 i_0_332 (.ZN (n_0_304), .A1 (A[14]), .A2 (n_0_433), .B1 (A[22]), .B2 (n_0_305));
OAI21_X1 i_0_331 (.ZN (n_0_303), .A (n_0_304), .B1 (n_0_309), .B2 (n_0_430));
AOI222_X1 i_0_330 (.ZN (n_0_302), .A1 (A[18]), .A2 (n_0_389), .B1 (A[10]), .B2 (n_0_394)
    , .C1 (n_0_442), .C2 (n_0_303));
AOI22_X1 i_0_329 (.ZN (n_0_301), .A1 (drc_ipo_n4), .A2 (n_0_302), .B1 (n_0_450), .B2 (n_0_374));
AOI222_X1 i_0_328 (.ZN (n_0_300), .A1 (A[6]), .A2 (n_100), .B1 (n_0_390), .B2 (n_0_391)
    , .C1 (n_0_484), .C2 (n_0_301));
INV_X1 i_0_327 (.ZN (n_61), .A (n_0_300));
AOI22_X1 i_0_326 (.ZN (n_0_299), .A1 (A[13]), .A2 (n_0_433), .B1 (A[21]), .B2 (n_0_305));
OAI21_X1 i_0_325 (.ZN (n_0_298), .A (n_0_299), .B1 (n_0_307), .B2 (n_0_430));
AOI222_X1 i_0_324 (.ZN (n_0_297), .A1 (A[17]), .A2 (n_0_389), .B1 (A[9]), .B2 (n_0_394)
    , .C1 (n_0_442), .C2 (n_0_298));
AOI22_X1 i_0_323 (.ZN (n_0_296), .A1 (drc_ipo_n4), .A2 (n_0_297), .B1 (n_0_450), .B2 (n_0_423));
AOI222_X1 i_0_322 (.ZN (n_0_295), .A1 (n_0_390), .A2 (n_0_301), .B1 (A[5]), .B2 (n_100)
    , .C1 (n_0_484), .C2 (n_0_296));
INV_X1 i_0_321 (.ZN (n_60), .A (n_0_295));
AOI22_X1 i_0_320 (.ZN (n_0_294), .A1 (A[12]), .A2 (n_0_433), .B1 (A[20]), .B2 (n_0_305));
OAI21_X1 i_0_319 (.ZN (n_0_293), .A (n_0_294), .B1 (n_0_306), .B2 (n_0_430));
AOI222_X1 i_0_318 (.ZN (n_0_292), .A1 (A[16]), .A2 (n_0_389), .B1 (A[8]), .B2 (n_0_394)
    , .C1 (n_0_442), .C2 (n_0_293));
AOI22_X1 i_0_317 (.ZN (n_0_291), .A1 (drc_ipo_n4), .A2 (n_0_292), .B1 (n_0_450), .B2 (n_0_302));
AOI222_X1 i_0_316 (.ZN (n_0_290), .A1 (n_0_390), .A2 (n_0_296), .B1 (A[4]), .B2 (n_100)
    , .C1 (n_0_484), .C2 (n_0_291));
INV_X1 i_0_315 (.ZN (n_59), .A (n_0_290));
NOR3_X1 i_0_314 (.ZN (n_0_289), .A1 (n_0_439), .A2 (n_0_435), .A3 (n_0_441));
AOI22_X1 i_0_313 (.ZN (n_0_288), .A1 (n_0_441), .A2 (n_0_424), .B1 (A[11]), .B2 (n_0_388));
INV_X1 i_0_312 (.ZN (n_0_287), .A (n_0_288));
AOI221_X1 i_0_311 (.ZN (n_0_286), .A (n_0_287), .B1 (A[19]), .B2 (n_0_289), .C1 (A[3]), .C2 (n_0_422));
AOI22_X1 i_0_310 (.ZN (n_0_285), .A1 (drc_ipo_n4), .A2 (n_0_286), .B1 (n_0_450), .B2 (n_0_297));
AOI222_X2 i_0_309 (.ZN (n_0_284), .A1 (n_0_390), .A2 (n_0_291), .B1 (A[3]), .B2 (n_100)
    , .C1 (n_0_484), .C2 (n_0_285));
INV_X1 i_0_345 (.ZN (n_58), .A (n_0_284));
AOI22_X1 i_0_308 (.ZN (n_0_283), .A1 (n_0_441), .A2 (n_0_303), .B1 (A[10]), .B2 (n_0_388));
INV_X1 i_0_307 (.ZN (n_0_282), .A (n_0_283));
AOI221_X1 i_0_306 (.ZN (n_0_281), .A (n_0_282), .B1 (A[18]), .B2 (n_0_289), .C1 (A[2]), .C2 (n_0_422));
AOI22_X1 i_0_305 (.ZN (n_0_280), .A1 (drc_ipo_n4), .A2 (n_0_281), .B1 (n_0_450), .B2 (n_0_292));
AOI222_X2 i_0_304 (.ZN (n_0_279), .A1 (n_0_484), .A2 (n_0_280), .B1 (A[2]), .B2 (n_100)
    , .C1 (n_0_390), .C2 (n_0_285));
INV_X1 i_0_303 (.ZN (n_57), .A (n_0_279));
NAND2_X1 i_0_302 (.ZN (n_0_278), .A1 (A[9]), .A2 (n_0_388));
OAI21_X1 i_0_301 (.ZN (n_0_277), .A (n_0_278), .B1 (n_0_198), .B2 (n_0_421));
AOI221_X1 i_0_300 (.ZN (n_0_276), .A (n_0_277), .B1 (A[17]), .B2 (n_0_289), .C1 (n_0_441), .C2 (n_0_298));
AOI22_X1 i_0_299 (.ZN (n_0_275), .A1 (n_0_450), .A2 (n_0_286), .B1 (drc_ipo_n4), .B2 (n_0_276));
AOI222_X2 i_0_298 (.ZN (n_0_274), .A1 (n_0_390), .A2 (n_0_280), .B1 (A[1]), .B2 (n_100)
    , .C1 (n_0_484), .C2 (n_0_275));
INV_X1 i_0_333 (.ZN (n_56), .A (n_0_274));
AOI22_X1 i_0_297 (.ZN (n_0_273), .A1 (n_0_441), .A2 (n_0_293), .B1 (A[0]), .B2 (n_0_422));
INV_X1 i_0_296 (.ZN (n_0_272), .A (n_0_273));
AOI221_X1 i_0_295 (.ZN (n_0_271), .A (n_0_272), .B1 (A[8]), .B2 (n_0_388), .C1 (A[16]), .C2 (n_0_289));
AOI221_X1 i_0_294 (.ZN (n_0_270), .A (n_0_471), .B1 (drc_ipo_n4), .B2 (n_0_271), .C1 (n_0_450), .C2 (n_0_281));
AOI221_X1 i_0_293 (.ZN (n_0_269), .A (n_0_270), .B1 (A[0]), .B2 (n_100), .C1 (n_0_390), .C2 (n_0_275));
INV_X1 i_0_292 (.ZN (n_55), .A (n_0_269));
AOI22_X1 i_0_291 (.ZN (n_0_268), .A1 (B[29]), .A2 (n_0_396), .B1 (A[29]), .B2 (n_100));
INV_X1 i_0_290 (.ZN (\exp_Sum[6] ), .A (n_0_268));
AOI22_X1 i_0_289 (.ZN (n_0_267), .A1 (B[28]), .A2 (n_0_396), .B1 (A[28]), .B2 (n_100));
INV_X1 i_0_288 (.ZN (\exp_Sum[5] ), .A (n_0_267));
AOI22_X1 i_0_287 (.ZN (n_0_266), .A1 (B[27]), .A2 (n_0_396), .B1 (A[27]), .B2 (n_100));
INV_X1 i_0_286 (.ZN (\exp_Sum[4] ), .A (n_0_266));
AOI22_X1 i_0_285 (.ZN (n_0_265), .A1 (B[26]), .A2 (n_0_396), .B1 (A[26]), .B2 (n_100));
INV_X1 i_0_284 (.ZN (\exp_Sum[3] ), .A (n_0_265));
AOI22_X1 i_0_283 (.ZN (n_0_264), .A1 (B[25]), .A2 (n_0_396), .B1 (A[25]), .B2 (n_100));
INV_X1 i_0_282 (.ZN (\exp_Sum[2] ), .A (n_0_264));
AOI22_X1 i_0_281 (.ZN (n_0_263), .A1 (B[24]), .A2 (n_0_396), .B1 (A[24]), .B2 (n_100));
INV_X1 i_0_280 (.ZN (\exp_Sum[1] ), .A (n_0_263));
AOI22_X1 i_0_279 (.ZN (n_0_262), .A1 (B[23]), .A2 (n_0_396), .B1 (A[23]), .B2 (n_100));
INV_X1 i_0_277 (.ZN (\exp_Sum[0] ), .A (n_0_262));
NAND2_X1 i_0_276 (.ZN (n_0_261), .A1 (n_78), .A2 (n_0_274));
XOR2_X1 i_0_275 (.Z (n_0_260), .A (n_88), .B (n_66));
NOR2_X1 i_0_274 (.ZN (n_0_259), .A1 (n_85), .A2 (n_0_317));
AOI222_X1 i_0_273 (.ZN (n_0_258), .A1 (n_0_501), .A2 (n_75), .B1 (n_0_496), .B2 (n_74)
    , .C1 (n_97), .C2 (n_0_379));
XOR2_X1 i_0_272 (.Z (n_0_257), .A (n_98), .B (n_0_381));
AOI211_X1 i_0_271 (.ZN (n_0_256), .A (n_0_506), .B (n_0_517), .C1 (n_96), .C2 (n_0_376));
NAND3_X1 i_0_270 (.ZN (n_0_255), .A1 (n_0_257), .A2 (n_0_256), .A3 (n_0_258));
AOI22_X1 i_0_269 (.ZN (n_0_254), .A1 (n_0_451), .A2 (n_65), .B1 (n_87), .B2 (n_0_328));
OAI22_X1 i_0_268 (.ZN (n_0_253), .A1 (n_0_431), .A2 (n_0_366), .B1 (n_83), .B2 (n_99));
AOI22_X1 i_0_267 (.ZN (n_0_252), .A1 (n_82), .A2 (n_0_300), .B1 (n_0_446), .B2 (n_64));
AOI222_X1 i_0_266 (.ZN (n_0_251), .A1 (n_93), .A2 (n_0_359), .B1 (n_92), .B2 (n_0_356)
    , .C1 (n_0_426), .C2 (n_61));
OAI221_X1 i_0_265 (.ZN (n_0_250), .A (n_0_251), .B1 (n_0_487), .B2 (n_73), .C1 (n_95), .C2 (n_0_367));
AOI221_X1 i_0_264 (.ZN (n_0_249), .A (n_0_250), .B1 (n_86), .B2 (n_0_320), .C1 (n_0_437), .C2 (n_62));
OAI211_X1 i_0_263 (.ZN (n_0_248), .A (n_0_252), .B (n_0_249), .C1 (n_0_437), .C2 (n_62));
AOI221_X1 i_0_262 (.ZN (n_0_247), .A (n_0_248), .B1 (n_0_550), .B2 (n_60), .C1 (n_101), .C2 (n_0_295));
OAI221_X1 i_0_261 (.ZN (n_0_246), .A (n_0_247), .B1 (n_0_397), .B2 (n_55), .C1 (n_77), .C2 (n_0_269));
OAI221_X1 i_0_260 (.ZN (n_0_245), .A (n_0_254), .B1 (n_79), .B2 (n_0_279), .C1 (n_78), .C2 (n_0_274));
OAI21_X1 i_0_259 (.ZN (n_0_244), .A (n_0_261), .B1 (n_81), .B2 (n_0_290));
AOI22_X1 i_0_258 (.ZN (n_0_243), .A1 (n_94), .A2 (n_0_363), .B1 (n_0_481), .B2 (n_72));
AOI22_X1 i_0_257 (.ZN (n_0_242), .A1 (n_91), .A2 (n_0_346), .B1 (n_90), .B2 (n_0_342));
AOI221_X1 i_0_256 (.ZN (n_0_241), .A (n_0_255), .B1 (n_0_477), .B2 (n_71), .C1 (n_0_473), .C2 (n_70));
AOI22_X1 i_0_255 (.ZN (n_0_240), .A1 (n_0_467), .A2 (n_69), .B1 (n_0_461), .B2 (n_68));
NAND4_X1 i_0_254 (.ZN (n_0_239), .A1 (n_0_243), .A2 (n_0_242), .A3 (n_0_241), .A4 (n_0_240));
NOR4_X1 i_0_253 (.ZN (n_0_238), .A1 (n_0_260), .A2 (n_0_245), .A3 (n_0_244), .A4 (n_0_239));
OAI222_X1 i_0_252 (.ZN (n_0_237), .A1 (n_80), .A2 (n_0_284), .B1 (n_0_406), .B2 (n_57)
    , .C1 (n_0_416), .C2 (n_59));
AOI221_X1 i_0_251 (.ZN (n_0_236), .A (n_0_237), .B1 (n_0_458), .B2 (n_67), .C1 (n_89), .C2 (n_0_337));
AOI221_X1 i_0_250 (.ZN (n_0_235), .A (n_0_259), .B1 (n_85), .B2 (n_0_317), .C1 (n_80), .C2 (n_0_284));
NAND4_X1 i_0_249 (.ZN (n_0_234), .A1 (n_0_253), .A2 (n_0_235), .A3 (n_0_236), .A4 (n_0_238));
XNOR2_X1 i_0_248 (.ZN (n_0_233), .A (n_0_94), .B (A[31]));
INV_X1 i_0_247 (.ZN (n_0_232), .A (n_0_233));
OAI21_X4 i_0_246 (.ZN (n_0_231), .A (n_0_233), .B1 (n_0_246), .B2 (n_0_234));
INV_X1 i_0_245 (.ZN (n_0_230), .A (n_0_231));
AOI21_X1 i_0_244 (.ZN (n_0_229), .A (n_0_231), .B1 (\num_leading_zeros[4] ), .B2 (\num_leading_zeros[3] ));
INV_X1 i_0_243 (.ZN (n_0_228), .A (n_0_229));
AND2_X1 i_0_278 (.ZN (underflow), .A1 (n_25), .A2 (n_0_229));
NAND3_X1 i_0_242 (.ZN (n_0_227), .A1 (\exp_Sum[3] ), .A2 (\exp_Sum[2] ), .A3 (\exp_Sum[1] ));
NOR4_X1 i_0_241 (.ZN (n_0_226), .A1 (\exp_Sum[0] ), .A2 (n_0_227), .A3 (n_0_267), .A4 (n_0_266));
NAND4_X1 i_0_240 (.ZN (n_0_225), .A1 (n_24), .A2 (\exp_Sum[7] ), .A3 (\exp_Sum[6] ), .A4 (n_0_226));
NOR2_X1 i_0_239 (.ZN (overflow), .A1 (n_0_233), .A2 (n_0_225));
AND2_X1 i_0_238 (.ZN (\mant_A[31] ), .A1 (n_54), .A2 (n_0_230));
AOI22_X1 i_0_237 (.ZN (\mant_A[23] ), .A1 (n_0_564), .A2 (n_0_230), .B1 (n_0_396), .B2 (n_0_232));
NOR2_X1 i_0_236 (.ZN (n_0_224), .A1 (n_52), .A2 (n_0_231));
AOI21_X1 i_0_235 (.ZN (\mant_A[22] ), .A (n_0_224), .B1 (n_0_381), .B2 (n_0_231));
NOR2_X1 i_0_234 (.ZN (n_0_223), .A1 (n_51), .A2 (n_0_231));
AOI21_X1 i_0_233 (.ZN (\mant_A[21] ), .A (n_0_223), .B1 (n_0_379), .B2 (n_0_231));
NOR2_X1 i_0_232 (.ZN (n_0_222), .A1 (n_50), .A2 (n_0_231));
AOI21_X1 i_0_231 (.ZN (\mant_A[20] ), .A (n_0_222), .B1 (n_0_376), .B2 (n_0_231));
NOR2_X1 i_0_230 (.ZN (n_0_221), .A1 (n_49), .A2 (n_0_231));
AOI21_X1 i_0_229 (.ZN (\mant_A[19] ), .A (n_0_221), .B1 (n_0_367), .B2 (n_0_231));
NOR2_X1 i_0_228 (.ZN (n_0_220), .A1 (n_48), .A2 (n_0_231));
AOI21_X1 i_0_227 (.ZN (\mant_A[18] ), .A (n_0_220), .B1 (n_0_363), .B2 (n_0_231));
NOR2_X1 i_0_226 (.ZN (n_0_219), .A1 (n_47), .A2 (n_0_231));
AOI21_X1 i_0_225 (.ZN (\mant_A[17] ), .A (n_0_219), .B1 (n_0_359), .B2 (n_0_231));
NOR2_X1 i_0_224 (.ZN (n_0_218), .A1 (n_46), .A2 (n_0_231));
AOI21_X1 i_0_223 (.ZN (\mant_A[16] ), .A (n_0_218), .B1 (n_0_356), .B2 (n_0_231));
NOR2_X1 i_0_222 (.ZN (n_0_217), .A1 (n_45), .A2 (n_0_231));
AOI21_X1 i_0_221 (.ZN (\mant_A[15] ), .A (n_0_217), .B1 (n_0_346), .B2 (n_0_231));
NOR2_X1 i_0_220 (.ZN (n_0_216), .A1 (n_44), .A2 (n_0_231));
AOI21_X1 i_0_219 (.ZN (\mant_A[14] ), .A (n_0_216), .B1 (n_0_342), .B2 (n_0_231));
NOR2_X1 i_0_218 (.ZN (n_0_215), .A1 (n_43), .A2 (n_0_231));
AOI21_X1 i_0_217 (.ZN (\mant_A[13] ), .A (n_0_215), .B1 (n_0_337), .B2 (n_0_231));
NOR2_X1 i_0_195 (.ZN (n_0_214), .A1 (n_42), .A2 (n_0_231));
AOI21_X1 i_0_194 (.ZN (\mant_A[12] ), .A (n_0_214), .B1 (n_0_334), .B2 (n_0_231));
NOR2_X1 i_0_193 (.ZN (n_0_213), .A1 (n_41), .A2 (n_0_231));
AOI21_X1 i_0_192 (.ZN (\mant_A[11] ), .A (n_0_213), .B1 (n_0_328), .B2 (n_0_231));
NOR2_X1 i_0_191 (.ZN (n_0_212), .A1 (n_40), .A2 (n_0_231));
AOI21_X1 i_0_190 (.ZN (\mant_A[10] ), .A (n_0_212), .B1 (n_0_320), .B2 (n_0_231));
NOR2_X1 i_0_189 (.ZN (n_0_211), .A1 (n_39), .A2 (n_0_231));
AOI21_X1 i_0_188 (.ZN (\mant_A[9] ), .A (n_0_211), .B1 (n_0_317), .B2 (n_0_231));
NOR2_X1 i_0_187 (.ZN (n_0_210), .A1 (n_38), .A2 (n_0_231));
AOI21_X1 i_0_186 (.ZN (\mant_A[8] ), .A (n_0_210), .B1 (n_0_311), .B2 (n_0_231));
NOR2_X1 i_0_185 (.ZN (n_0_209), .A1 (n_37), .A2 (n_0_231));
AOI21_X1 i_0_184 (.ZN (\mant_A[7] ), .A (n_0_209), .B1 (n_0_366), .B2 (n_0_231));
NOR2_X1 i_0_183 (.ZN (n_0_208), .A1 (n_36), .A2 (n_0_231));
AOI21_X1 i_0_182 (.ZN (\mant_A[6] ), .A (n_0_208), .B1 (n_0_300), .B2 (n_0_231));
NOR2_X1 i_0_181 (.ZN (n_0_207), .A1 (n_35), .A2 (n_0_231));
AOI21_X1 i_0_180 (.ZN (\mant_A[5] ), .A (n_0_207), .B1 (n_0_295), .B2 (n_0_231));
NOR2_X1 i_0_179 (.ZN (n_0_206), .A1 (n_34), .A2 (n_0_231));
AOI21_X1 i_0_178 (.ZN (\mant_A[4] ), .A (n_0_206), .B1 (n_0_290), .B2 (n_0_231));
NOR2_X1 i_0_177 (.ZN (n_0_205), .A1 (n_33), .A2 (n_0_231));
AOI21_X1 i_0_176 (.ZN (\mant_A[3] ), .A (n_0_205), .B1 (n_0_284), .B2 (n_0_231));
NOR2_X1 i_0_175 (.ZN (n_0_204), .A1 (n_32), .A2 (n_0_231));
AOI21_X1 i_0_174 (.ZN (\mant_A[2] ), .A (n_0_204), .B1 (n_0_279), .B2 (n_0_231));
NOR2_X1 i_0_173 (.ZN (n_0_203), .A1 (n_31), .A2 (n_0_231));
AOI21_X1 i_0_172 (.ZN (\mant_A[1] ), .A (n_0_203), .B1 (n_0_274), .B2 (n_0_231));
AOI221_X1 i_0_216 (.ZN (n_0_191), .A (n_0_362), .B1 (n_0_603), .B2 (A[9]), .C1 (n_0_604), .C2 (A[10]));
INV_X1 i_0_215 (.ZN (n_0_190), .A (n_0_191));
OAI221_X1 i_0_214 (.ZN (n_0_189), .A (n_0_190), .B1 (n_0_604), .B2 (A[10]), .C1 (n_0_605), .C2 (A[11]));
AOI22_X1 i_0_213 (.ZN (n_0_188), .A1 (n_0_606), .A2 (A[12]), .B1 (n_0_605), .B2 (A[11]));
AOI22_X1 i_0_212 (.ZN (n_0_187), .A1 (n_0_189), .A2 (n_0_188), .B1 (B[12]), .B2 (n_0_578));
AOI21_X1 i_0_211 (.ZN (n_0_186), .A (n_0_187), .B1 (n_0_607), .B2 (A[13]));
AOI221_X1 i_0_210 (.ZN (n_0_185), .A (n_0_186), .B1 (B[13]), .B2 (n_0_579), .C1 (B[14]), .C2 (n_0_580));
INV_X1 i_0_209 (.ZN (n_0_184), .A (n_0_185));
OAI221_X1 i_0_208 (.ZN (n_0_183), .A (n_0_184), .B1 (B[14]), .B2 (n_0_580), .C1 (B[15]), .C2 (n_0_581));
AOI22_X1 i_0_207 (.ZN (n_0_182), .A1 (B[16]), .A2 (n_0_582), .B1 (B[15]), .B2 (n_0_581));
AOI22_X1 i_0_206 (.ZN (n_0_181), .A1 (n_0_183), .A2 (n_0_182), .B1 (n_0_608), .B2 (A[16]));
AOI21_X1 i_0_205 (.ZN (n_0_180), .A (n_0_181), .B1 (B[17]), .B2 (n_0_583));
AOI221_X1 i_0_204 (.ZN (n_0_179), .A (n_0_180), .B1 (n_0_609), .B2 (A[17]), .C1 (n_0_610), .C2 (A[18]));
AOI221_X1 i_0_203 (.ZN (n_0_178), .A (n_0_179), .B1 (B[19]), .B2 (n_0_585), .C1 (B[18]), .C2 (n_0_584));
AOI221_X1 i_0_202 (.ZN (n_0_177), .A (n_0_178), .B1 (n_0_611), .B2 (A[19]), .C1 (n_0_612), .C2 (A[20]));
AOI221_X1 i_0_201 (.ZN (n_0_176), .A (n_0_177), .B1 (B[21]), .B2 (n_0_587), .C1 (B[20]), .C2 (n_0_586));
OAI22_X1 i_0_200 (.ZN (n_0_175), .A1 (B[21]), .A2 (n_0_587), .B1 (B[22]), .B2 (n_0_588));
OAI22_X1 i_0_199 (.ZN (n_0_174), .A1 (n_0_613), .A2 (A[22]), .B1 (n_0_176), .B2 (n_0_175));
AOI21_X1 i_0_198 (.ZN (n_0_173), .A (n_0_396), .B1 (n_102), .B2 (n_0_174));
NAND2_X1 i_0_197 (.ZN (n_0_172), .A1 (A[31]), .A2 (n_0_173));
OAI21_X1 i_0_196 (.ZN (Sum[31]), .A (n_0_172), .B1 (n_0_94), .B2 (n_0_173));
NOR2_X1 i_0_171 (.ZN (n_0_171), .A1 (n_25), .A2 (n_0_228));
AOI22_X1 i_0_170 (.ZN (n_0_170), .A1 (n_0_129), .A2 (\exp_Sum[4] ), .B1 (n_30), .B2 (n_0_266));
AOI22_X1 i_0_169 (.ZN (n_0_169), .A1 (n_29), .A2 (n_0_265), .B1 (n_0_128), .B2 (\exp_Sum[3] ));
AOI22_X1 i_0_168 (.ZN (n_0_168), .A1 (n_28), .A2 (n_0_264), .B1 (n_0_126), .B2 (\exp_Sum[2] ));
INV_X1 i_0_167 (.ZN (n_0_167), .A (n_0_168));
NAND2_X1 i_0_166 (.ZN (n_0_166), .A1 (n_26), .A2 (n_0_262));
INV_X1 i_0_165 (.ZN (n_0_165), .A (n_0_166));
AOI22_X1 i_0_164 (.ZN (n_0_164), .A1 (n_27), .A2 (n_0_263), .B1 (n_0_125), .B2 (\exp_Sum[1] ));
AOI22_X1 i_0_163 (.ZN (n_0_163), .A1 (n_27), .A2 (n_0_263), .B1 (n_0_165), .B2 (n_0_164));
OAI22_X1 i_0_162 (.ZN (n_0_162), .A1 (n_0_126), .A2 (\exp_Sum[2] ), .B1 (n_0_167), .B2 (n_0_163));
AOI22_X1 i_0_161 (.ZN (n_0_161), .A1 (n_29), .A2 (n_0_265), .B1 (n_0_169), .B2 (n_0_162));
AOI22_X1 i_0_160 (.ZN (n_0_160), .A1 (n_0_129), .A2 (\exp_Sum[4] ), .B1 (n_0_170), .B2 (n_0_161));
NAND2_X1 i_0_159 (.ZN (n_0_159), .A1 (n_0_267), .A2 (n_0_160));
NOR2_X1 i_0_158 (.ZN (n_0_158), .A1 (\exp_Sum[6] ), .A2 (n_0_159));
INV_X1 i_0_157 (.ZN (n_0_157), .A (n_0_158));
NAND2_X1 i_0_156 (.ZN (n_0_156), .A1 (n_0_171), .A2 (n_0_158));
AOI21_X1 i_0_155 (.ZN (n_0_155), .A (\exp_Sum[7] ), .B1 (n_0_6), .B2 (n_0_232));
NAND3_X1 i_0_154 (.ZN (n_0_154), .A1 (\num_leading_zeros[4] ), .A2 (\num_leading_zeros[3] ), .A3 (n_0_230));
INV_X1 i_0_153 (.ZN (n_0_153), .A (n_0_154));
AOI221_X1 i_0_152 (.ZN (n_0_152), .A (n_0_153), .B1 (n_0_171), .B2 (n_0_157), .C1 (n_0_563), .C2 (n_0_232));
AOI22_X1 i_0_151 (.ZN (Sum[30]), .A1 (n_0_156), .A2 (n_0_155), .B1 (\exp_Sum[7] ), .B2 (n_0_152));
AOI21_X1 i_0_150 (.ZN (n_0_151), .A (n_0_153), .B1 (n_0_171), .B2 (n_0_159));
NAND2_X1 i_0_149 (.ZN (n_0_150), .A1 (n_0_13), .A2 (n_0_232));
OAI211_X1 i_0_148 (.ZN (Sum[29]), .A (n_0_156), .B (n_0_150), .C1 (n_0_268), .C2 (n_0_151));
OAI21_X1 i_0_147 (.ZN (n_0_149), .A (n_0_159), .B1 (n_0_267), .B2 (n_0_160));
AOI22_X1 i_0_146 (.ZN (n_0_148), .A1 (n_0_12), .A2 (n_0_232), .B1 (n_0_171), .B2 (n_0_149));
OAI21_X1 i_0_145 (.ZN (Sum[28]), .A (n_0_148), .B1 (n_0_267), .B2 (n_0_154));
XOR2_X1 i_0_144 (.Z (n_0_147), .A (n_0_170), .B (n_0_161));
AOI222_X1 i_0_143 (.ZN (n_0_146), .A1 (n_0_11), .A2 (n_0_232), .B1 (\exp_Sum[4] )
    , .B2 (n_0_153), .C1 (n_0_171), .C2 (n_0_147));
INV_X1 i_0_142 (.ZN (Sum[27]), .A (n_0_146));
XNOR2_X1 i_0_141 (.ZN (n_0_145), .A (n_0_169), .B (n_0_162));
AOI222_X1 i_0_140 (.ZN (n_0_144), .A1 (n_0_10), .A2 (n_0_232), .B1 (\exp_Sum[3] )
    , .B2 (n_0_153), .C1 (n_0_171), .C2 (n_0_145));
INV_X1 i_0_139 (.ZN (Sum[26]), .A (n_0_144));
XOR2_X1 i_0_138 (.Z (n_0_143), .A (n_0_168), .B (n_0_163));
AOI222_X1 i_0_137 (.ZN (n_0_142), .A1 (n_0_9), .A2 (n_0_232), .B1 (\exp_Sum[2] ), .B2 (n_0_153)
    , .C1 (n_0_171), .C2 (n_0_143));
INV_X1 i_0_136 (.ZN (Sum[25]), .A (n_0_142));
XOR2_X1 i_0_135 (.Z (n_0_141), .A (n_0_166), .B (n_0_164));
AOI222_X1 i_0_134 (.ZN (n_0_140), .A1 (n_0_8), .A2 (n_0_232), .B1 (\exp_Sum[1] ), .B2 (n_0_153)
    , .C1 (n_0_171), .C2 (n_0_141));
INV_X1 i_0_133 (.ZN (Sum[24]), .A (n_0_140));
OAI21_X1 i_0_132 (.ZN (n_0_139), .A (n_0_166), .B1 (n_26), .B2 (n_0_262));
AOI222_X1 i_0_131 (.ZN (n_0_138), .A1 (n_0_7), .A2 (n_0_232), .B1 (\exp_Sum[0] ), .B2 (n_0_153)
    , .C1 (n_0_171), .C2 (n_0_139));
INV_X1 i_0_130 (.ZN (Sum[23]), .A (n_0_138));
OAI21_X2 i_0_129 (.ZN (n_0_137), .A (n_0_154), .B1 (n_24), .B2 (n_0_233));
AND3_X1 i_0_128 (.ZN (n_0_136), .A1 (n_24), .A2 (n_0_232), .A3 (n_0_225));
AOI22_X1 i_0_127 (.ZN (n_0_135), .A1 (n_22), .A2 (n_0_137), .B1 (n_23), .B2 (n_0_136));
NAND2_X1 i_0_126 (.ZN (n_0_134), .A1 (n_26), .A2 (n_0_229));
INV_X1 i_0_125 (.ZN (n_0_133), .A (n_0_134));
NAND2_X1 i_0_124 (.ZN (n_0_127), .A1 (n_13), .A2 (n_0_119));
AOI22_X1 i_0_123 (.ZN (n_0_124), .A1 (n_21), .A2 (n_0_113), .B1 (n_5), .B2 (n_0_121));
OAI211_X1 i_0_122 (.ZN (n_0_123), .A (n_0_127), .B (n_0_124), .C1 (n_0_126), .C2 (n_0_102));
OAI22_X1 i_0_121 (.ZN (n_0_118), .A1 (n_0_125), .A2 (n_0_110), .B1 (n_27), .B2 (n_0_123));
INV_X1 i_0_120 (.ZN (n_0_117), .A (n_0_118));
NOR2_X2 i_0_119 (.ZN (n_0_116), .A1 (n_26), .A2 (n_0_228));
INV_X1 i_0_118 (.ZN (n_0_115), .A (n_0_116));
AOI22_X1 i_0_117 (.ZN (n_0_108), .A1 (n_14), .A2 (n_0_119), .B1 (n_6), .B2 (n_0_121));
OAI21_X1 i_0_116 (.ZN (n_0_107), .A (n_0_108), .B1 (n_0_126), .B2 (n_0_197));
AOI21_X1 i_0_115 (.ZN (n_0_106), .A (n_0_107), .B1 (n_22), .B2 (n_0_113));
AOI221_X1 i_0_114 (.ZN (n_0_105), .A (n_0_115), .B1 (n_0_125), .B2 (n_0_106), .C1 (n_27), .C2 (n_0_132));
AOI21_X1 i_0_113 (.ZN (n_0_104), .A (n_0_105), .B1 (n_0_133), .B2 (n_0_117));
NAND2_X1 i_0_112 (.ZN (Sum[22]), .A1 (n_0_135), .A2 (n_0_104));
AOI22_X1 i_0_111 (.ZN (n_0_103), .A1 (n_22), .A2 (n_0_136), .B1 (n_0_117), .B2 (n_0_116));
AOI22_X1 i_0_110 (.ZN (n_0_98), .A1 (n_0_133), .A2 (n_0_130), .B1 (n_21), .B2 (n_0_137));
NAND2_X1 i_0_109 (.ZN (Sum[21]), .A1 (n_0_103), .A2 (n_0_98));
NAND2_X1 i_0_108 (.ZN (n_0_97), .A1 (n_21), .A2 (n_0_136));
AOI22_X1 i_0_107 (.ZN (n_0_93), .A1 (n_20), .A2 (n_0_137), .B1 (n_0_116), .B2 (n_0_130));
OAI211_X1 i_0_106 (.ZN (Sum[20]), .A (n_0_97), .B (n_0_93), .C1 (n_0_134), .C2 (n_0_100));
AOI22_X1 i_0_105 (.ZN (n_0_92), .A1 (n_4), .A2 (n_0_120), .B1 (n_12), .B2 (n_0_114));
OAI22_X1 i_0_104 (.ZN (n_0_91), .A1 (n_28), .A2 (n_0_194), .B1 (n_0_126), .B2 (n_0_92));
AOI22_X1 i_0_103 (.ZN (n_0_90), .A1 (n_0_125), .A2 (n_0_195), .B1 (n_27), .B2 (n_0_91));
AOI22_X1 i_0_102 (.ZN (n_0_89), .A1 (n_20), .A2 (n_0_136), .B1 (n_19), .B2 (n_0_137));
OAI221_X1 i_0_101 (.ZN (Sum[19]), .A (n_0_89), .B1 (n_0_134), .B2 (n_0_90), .C1 (n_0_115), .C2 (n_0_100));
AOI22_X1 i_0_100 (.ZN (n_0_88), .A1 (n_19), .A2 (n_0_136), .B1 (n_18), .B2 (n_0_137));
NOR3_X2 i_0_99 (.ZN (n_0_87), .A1 (n_30), .A2 (n_29), .A3 (n_0_126));
NOR3_X1 i_0_98 (.ZN (n_0_86), .A1 (n_30), .A2 (n_0_128), .A3 (n_0_126));
AOI22_X1 i_0_97 (.ZN (n_0_85), .A1 (n_11), .A2 (n_0_87), .B1 (n_3), .B2 (n_0_86));
OAI21_X1 i_0_96 (.ZN (n_0_84), .A (n_0_85), .B1 (n_28), .B2 (n_0_112));
AOI22_X1 i_0_95 (.ZN (n_0_83), .A1 (n_27), .A2 (n_0_84), .B1 (n_0_125), .B2 (n_0_101));
OAI221_X1 i_0_94 (.ZN (Sum[18]), .A (n_0_88), .B1 (n_0_115), .B2 (n_0_90), .C1 (n_0_134), .C2 (n_0_83));
AOI22_X1 i_0_93 (.ZN (n_0_82), .A1 (n_17), .A2 (n_0_137), .B1 (n_18), .B2 (n_0_136));
AOI22_X1 i_0_92 (.ZN (n_0_81), .A1 (n_10), .A2 (n_0_87), .B1 (n_2), .B2 (n_0_86));
OAI21_X1 i_0_91 (.ZN (n_0_80), .A (n_0_81), .B1 (n_28), .B2 (n_0_196));
AOI22_X1 i_0_90 (.ZN (n_0_79), .A1 (n_0_125), .A2 (n_0_91), .B1 (n_27), .B2 (n_0_80));
OAI221_X1 i_0_89 (.ZN (Sum[17]), .A (n_0_82), .B1 (n_0_134), .B2 (n_0_79), .C1 (n_0_115), .C2 (n_0_83));
AOI22_X1 i_0_88 (.ZN (n_0_78), .A1 (n_1), .A2 (n_0_86), .B1 (n_9), .B2 (n_0_87));
OAI21_X1 i_0_87 (.ZN (n_0_77), .A (n_0_78), .B1 (n_28), .B2 (n_0_109));
AOI22_X1 i_0_86 (.ZN (n_0_76), .A1 (n_0_125), .A2 (n_0_84), .B1 (n_27), .B2 (n_0_77));
INV_X1 i_0_85 (.ZN (n_0_75), .A (n_0_76));
AOI22_X1 i_0_84 (.ZN (n_0_74), .A1 (n_0_133), .A2 (n_0_75), .B1 (n_17), .B2 (n_0_136));
NAND2_X1 i_0_83 (.ZN (n_0_73), .A1 (n_16), .A2 (n_0_137));
OAI211_X1 i_0_82 (.ZN (Sum[16]), .A (n_0_74), .B (n_0_73), .C1 (n_0_115), .C2 (n_0_79));
AOI22_X1 i_0_81 (.ZN (n_0_72), .A1 (n_0), .A2 (n_0_86), .B1 (n_8), .B2 (n_0_87));
OAI21_X1 i_0_80 (.ZN (n_0_71), .A (n_0_72), .B1 (n_28), .B2 (n_0_92));
AOI22_X1 i_0_79 (.ZN (n_0_70), .A1 (n_0_125), .A2 (n_0_80), .B1 (n_27), .B2 (n_0_71));
AOI22_X1 i_0_78 (.ZN (n_0_69), .A1 (n_16), .A2 (n_0_136), .B1 (n_15), .B2 (n_0_137));
OAI221_X1 i_0_77 (.ZN (Sum[15]), .A (n_0_69), .B1 (n_0_134), .B2 (n_0_70), .C1 (n_0_115), .C2 (n_0_76));
AOI222_X1 i_0_76 (.ZN (n_0_68), .A1 (n_11), .A2 (n_0_113), .B1 (n_3), .B2 (n_0_119)
    , .C1 (n_7), .C2 (n_0_87));
NAND2_X1 i_0_75 (.ZN (n_0_67), .A1 (n_0_125), .A2 (n_0_77));
OAI21_X1 i_0_74 (.ZN (n_0_66), .A (n_0_67), .B1 (n_0_125), .B2 (n_0_68));
AOI22_X1 i_0_73 (.ZN (n_0_65), .A1 (n_15), .A2 (n_0_136), .B1 (n_0_133), .B2 (n_0_66));
NAND2_X1 i_0_72 (.ZN (n_0_64), .A1 (n_14), .A2 (n_0_137));
OAI211_X1 i_0_71 (.ZN (Sum[14]), .A (n_0_64), .B (n_0_65), .C1 (n_0_115), .C2 (n_0_70));
AOI22_X1 i_0_70 (.ZN (n_0_63), .A1 (n_0_116), .A2 (n_0_66), .B1 (n_14), .B2 (n_0_136));
AOI222_X1 i_0_69 (.ZN (n_0_62), .A1 (n_10), .A2 (n_0_113), .B1 (n_2), .B2 (n_0_119)
    , .C1 (n_6), .C2 (n_0_87));
NAND2_X1 i_0_68 (.ZN (n_0_61), .A1 (n_0_125), .A2 (n_0_71));
OAI21_X1 i_0_67 (.ZN (n_0_60), .A (n_0_61), .B1 (n_0_125), .B2 (n_0_62));
AOI22_X1 i_0_66 (.ZN (n_0_59), .A1 (n_13), .A2 (n_0_137), .B1 (n_0_133), .B2 (n_0_60));
NAND2_X1 i_0_65 (.ZN (Sum[13]), .A1 (n_0_63), .A2 (n_0_59));
AOI222_X1 i_0_64 (.ZN (n_0_58), .A1 (n_9), .A2 (n_0_113), .B1 (n_1), .B2 (n_0_119)
    , .C1 (n_5), .C2 (n_0_87));
OAI22_X1 i_0_63 (.ZN (n_0_57), .A1 (n_27), .A2 (n_0_68), .B1 (n_0_125), .B2 (n_0_58));
AOI22_X1 i_0_62 (.ZN (n_0_56), .A1 (n_0_133), .A2 (n_0_57), .B1 (n_13), .B2 (n_0_136));
AOI22_X1 i_0_61 (.ZN (n_0_55), .A1 (n_12), .A2 (n_0_137), .B1 (n_0_116), .B2 (n_0_60));
NAND2_X1 i_0_60 (.ZN (Sum[12]), .A1 (n_0_56), .A2 (n_0_55));
AOI22_X1 i_0_59 (.ZN (n_0_54), .A1 (n_11), .A2 (n_0_137), .B1 (n_12), .B2 (n_0_136));
AOI222_X1 i_0_58 (.ZN (n_0_53), .A1 (n_8), .A2 (n_0_113), .B1 (n_0), .B2 (n_0_119)
    , .C1 (n_4), .C2 (n_0_87));
OAI22_X1 i_0_57 (.ZN (n_0_52), .A1 (n_27), .A2 (n_0_62), .B1 (n_0_125), .B2 (n_0_53));
AOI22_X1 i_0_56 (.ZN (n_0_51), .A1 (n_0_133), .A2 (n_0_52), .B1 (n_0_116), .B2 (n_0_57));
NAND2_X1 i_0_55 (.ZN (Sum[11]), .A1 (n_0_54), .A2 (n_0_51));
AOI22_X1 i_0_54 (.ZN (n_0_50), .A1 (n_0_116), .A2 (n_0_52), .B1 (n_11), .B2 (n_0_136));
AOI22_X1 i_0_53 (.ZN (n_0_49), .A1 (n_7), .A2 (n_0_113), .B1 (n_3), .B2 (n_0_87));
OAI22_X1 i_0_52 (.ZN (n_0_48), .A1 (n_0_125), .A2 (n_0_49), .B1 (n_27), .B2 (n_0_58));
AOI22_X1 i_0_51 (.ZN (n_0_47), .A1 (n_10), .A2 (n_0_137), .B1 (n_0_133), .B2 (n_0_48));
NAND2_X1 i_0_50 (.ZN (Sum[10]), .A1 (n_0_50), .A2 (n_0_47));
AOI22_X1 i_0_49 (.ZN (n_0_46), .A1 (n_6), .A2 (n_0_113), .B1 (n_2), .B2 (n_0_87));
OAI22_X1 i_0_48 (.ZN (n_0_45), .A1 (n_27), .A2 (n_0_53), .B1 (n_0_125), .B2 (n_0_46));
AOI22_X1 i_0_47 (.ZN (n_0_44), .A1 (n_0_133), .A2 (n_0_45), .B1 (n_10), .B2 (n_0_136));
AOI22_X1 i_0_46 (.ZN (n_0_43), .A1 (n_9), .A2 (n_0_137), .B1 (n_0_116), .B2 (n_0_48));
NAND2_X1 i_0_45 (.ZN (Sum[9]), .A1 (n_0_44), .A2 (n_0_43));
AOI22_X1 i_0_44 (.ZN (n_0_42), .A1 (n_9), .A2 (n_0_136), .B1 (n_8), .B2 (n_0_137));
AOI22_X1 i_0_43 (.ZN (n_0_41), .A1 (n_5), .A2 (n_0_113), .B1 (n_1), .B2 (n_0_87));
OAI22_X1 i_0_42 (.ZN (n_0_40), .A1 (n_27), .A2 (n_0_49), .B1 (n_0_125), .B2 (n_0_41));
AOI22_X1 i_0_41 (.ZN (n_0_39), .A1 (n_0_116), .A2 (n_0_45), .B1 (n_0_133), .B2 (n_0_40));
NAND2_X1 i_0_40 (.ZN (Sum[8]), .A1 (n_0_42), .A2 (n_0_39));
AOI22_X1 i_0_39 (.ZN (n_0_38), .A1 (n_8), .A2 (n_0_136), .B1 (n_0_116), .B2 (n_0_40));
AOI22_X1 i_0_38 (.ZN (n_0_37), .A1 (n_4), .A2 (n_0_113), .B1 (n_0), .B2 (n_0_87));
OAI22_X1 i_0_37 (.ZN (n_0_36), .A1 (n_27), .A2 (n_0_46), .B1 (n_0_125), .B2 (n_0_37));
AOI22_X1 i_0_36 (.ZN (n_0_35), .A1 (n_0_133), .A2 (n_0_36), .B1 (n_7), .B2 (n_0_137));
NAND2_X1 i_0_35 (.ZN (Sum[7]), .A1 (n_0_38), .A2 (n_0_35));
AND2_X1 i_0_34 (.ZN (n_0_34), .A1 (n_27), .A2 (n_0_113));
NAND2_X1 i_0_33 (.ZN (n_0_33), .A1 (n_3), .A2 (n_0_34));
OAI21_X1 i_0_32 (.ZN (n_0_32), .A (n_0_33), .B1 (n_27), .B2 (n_0_41));
AOI22_X1 i_0_31 (.ZN (n_0_31), .A1 (n_0_133), .A2 (n_0_32), .B1 (n_7), .B2 (n_0_136));
AOI22_X1 i_0_30 (.ZN (n_0_30), .A1 (n_6), .A2 (n_0_137), .B1 (n_0_116), .B2 (n_0_36));
NAND2_X1 i_0_29 (.ZN (Sum[6]), .A1 (n_0_31), .A2 (n_0_30));
AOI22_X1 i_0_28 (.ZN (n_0_29), .A1 (n_6), .A2 (n_0_136), .B1 (n_0_116), .B2 (n_0_32));
NAND2_X1 i_0_27 (.ZN (n_0_28), .A1 (n_2), .A2 (n_0_34));
OAI21_X1 i_0_26 (.ZN (n_0_27), .A (n_0_28), .B1 (n_27), .B2 (n_0_37));
AOI22_X1 i_0_25 (.ZN (n_0_26), .A1 (n_0_133), .A2 (n_0_27), .B1 (n_5), .B2 (n_0_137));
NAND2_X1 i_0_24 (.ZN (Sum[5]), .A1 (n_0_29), .A2 (n_0_26));
AND2_X1 i_0_23 (.ZN (n_0_25), .A1 (n_0_125), .A2 (n_0_113));
AOI22_X1 i_0_22 (.ZN (n_0_24), .A1 (n_1), .A2 (n_0_34), .B1 (n_3), .B2 (n_0_25));
AOI222_X1 i_0_21 (.ZN (n_0_23), .A1 (n_5), .A2 (n_0_136), .B1 (n_4), .B2 (n_0_137)
    , .C1 (n_0_116), .C2 (n_0_27));
OAI21_X1 i_0_20 (.ZN (Sum[4]), .A (n_0_23), .B1 (n_0_134), .B2 (n_0_24));
AOI22_X1 i_0_19 (.ZN (n_0_22), .A1 (n_3), .A2 (n_0_137), .B1 (n_4), .B2 (n_0_136));
AOI22_X1 i_0_18 (.ZN (n_0_21), .A1 (n_0), .A2 (n_0_34), .B1 (n_2), .B2 (n_0_25));
OAI221_X1 i_0_17 (.ZN (Sum[3]), .A (n_0_22), .B1 (n_0_134), .B2 (n_0_21), .C1 (n_0_115), .C2 (n_0_24));
NAND2_X1 i_0_16 (.ZN (n_0_20), .A1 (n_1), .A2 (n_0_25));
AOI22_X1 i_0_15 (.ZN (n_0_19), .A1 (n_3), .A2 (n_0_136), .B1 (n_2), .B2 (n_0_137));
OAI221_X1 i_0_14 (.ZN (Sum[2]), .A (n_0_19), .B1 (n_0_134), .B2 (n_0_20), .C1 (n_0_115), .C2 (n_0_21));
AOI21_X1 i_0_13 (.ZN (n_0_18), .A (n_0_137), .B1 (n_0_116), .B2 (n_0_25));
INV_X1 i_0_12 (.ZN (n_0_17), .A (n_0_18));
NAND2_X1 i_0_11 (.ZN (n_0_16), .A1 (n_0), .A2 (n_0_25));
AOI22_X1 i_0_10 (.ZN (n_0_15), .A1 (n_1), .A2 (n_0_17), .B1 (n_2), .B2 (n_0_136));
OAI21_X1 i_0_9 (.ZN (Sum[1]), .A (n_0_15), .B1 (n_0_134), .B2 (n_0_16));
AOI22_X1 i_0_8 (.ZN (n_0_14), .A1 (n_0), .A2 (n_0_17), .B1 (n_1), .B2 (n_0_136));
INV_X1 i_0_7 (.ZN (Sum[0]), .A (n_0_14));
HA_X1 i_0_6 (.CO (n_0_6), .S (n_0_13), .A (\exp_Sum[6] ), .B (n_0_5));
HA_X1 i_0_5 (.CO (n_0_5), .S (n_0_12), .A (\exp_Sum[5] ), .B (n_0_4));
HA_X1 i_0_4 (.CO (n_0_4), .S (n_0_11), .A (\exp_Sum[4] ), .B (n_0_3));
HA_X1 i_0_3 (.CO (n_0_3), .S (n_0_10), .A (\exp_Sum[3] ), .B (n_0_2));
HA_X1 i_0_2 (.CO (n_0_2), .S (n_0_9), .A (\exp_Sum[2] ), .B (n_0_1));
HA_X1 i_0_1 (.CO (n_0_1), .S (n_0_8), .A (\exp_Sum[1] ), .B (n_0_0));
HA_X1 i_0_0 (.CO (n_0_0), .S (n_0_7), .A (n_24), .B (\exp_Sum[0] ));
datapath__0_43 i_22 (.p_0 ({n_54, uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, 
    n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
    n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, uc_35}), .mant_A ({
    n_100, n_76, n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, 
    n_64, n_63, n_62, n_99, n_61, n_60, n_59, n_58, n_57, n_56, n_55}));
datapath__0_38 i_17 (.p_1 ({uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, n_30, n_29, 
    n_28, n_27, n_26}), .p_0 ({1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 
    1'b0 , 1'b0 , \num_leading_zeros[0] , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 
    \num_leading_zeros[4] , \num_leading_zeros[3] , \num_leading_zeros[2] , \num_leading_zeros[1] , 
    1'b1 }));
datapath__0_25 i_5 (.p_0 (n_25), .exp_Sum ({\exp_Sum[7] , \exp_Sum[6] , \exp_Sum[5] , 
    \exp_Sum[4] , \exp_Sum[3] , \exp_Sum[2] , \exp_Sum[1] , \exp_Sum[0] }), .p_1 ({
    1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , \num_leading_zeros[0] , 
    1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , \num_leading_zeros[4] , \num_leading_zeros[3] , 
    \num_leading_zeros[2] , \num_leading_zeros[1] , 1'b1 }));
count_leading_zeros count_leading_zeros_instance (.result ({\num_leading_zeros[4] , 
    \num_leading_zeros[3] , \num_leading_zeros[2] , \num_leading_zeros[1] , \num_leading_zeros[0] })
    , .valueIn ({n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
    n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}));
CLA CLA_dut (.sum ({uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, n_24, n_23, 
    n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, 
    n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}), .in1 ({\mant_A[31] , uc_0, 
    uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, \mant_A[23] , \mant_A[22] , \mant_A[21] , 
    \mant_A[20] , \mant_A[19] , \mant_A[18] , \mant_A[17] , \mant_A[16] , \mant_A[15] , 
    \mant_A[14] , \mant_A[13] , \mant_A[12] , \mant_A[11] , \mant_A[10] , \mant_A[9] , 
    \mant_A[8] , \mant_A[7] , \mant_A[6] , \mant_A[5] , \mant_A[4] , \mant_A[3] , 
    \mant_A[2] , \mant_A[1] , n_55}), .in2 ({uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, 
    uc_13, uc_14, n_102, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, n_89, 
    n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_101, n_81, n_80, n_79, n_78, n_77}));
CLKBUF_X1 drc_ipo_c4 (.Z (drc_ipo_n4), .A (n_0_470));

endmodule //fp_adder

module buffer__0_58 (clk_CTS_1_PP_0, clk, rst, en, D, Q);

output [31:0] Q;
input [31:0] D;
input clk;
input en;
input rst;
input clk_CTS_1_PP_0;
wire n_0_0;
wire n_1;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid1_48;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (D[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (D[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (D[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (D[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (D[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (D[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (D[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (D[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (D[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (D[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (D[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (D[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (D[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (D[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (D[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (D[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (D[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (D[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (D[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (D[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (D[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (D[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (D[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (D[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (D[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (D[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (D[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (D[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (D[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (D[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (D[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (D[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (rst));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (rst));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (CTS_n_tid1_48), .D (n_2));
DFF_X1 \Q_reg[1]  (.Q (Q[1]), .CK (CTS_n_tid1_48), .D (n_3));
DFF_X1 \Q_reg[2]  (.Q (Q[2]), .CK (CTS_n_tid1_48), .D (n_4));
DFF_X1 \Q_reg[3]  (.Q (Q[3]), .CK (CTS_n_tid1_48), .D (n_5));
DFF_X1 \Q_reg[4]  (.Q (Q[4]), .CK (CTS_n_tid1_48), .D (n_6));
DFF_X1 \Q_reg[5]  (.Q (Q[5]), .CK (CTS_n_tid1_48), .D (n_7));
DFF_X1 \Q_reg[6]  (.Q (Q[6]), .CK (CTS_n_tid1_48), .D (n_8));
DFF_X1 \Q_reg[7]  (.Q (Q[7]), .CK (CTS_n_tid1_48), .D (n_9));
DFF_X1 \Q_reg[8]  (.Q (Q[8]), .CK (CTS_n_tid1_48), .D (n_10));
DFF_X1 \Q_reg[9]  (.Q (Q[9]), .CK (CTS_n_tid1_48), .D (n_11));
DFF_X1 \Q_reg[10]  (.Q (Q[10]), .CK (CTS_n_tid1_48), .D (n_12));
DFF_X1 \Q_reg[11]  (.Q (Q[11]), .CK (CTS_n_tid1_48), .D (n_13));
DFF_X1 \Q_reg[12]  (.Q (Q[12]), .CK (CTS_n_tid1_48), .D (n_14));
DFF_X1 \Q_reg[13]  (.Q (Q[13]), .CK (CTS_n_tid1_48), .D (n_15));
DFF_X1 \Q_reg[14]  (.Q (Q[14]), .CK (CTS_n_tid1_48), .D (n_16));
DFF_X1 \Q_reg[15]  (.Q (Q[15]), .CK (CTS_n_tid1_48), .D (n_17));
DFF_X1 \Q_reg[16]  (.Q (Q[16]), .CK (CTS_n_tid1_48), .D (n_18));
DFF_X1 \Q_reg[17]  (.Q (Q[17]), .CK (CTS_n_tid1_48), .D (n_19));
DFF_X1 \Q_reg[18]  (.Q (Q[18]), .CK (CTS_n_tid1_48), .D (n_20));
DFF_X1 \Q_reg[19]  (.Q (Q[19]), .CK (CTS_n_tid1_48), .D (n_21));
DFF_X1 \Q_reg[20]  (.Q (Q[20]), .CK (CTS_n_tid1_48), .D (n_22));
DFF_X1 \Q_reg[21]  (.Q (Q[21]), .CK (CTS_n_tid1_48), .D (n_23));
DFF_X1 \Q_reg[22]  (.Q (Q[22]), .CK (CTS_n_tid1_48), .D (n_24));
DFF_X1 \Q_reg[23]  (.Q (Q[23]), .CK (CTS_n_tid1_48), .D (n_25));
DFF_X1 \Q_reg[24]  (.Q (Q[24]), .CK (CTS_n_tid1_48), .D (n_26));
DFF_X1 \Q_reg[25]  (.Q (Q[25]), .CK (CTS_n_tid1_48), .D (n_27));
DFF_X1 \Q_reg[26]  (.Q (Q[26]), .CK (CTS_n_tid1_48), .D (n_28));
DFF_X1 \Q_reg[27]  (.Q (Q[27]), .CK (CTS_n_tid1_48), .D (n_29));
DFF_X1 \Q_reg[28]  (.Q (Q[28]), .CK (CTS_n_tid1_48), .D (n_30));
DFF_X1 \Q_reg[29]  (.Q (Q[29]), .CK (CTS_n_tid1_48), .D (n_31));
DFF_X1 \Q_reg[30]  (.Q (Q[30]), .CK (CTS_n_tid1_48), .D (n_32));
DFF_X1 \Q_reg[31]  (.Q (Q[31]), .CK (CTS_n_tid1_48), .D (n_33));
CLKGATETST_X8 clk_gate_Q_reg (.GCK (CTS_n_tid1_48), .CK (clk_CTS_1_PP_0), .E (n_1), .SE (1'b0 ));

endmodule //buffer__0_58

module buffer__0_55 (clk_CTS_1_PP_0, clk, rst, en, D, Q);

output [31:0] Q;
input [31:0] D;
input clk;
input en;
input rst;
input clk_CTS_1_PP_0;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (D[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (D[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (D[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (D[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (D[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (D[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (D[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (D[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (D[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (D[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (D[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (D[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (D[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (D[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (D[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (D[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (D[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (D[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (D[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (D[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (D[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (D[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (D[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (D[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (D[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (D[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (D[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (D[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (D[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (D[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (D[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (D[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (rst));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (rst));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (n_0), .D (n_2));
DFF_X1 \Q_reg[1]  (.Q (Q[1]), .CK (n_0), .D (n_3));
DFF_X1 \Q_reg[2]  (.Q (Q[2]), .CK (n_0), .D (n_4));
DFF_X1 \Q_reg[3]  (.Q (Q[3]), .CK (n_0), .D (n_5));
DFF_X1 \Q_reg[4]  (.Q (Q[4]), .CK (n_0), .D (n_6));
DFF_X1 \Q_reg[5]  (.Q (Q[5]), .CK (n_0), .D (n_7));
DFF_X1 \Q_reg[6]  (.Q (Q[6]), .CK (n_0), .D (n_8));
DFF_X1 \Q_reg[7]  (.Q (Q[7]), .CK (n_0), .D (n_9));
DFF_X1 \Q_reg[8]  (.Q (Q[8]), .CK (n_0), .D (n_10));
DFF_X1 \Q_reg[9]  (.Q (Q[9]), .CK (n_0), .D (n_11));
DFF_X1 \Q_reg[10]  (.Q (Q[10]), .CK (n_0), .D (n_12));
DFF_X1 \Q_reg[11]  (.Q (Q[11]), .CK (n_0), .D (n_13));
DFF_X1 \Q_reg[12]  (.Q (Q[12]), .CK (n_0), .D (n_14));
DFF_X1 \Q_reg[13]  (.Q (Q[13]), .CK (n_0), .D (n_15));
DFF_X1 \Q_reg[14]  (.Q (Q[14]), .CK (n_0), .D (n_16));
DFF_X1 \Q_reg[15]  (.Q (Q[15]), .CK (n_0), .D (n_17));
DFF_X1 \Q_reg[16]  (.Q (Q[16]), .CK (n_0), .D (n_18));
DFF_X1 \Q_reg[17]  (.Q (Q[17]), .CK (n_0), .D (n_19));
DFF_X1 \Q_reg[18]  (.Q (Q[18]), .CK (n_0), .D (n_20));
DFF_X1 \Q_reg[19]  (.Q (Q[19]), .CK (n_0), .D (n_21));
DFF_X1 \Q_reg[20]  (.Q (Q[20]), .CK (n_0), .D (n_22));
DFF_X1 \Q_reg[21]  (.Q (Q[21]), .CK (n_0), .D (n_23));
DFF_X1 \Q_reg[22]  (.Q (Q[22]), .CK (n_0), .D (n_24));
DFF_X1 \Q_reg[23]  (.Q (Q[23]), .CK (n_0), .D (n_25));
DFF_X1 \Q_reg[24]  (.Q (Q[24]), .CK (n_0), .D (n_26));
DFF_X1 \Q_reg[25]  (.Q (Q[25]), .CK (n_0), .D (n_27));
DFF_X1 \Q_reg[26]  (.Q (Q[26]), .CK (n_0), .D (n_28));
DFF_X1 \Q_reg[27]  (.Q (Q[27]), .CK (n_0), .D (n_29));
DFF_X1 \Q_reg[28]  (.Q (Q[28]), .CK (n_0), .D (n_30));
DFF_X1 \Q_reg[29]  (.Q (Q[29]), .CK (n_0), .D (n_31));
DFF_X1 \Q_reg[30]  (.Q (Q[30]), .CK (n_0), .D (n_32));
DFF_X1 \Q_reg[31]  (.Q (Q[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_Q_reg (.GCK (n_0), .CK (clk_CTS_1_PP_0), .E (n_1), .SE (1'b0 ));

endmodule //buffer__0_55

module fp_adder_buff (clk, rst, en, a, b, sum, overflow, underflow);

output overflow;
output [31:0] sum;
output underflow;
input [31:0] a;
input [31:0] b;
input clk;
input en;
input rst;
wire CTS_n_tid1_3;
wire \a_out[31] ;
wire \a_out[30] ;
wire \a_out[29] ;
wire \a_out[28] ;
wire \a_out[27] ;
wire \a_out[26] ;
wire \a_out[25] ;
wire \a_out[24] ;
wire \a_out[23] ;
wire \a_out[22] ;
wire \a_out[21] ;
wire \a_out[20] ;
wire \a_out[19] ;
wire \a_out[18] ;
wire \a_out[17] ;
wire \a_out[16] ;
wire \a_out[15] ;
wire \a_out[14] ;
wire \a_out[13] ;
wire \a_out[12] ;
wire \a_out[11] ;
wire \a_out[10] ;
wire \a_out[9] ;
wire \a_out[8] ;
wire \a_out[7] ;
wire \a_out[6] ;
wire \a_out[5] ;
wire \a_out[4] ;
wire \a_out[3] ;
wire \a_out[2] ;
wire \a_out[1] ;
wire \a_out[0] ;
wire \b_out[31] ;
wire \b_out[30] ;
wire \b_out[29] ;
wire \b_out[28] ;
wire \b_out[27] ;
wire \b_out[26] ;
wire \b_out[25] ;
wire \b_out[24] ;
wire \b_out[23] ;
wire \b_out[22] ;
wire \b_out[21] ;
wire \b_out[20] ;
wire \b_out[19] ;
wire \b_out[18] ;
wire \b_out[17] ;
wire \b_out[16] ;
wire \b_out[15] ;
wire \b_out[14] ;
wire \b_out[13] ;
wire \b_out[12] ;
wire \b_out[11] ;
wire \b_out[10] ;
wire \b_out[9] ;
wire \b_out[8] ;
wire \b_out[7] ;
wire \b_out[6] ;
wire \b_out[5] ;
wire \b_out[4] ;
wire \b_out[3] ;
wire \b_out[2] ;
wire \b_out[1] ;
wire \b_out[0] ;
wire underflow_out;
wire overflow_out;
wire \sum_out[31] ;
wire \sum_out[30] ;
wire \sum_out[29] ;
wire \sum_out[28] ;
wire \sum_out[27] ;
wire \sum_out[26] ;
wire \sum_out[25] ;
wire \sum_out[24] ;
wire \sum_out[23] ;
wire \sum_out[22] ;
wire \sum_out[21] ;
wire \sum_out[20] ;
wire \sum_out[19] ;
wire \sum_out[18] ;
wire \sum_out[17] ;
wire \sum_out[16] ;
wire \sum_out[15] ;
wire \sum_out[14] ;
wire \sum_out[13] ;
wire \sum_out[12] ;
wire \sum_out[11] ;
wire \sum_out[10] ;
wire \sum_out[9] ;
wire \sum_out[8] ;
wire \sum_out[7] ;
wire \sum_out[6] ;
wire \sum_out[5] ;
wire \sum_out[4] ;
wire \sum_out[3] ;
wire \sum_out[2] ;
wire \sum_out[1] ;
wire \sum_out[0] ;


buffer__parameterized0 outRegU (.Q ({underflow}), .D ({underflow_out}), .en (en), .rst (rst)
    , .clk_CTS_1_PP_0 (CTS_n_tid1_3));
buffer__parameterized0__0_52 outRegO (.Q ({overflow}), .clk_CTS_1_PP_0 (CTS_n_tid1_3)
    , .D ({overflow_out}), .en (en), .rst (rst), .clk_CTS_1_PP_8 (clk));
buffer outRegS (.Q ({sum[31], sum[30], sum[29], sum[28], sum[27], sum[26], sum[25], 
    sum[24], sum[23], sum[22], sum[21], sum[20], sum[19], sum[18], sum[17], sum[16], 
    sum[15], sum[14], sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], sum[7], 
    sum[6], sum[5], sum[4], sum[3], sum[2], sum[1], sum[0]}), .D ({\sum_out[31] , 
    \sum_out[30] , \sum_out[29] , \sum_out[28] , \sum_out[27] , \sum_out[26] , \sum_out[25] , 
    \sum_out[24] , \sum_out[23] , \sum_out[22] , \sum_out[21] , \sum_out[20] , \sum_out[19] , 
    \sum_out[18] , \sum_out[17] , \sum_out[16] , \sum_out[15] , \sum_out[14] , \sum_out[13] , 
    \sum_out[12] , \sum_out[11] , \sum_out[10] , \sum_out[9] , \sum_out[8] , \sum_out[7] , 
    \sum_out[6] , \sum_out[5] , \sum_out[4] , \sum_out[3] , \sum_out[2] , \sum_out[1] , 
    \sum_out[0] }), .en (en), .rst (rst), .clk_CTS_1_PP_3 (clk));
fp_adder A32 (.Sum ({\sum_out[31] , \sum_out[30] , \sum_out[29] , \sum_out[28] , 
    \sum_out[27] , \sum_out[26] , \sum_out[25] , \sum_out[24] , \sum_out[23] , \sum_out[22] , 
    \sum_out[21] , \sum_out[20] , \sum_out[19] , \sum_out[18] , \sum_out[17] , \sum_out[16] , 
    \sum_out[15] , \sum_out[14] , \sum_out[13] , \sum_out[12] , \sum_out[11] , \sum_out[10] , 
    \sum_out[9] , \sum_out[8] , \sum_out[7] , \sum_out[6] , \sum_out[5] , \sum_out[4] , 
    \sum_out[3] , \sum_out[2] , \sum_out[1] , \sum_out[0] }), .overflow (overflow_out)
    , .underflow (underflow_out), .A ({\a_out[31] , \a_out[30] , \a_out[29] , \a_out[28] , 
    \a_out[27] , \a_out[26] , \a_out[25] , \a_out[24] , \a_out[23] , \a_out[22] , 
    \a_out[21] , \a_out[20] , \a_out[19] , \a_out[18] , \a_out[17] , \a_out[16] , 
    \a_out[15] , \a_out[14] , \a_out[13] , \a_out[12] , \a_out[11] , \a_out[10] , 
    \a_out[9] , \a_out[8] , \a_out[7] , \a_out[6] , \a_out[5] , \a_out[4] , \a_out[3] , 
    \a_out[2] , \a_out[1] , \a_out[0] }), .B ({\b_out[31] , \b_out[30] , \b_out[29] , 
    \b_out[28] , \b_out[27] , \b_out[26] , \b_out[25] , \b_out[24] , \b_out[23] , 
    \b_out[22] , \b_out[21] , \b_out[20] , \b_out[19] , \b_out[18] , \b_out[17] , 
    \b_out[16] , \b_out[15] , \b_out[14] , \b_out[13] , \b_out[12] , \b_out[11] , 
    \b_out[10] , \b_out[9] , \b_out[8] , \b_out[7] , \b_out[6] , \b_out[5] , \b_out[4] , 
    \b_out[3] , \b_out[2] , \b_out[1] , \b_out[0] }));
buffer__0_58 inRegB (.Q ({\b_out[31] , \b_out[30] , \b_out[29] , \b_out[28] , \b_out[27] , 
    \b_out[26] , \b_out[25] , \b_out[24] , \b_out[23] , \b_out[22] , \b_out[21] , 
    \b_out[20] , \b_out[19] , \b_out[18] , \b_out[17] , \b_out[16] , \b_out[15] , 
    \b_out[14] , \b_out[13] , \b_out[12] , \b_out[11] , \b_out[10] , \b_out[9] , 
    \b_out[8] , \b_out[7] , \b_out[6] , \b_out[5] , \b_out[4] , \b_out[3] , \b_out[2] , 
    \b_out[1] , \b_out[0] }), .D ({b[31], b[30], b[29], b[28], b[27], b[26], b[25], 
    b[24], b[23], b[22], b[21], b[20], b[19], b[18], b[17], b[16], b[15], b[14], 
    b[13], b[12], b[11], b[10], b[9], b[8], b[7], b[6], b[5], b[4], b[3], b[2], b[1], 
    b[0]}), .en (en), .rst (rst), .clk_CTS_1_PP_0 (CTS_n_tid1_3));
buffer__0_55 inRegA (.Q ({\a_out[31] , \a_out[30] , \a_out[29] , \a_out[28] , \a_out[27] , 
    \a_out[26] , \a_out[25] , \a_out[24] , \a_out[23] , \a_out[22] , \a_out[21] , 
    \a_out[20] , \a_out[19] , \a_out[18] , \a_out[17] , \a_out[16] , \a_out[15] , 
    \a_out[14] , \a_out[13] , \a_out[12] , \a_out[11] , \a_out[10] , \a_out[9] , 
    \a_out[8] , \a_out[7] , \a_out[6] , \a_out[5] , \a_out[4] , \a_out[3] , \a_out[2] , 
    \a_out[1] , \a_out[0] }), .D ({a[31], a[30], a[29], a[28], a[27], a[26], a[25], 
    a[24], a[23], a[22], a[21], a[20], a[19], a[18], a[17], a[16], a[15], a[14], 
    a[13], a[12], a[11], a[10], a[9], a[8], a[7], a[6], a[5], a[4], a[3], a[2], a[1], 
    a[0]}), .en (en), .rst (rst), .clk_CTS_1_PP_0 (CTS_n_tid1_3));

endmodule //fp_adder_buff


