/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 16 17:42:20 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2338596271 */

module datapath(p_0, b);
   output [31:0]p_0;
   input [31:0]b;

   XOR2_X1 i_0 (.A(b[1]), .B(b[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(b[2]), .B1(b[1]), .B2(b[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(b[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(b[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(b[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(b[6]), .B1(n_27), .B2(b[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(b[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(b[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(b[9]), .B1(n_25), .B2(b[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(b[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(b[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(b[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(b[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(b[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(b[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(b[16]), .B1(n_19), .B2(b[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(b[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(b[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(b[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(b[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(b[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(b[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(b[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(b[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(b[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(b[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(b[27]), .B1(n_9), .B2(b[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(b[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(b[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(b[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(b[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(b[28]), .A3(b[29]), .A4(b[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(b[28]), .A3(b[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(b[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(b[26]), .A3(b[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(b[23]), .A3(b[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(b[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(b[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(b[18]), .A3(b[19]), .A4(b[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(b[18]), .A3(b[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(b[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(b[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(b[15]), .A3(b[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(b[12]), .A3(b[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(b[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(b[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(b[8]), .A3(b[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(b[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(b[5]), .A3(b[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(b[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(b[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(b[2]), .A2(b[1]), .A3(b[0]), .ZN(n_29));
   INV_X1 i_61 (.A(b[11]), .ZN(n_30));
   INV_X1 i_62 (.A(b[14]), .ZN(n_31));
   INV_X1 i_63 (.A(b[21]), .ZN(n_32));
   INV_X1 i_64 (.A(b[25]), .ZN(n_33));
endmodule

module datapath__0_1(p_0, a);
   output [31:0]p_0;
   input [31:0]a;

   XOR2_X1 i_0 (.A(a[1]), .B(a[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(a[2]), .B1(a[1]), .B2(a[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(a[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(a[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(a[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(a[6]), .B1(n_27), .B2(a[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(a[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(a[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(a[9]), .B1(n_25), .B2(a[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(a[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(a[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(a[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(a[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(a[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(a[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(a[16]), .B1(n_19), .B2(a[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(a[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(a[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(a[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(a[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(a[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(a[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(a[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(a[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(a[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(a[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(a[27]), .B1(n_9), .B2(a[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(a[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(a[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(a[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(a[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(a[28]), .A3(a[29]), .A4(a[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(a[28]), .A3(a[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(a[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(a[26]), .A3(a[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(a[23]), .A3(a[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(a[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(a[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(a[18]), .A3(a[19]), .A4(a[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(a[18]), .A3(a[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(a[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(a[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(a[15]), .A3(a[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(a[12]), .A3(a[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(a[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(a[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(a[8]), .A3(a[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(a[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(a[5]), .A3(a[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(a[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(a[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(a[2]), .A2(a[1]), .A3(a[0]), .ZN(n_29));
   INV_X1 i_61 (.A(a[11]), .ZN(n_30));
   INV_X1 i_62 (.A(a[14]), .ZN(n_31));
   INV_X1 i_63 (.A(a[21]), .ZN(n_32));
   INV_X1 i_64 (.A(a[25]), .ZN(n_33));
endmodule

module datapath__0_3(A, p_0, multiplicand);
   input [31:0]A;
   output [31:0]p_0;
   input [31:0]multiplicand;

   INV_X1 i_0 (.A(A[0]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_0), .A2(multiplicand[0]), .ZN(n_1));
   OAI21_X1 i_2 (.A(n_1), .B1(multiplicand[0]), .B2(n_0), .ZN(p_0[0]));
   XNOR2_X1 i_3 (.A(A[1]), .B(multiplicand[1]), .ZN(n_2));
   XOR2_X1 i_4 (.A(n_2), .B(n_1), .Z(p_0[1]));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   INV_X1 i_6 (.A(A[1]), .ZN(n_4));
   AOI22_X1 i_7 (.A1(n_2), .A2(n_3), .B1(n_4), .B2(multiplicand[1]), .ZN(n_5));
   XOR2_X1 i_8 (.A(multiplicand[2]), .B(A[2]), .Z(n_6));
   XNOR2_X1 i_9 (.A(n_5), .B(n_6), .ZN(p_0[2]));
   INV_X1 i_10 (.A(multiplicand[2]), .ZN(n_7));
   OAI22_X1 i_11 (.A1(n_5), .A2(n_6), .B1(n_7), .B2(A[2]), .ZN(n_8));
   XNOR2_X1 i_12 (.A(A[3]), .B(multiplicand[3]), .ZN(n_9));
   XNOR2_X1 i_13 (.A(n_8), .B(n_9), .ZN(p_0[3]));
   INV_X1 i_14 (.A(A[3]), .ZN(n_10));
   AOI22_X1 i_15 (.A1(n_8), .A2(n_9), .B1(n_10), .B2(multiplicand[3]), .ZN(n_11));
   XOR2_X1 i_16 (.A(multiplicand[4]), .B(A[4]), .Z(n_12));
   XNOR2_X1 i_17 (.A(n_11), .B(n_12), .ZN(p_0[4]));
   INV_X1 i_18 (.A(multiplicand[4]), .ZN(n_13));
   OAI22_X1 i_19 (.A1(n_11), .A2(n_12), .B1(n_13), .B2(A[4]), .ZN(n_14));
   XNOR2_X1 i_20 (.A(A[5]), .B(multiplicand[5]), .ZN(n_15));
   XNOR2_X1 i_21 (.A(n_14), .B(n_15), .ZN(p_0[5]));
   INV_X1 i_22 (.A(A[5]), .ZN(n_16));
   AOI22_X1 i_23 (.A1(n_14), .A2(n_15), .B1(n_16), .B2(multiplicand[5]), 
      .ZN(n_17));
   XOR2_X1 i_24 (.A(multiplicand[6]), .B(A[6]), .Z(n_18));
   XNOR2_X1 i_25 (.A(n_17), .B(n_18), .ZN(p_0[6]));
   INV_X1 i_26 (.A(multiplicand[6]), .ZN(n_19));
   OAI22_X1 i_27 (.A1(n_17), .A2(n_18), .B1(n_19), .B2(A[6]), .ZN(n_20));
   XNOR2_X1 i_28 (.A(A[7]), .B(multiplicand[7]), .ZN(n_21));
   XNOR2_X1 i_29 (.A(n_20), .B(n_21), .ZN(p_0[7]));
   INV_X1 i_30 (.A(A[7]), .ZN(n_22));
   AOI22_X1 i_31 (.A1(n_20), .A2(n_21), .B1(n_22), .B2(multiplicand[7]), 
      .ZN(n_23));
   XOR2_X1 i_32 (.A(multiplicand[8]), .B(A[8]), .Z(n_24));
   XNOR2_X1 i_33 (.A(n_23), .B(n_24), .ZN(p_0[8]));
   INV_X1 i_34 (.A(multiplicand[8]), .ZN(n_25));
   OAI22_X1 i_35 (.A1(n_23), .A2(n_24), .B1(n_25), .B2(A[8]), .ZN(n_26));
   XNOR2_X1 i_36 (.A(A[9]), .B(multiplicand[9]), .ZN(n_27));
   XNOR2_X1 i_37 (.A(n_26), .B(n_27), .ZN(p_0[9]));
   INV_X1 i_38 (.A(A[9]), .ZN(n_28));
   AOI22_X1 i_39 (.A1(n_26), .A2(n_27), .B1(n_28), .B2(multiplicand[9]), 
      .ZN(n_29));
   XOR2_X1 i_40 (.A(multiplicand[10]), .B(A[10]), .Z(n_30));
   XNOR2_X1 i_41 (.A(n_29), .B(n_30), .ZN(p_0[10]));
   INV_X1 i_42 (.A(multiplicand[10]), .ZN(n_31));
   OAI22_X1 i_43 (.A1(n_29), .A2(n_30), .B1(n_31), .B2(A[10]), .ZN(n_32));
   XNOR2_X1 i_44 (.A(A[11]), .B(multiplicand[11]), .ZN(n_33));
   XNOR2_X1 i_45 (.A(n_32), .B(n_33), .ZN(p_0[11]));
   INV_X1 i_46 (.A(A[11]), .ZN(n_34));
   AOI22_X1 i_47 (.A1(n_32), .A2(n_33), .B1(n_34), .B2(multiplicand[11]), 
      .ZN(n_35));
   XOR2_X1 i_48 (.A(multiplicand[12]), .B(A[12]), .Z(n_36));
   XNOR2_X1 i_49 (.A(n_35), .B(n_36), .ZN(p_0[12]));
   INV_X1 i_50 (.A(multiplicand[12]), .ZN(n_37));
   OAI22_X1 i_51 (.A1(n_35), .A2(n_36), .B1(n_37), .B2(A[12]), .ZN(n_38));
   XNOR2_X1 i_52 (.A(A[13]), .B(multiplicand[13]), .ZN(n_39));
   XNOR2_X1 i_53 (.A(n_38), .B(n_39), .ZN(p_0[13]));
   INV_X1 i_54 (.A(A[13]), .ZN(n_40));
   AOI22_X1 i_55 (.A1(n_38), .A2(n_39), .B1(n_40), .B2(multiplicand[13]), 
      .ZN(n_41));
   XOR2_X1 i_56 (.A(multiplicand[14]), .B(A[14]), .Z(n_42));
   XNOR2_X1 i_57 (.A(n_41), .B(n_42), .ZN(p_0[14]));
   INV_X1 i_58 (.A(multiplicand[14]), .ZN(n_43));
   OAI22_X1 i_59 (.A1(n_41), .A2(n_42), .B1(n_43), .B2(A[14]), .ZN(n_44));
   XNOR2_X1 i_60 (.A(A[15]), .B(multiplicand[15]), .ZN(n_45));
   XNOR2_X1 i_61 (.A(n_44), .B(n_45), .ZN(p_0[15]));
   INV_X1 i_62 (.A(A[15]), .ZN(n_46));
   AOI22_X1 i_63 (.A1(n_44), .A2(n_45), .B1(n_46), .B2(multiplicand[15]), 
      .ZN(n_47));
   XOR2_X1 i_64 (.A(multiplicand[16]), .B(A[16]), .Z(n_48));
   XNOR2_X1 i_65 (.A(n_47), .B(n_48), .ZN(p_0[16]));
   INV_X1 i_66 (.A(multiplicand[16]), .ZN(n_49));
   OAI22_X1 i_67 (.A1(n_47), .A2(n_48), .B1(n_49), .B2(A[16]), .ZN(n_50));
   XNOR2_X1 i_68 (.A(A[17]), .B(multiplicand[17]), .ZN(n_51));
   XNOR2_X1 i_69 (.A(n_50), .B(n_51), .ZN(p_0[17]));
   INV_X1 i_70 (.A(A[17]), .ZN(n_52));
   AOI22_X1 i_71 (.A1(n_50), .A2(n_51), .B1(n_52), .B2(multiplicand[17]), 
      .ZN(n_53));
   XOR2_X1 i_72 (.A(multiplicand[18]), .B(A[18]), .Z(n_54));
   XNOR2_X1 i_73 (.A(n_53), .B(n_54), .ZN(p_0[18]));
   INV_X1 i_74 (.A(multiplicand[18]), .ZN(n_55));
   OAI22_X1 i_75 (.A1(n_53), .A2(n_54), .B1(n_55), .B2(A[18]), .ZN(n_56));
   XNOR2_X1 i_76 (.A(A[19]), .B(multiplicand[19]), .ZN(n_57));
   XNOR2_X1 i_77 (.A(n_56), .B(n_57), .ZN(p_0[19]));
   INV_X1 i_78 (.A(A[19]), .ZN(n_58));
   AOI22_X1 i_79 (.A1(n_56), .A2(n_57), .B1(n_58), .B2(multiplicand[19]), 
      .ZN(n_59));
   XOR2_X1 i_80 (.A(multiplicand[20]), .B(A[20]), .Z(n_60));
   XNOR2_X1 i_81 (.A(n_59), .B(n_60), .ZN(p_0[20]));
   INV_X1 i_82 (.A(multiplicand[20]), .ZN(n_61));
   OAI22_X1 i_83 (.A1(n_59), .A2(n_60), .B1(n_61), .B2(A[20]), .ZN(n_62));
   XNOR2_X1 i_84 (.A(A[21]), .B(multiplicand[21]), .ZN(n_63));
   XNOR2_X1 i_85 (.A(n_62), .B(n_63), .ZN(p_0[21]));
   INV_X1 i_86 (.A(A[21]), .ZN(n_64));
   AOI22_X1 i_87 (.A1(n_62), .A2(n_63), .B1(n_64), .B2(multiplicand[21]), 
      .ZN(n_65));
   XOR2_X1 i_88 (.A(multiplicand[22]), .B(A[22]), .Z(n_66));
   XNOR2_X1 i_89 (.A(n_65), .B(n_66), .ZN(p_0[22]));
   INV_X1 i_90 (.A(multiplicand[22]), .ZN(n_67));
   OAI22_X1 i_91 (.A1(n_65), .A2(n_66), .B1(n_67), .B2(A[22]), .ZN(n_68));
   XNOR2_X1 i_92 (.A(A[23]), .B(multiplicand[23]), .ZN(n_69));
   XNOR2_X1 i_93 (.A(n_68), .B(n_69), .ZN(p_0[23]));
   INV_X1 i_94 (.A(A[23]), .ZN(n_70));
   AOI22_X1 i_95 (.A1(n_68), .A2(n_69), .B1(n_70), .B2(multiplicand[23]), 
      .ZN(n_71));
   XOR2_X1 i_96 (.A(multiplicand[24]), .B(A[24]), .Z(n_72));
   XNOR2_X1 i_97 (.A(n_71), .B(n_72), .ZN(p_0[24]));
   INV_X1 i_98 (.A(multiplicand[24]), .ZN(n_73));
   OAI22_X1 i_99 (.A1(n_71), .A2(n_72), .B1(n_73), .B2(A[24]), .ZN(n_74));
   XNOR2_X1 i_100 (.A(A[25]), .B(multiplicand[25]), .ZN(n_75));
   XNOR2_X1 i_101 (.A(n_74), .B(n_75), .ZN(p_0[25]));
   INV_X1 i_102 (.A(A[25]), .ZN(n_76));
   AOI22_X1 i_103 (.A1(n_74), .A2(n_75), .B1(n_76), .B2(multiplicand[25]), 
      .ZN(n_77));
   XOR2_X1 i_104 (.A(multiplicand[26]), .B(A[26]), .Z(n_78));
   XNOR2_X1 i_105 (.A(n_77), .B(n_78), .ZN(p_0[26]));
   INV_X1 i_106 (.A(multiplicand[26]), .ZN(n_79));
   OAI22_X1 i_107 (.A1(n_77), .A2(n_78), .B1(n_79), .B2(A[26]), .ZN(n_80));
   XNOR2_X1 i_108 (.A(A[27]), .B(multiplicand[27]), .ZN(n_81));
   XNOR2_X1 i_109 (.A(n_80), .B(n_81), .ZN(p_0[27]));
   INV_X1 i_110 (.A(A[27]), .ZN(n_82));
   AOI22_X1 i_111 (.A1(n_80), .A2(n_81), .B1(n_82), .B2(multiplicand[27]), 
      .ZN(n_83));
   XOR2_X1 i_112 (.A(multiplicand[28]), .B(A[28]), .Z(n_84));
   XNOR2_X1 i_113 (.A(n_83), .B(n_84), .ZN(p_0[28]));
   INV_X1 i_114 (.A(multiplicand[28]), .ZN(n_85));
   OAI22_X1 i_115 (.A1(n_83), .A2(n_84), .B1(n_85), .B2(A[28]), .ZN(n_86));
   XNOR2_X1 i_116 (.A(A[29]), .B(multiplicand[29]), .ZN(n_87));
   XNOR2_X1 i_117 (.A(n_86), .B(n_87), .ZN(p_0[29]));
   INV_X1 i_118 (.A(A[29]), .ZN(n_88));
   AOI22_X1 i_119 (.A1(n_86), .A2(n_87), .B1(n_88), .B2(multiplicand[29]), 
      .ZN(n_89));
   INV_X1 i_120 (.A(multiplicand[30]), .ZN(n_90));
   OR2_X1 i_121 (.A1(n_90), .A2(A[30]), .ZN(n_91));
   NAND2_X1 i_122 (.A1(n_90), .A2(A[30]), .ZN(n_92));
   NAND2_X1 i_123 (.A1(n_91), .A2(n_92), .ZN(n_93));
   XNOR2_X1 i_124 (.A(n_89), .B(n_93), .ZN(p_0[30]));
   INV_X1 i_125 (.A(n_92), .ZN(n_94));
   AOI21_X1 i_126 (.A(n_94), .B1(n_89), .B2(n_91), .ZN(n_95));
   XNOR2_X1 i_127 (.A(A[31]), .B(multiplicand[31]), .ZN(n_96));
   XNOR2_X1 i_128 (.A(n_95), .B(n_96), .ZN(p_0[31]));
endmodule

module datapath__0_4(multiplicand, A, p_0);
   input [31:0]multiplicand;
   input [31:0]A;
   output [31:0]p_0;

   HA_X1 i_0 (.A(multiplicand[0]), .B(A[0]), .CO(n_0), .S(p_0[0]));
   FA_X1 i_1 (.A(multiplicand[1]), .B(A[1]), .CI(n_0), .CO(n_1), .S(p_0[1]));
   FA_X1 i_2 (.A(multiplicand[2]), .B(A[2]), .CI(n_1), .CO(n_2), .S(p_0[2]));
   FA_X1 i_3 (.A(multiplicand[3]), .B(A[3]), .CI(n_2), .CO(n_3), .S(p_0[3]));
   FA_X1 i_4 (.A(multiplicand[4]), .B(A[4]), .CI(n_3), .CO(n_4), .S(p_0[4]));
   FA_X1 i_5 (.A(multiplicand[5]), .B(A[5]), .CI(n_4), .CO(n_5), .S(p_0[5]));
   FA_X1 i_6 (.A(multiplicand[6]), .B(A[6]), .CI(n_5), .CO(n_6), .S(p_0[6]));
   FA_X1 i_7 (.A(multiplicand[7]), .B(A[7]), .CI(n_6), .CO(n_7), .S(p_0[7]));
   FA_X1 i_8 (.A(multiplicand[8]), .B(A[8]), .CI(n_7), .CO(n_8), .S(p_0[8]));
   FA_X1 i_9 (.A(multiplicand[9]), .B(A[9]), .CI(n_8), .CO(n_9), .S(p_0[9]));
   FA_X1 i_10 (.A(multiplicand[10]), .B(A[10]), .CI(n_9), .CO(n_10), .S(p_0[10]));
   FA_X1 i_11 (.A(multiplicand[11]), .B(A[11]), .CI(n_10), .CO(n_11), .S(p_0[11]));
   FA_X1 i_12 (.A(multiplicand[12]), .B(A[12]), .CI(n_11), .CO(n_12), .S(p_0[12]));
   FA_X1 i_13 (.A(multiplicand[13]), .B(A[13]), .CI(n_12), .CO(n_13), .S(p_0[13]));
   FA_X1 i_14 (.A(multiplicand[14]), .B(A[14]), .CI(n_13), .CO(n_14), .S(p_0[14]));
   FA_X1 i_15 (.A(multiplicand[15]), .B(A[15]), .CI(n_14), .CO(n_15), .S(p_0[15]));
   FA_X1 i_16 (.A(multiplicand[16]), .B(A[16]), .CI(n_15), .CO(n_16), .S(p_0[16]));
   FA_X1 i_17 (.A(multiplicand[17]), .B(A[17]), .CI(n_16), .CO(n_17), .S(p_0[17]));
   FA_X1 i_18 (.A(multiplicand[18]), .B(A[18]), .CI(n_17), .CO(n_18), .S(p_0[18]));
   FA_X1 i_19 (.A(multiplicand[19]), .B(A[19]), .CI(n_18), .CO(n_19), .S(p_0[19]));
   FA_X1 i_20 (.A(multiplicand[20]), .B(A[20]), .CI(n_19), .CO(n_20), .S(p_0[20]));
   FA_X1 i_21 (.A(multiplicand[21]), .B(A[21]), .CI(n_20), .CO(n_21), .S(p_0[21]));
   FA_X1 i_22 (.A(multiplicand[22]), .B(A[22]), .CI(n_21), .CO(n_22), .S(p_0[22]));
   FA_X1 i_23 (.A(multiplicand[23]), .B(A[23]), .CI(n_22), .CO(n_23), .S(p_0[23]));
   FA_X1 i_24 (.A(multiplicand[24]), .B(A[24]), .CI(n_23), .CO(n_24), .S(p_0[24]));
   FA_X1 i_25 (.A(multiplicand[25]), .B(A[25]), .CI(n_24), .CO(n_25), .S(p_0[25]));
   FA_X1 i_26 (.A(multiplicand[26]), .B(A[26]), .CI(n_25), .CO(n_26), .S(p_0[26]));
   FA_X1 i_27 (.A(multiplicand[27]), .B(A[27]), .CI(n_26), .CO(n_27), .S(p_0[27]));
   FA_X1 i_28 (.A(multiplicand[28]), .B(A[28]), .CI(n_27), .CO(n_28), .S(p_0[28]));
   FA_X1 i_29 (.A(multiplicand[29]), .B(A[29]), .CI(n_28), .CO(n_29), .S(p_0[29]));
   FA_X1 i_30 (.A(multiplicand[30]), .B(A[30]), .CI(n_29), .CO(n_30), .S(p_0[30]));
   XNOR2_X1 i_31 (.A(multiplicand[31]), .B(A[31]), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(p_0[31]));
endmodule

module datapath__0_7(p_0, p_1);
   output [63:0]p_0;
   input [63:0]p_1;

   XOR2_X1 i_0 (.A(p_1[1]), .B(p_1[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_60), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(p_1[2]), .B1(p_1[1]), .B2(p_1[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_1[3]), .B(n_60), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(p_1[4]), .B(n_59), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(p_1[5]), .B(n_58), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_57), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(p_1[6]), .B1(n_58), .B2(p_1[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_1[7]), .B(n_57), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(p_1[8]), .B(n_56), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_55), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(p_1[9]), .B1(n_56), .B2(p_1[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_1[10]), .B(n_55), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(p_1[11]), .B(n_54), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(p_1[12]), .B(n_53), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(p_1[13]), .B(n_52), .ZN(p_0[13]));
   XOR2_X1 i_16 (.A(p_1[14]), .B(n_51), .Z(p_0[14]));
   AND2_X1 i_17 (.A1(n_50), .A2(n_3), .ZN(p_0[15]));
   OAI21_X1 i_18 (.A(p_1[15]), .B1(n_51), .B2(p_1[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(p_1[16]), .B(n_50), .Z(p_0[16]));
   XOR2_X1 i_20 (.A(p_1[17]), .B(n_49), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(p_1[18]), .B(n_48), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(p_1[19]), .B(n_47), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(p_1[20]), .B(n_46), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(p_1[21]), .B(n_45), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(p_1[22]), .B(n_44), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(p_1[23]), .B(n_43), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(p_1[24]), .B(n_42), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(p_1[25]), .B(n_41), .ZN(p_0[25]));
   XNOR2_X1 i_29 (.A(p_1[26]), .B(n_40), .ZN(p_0[26]));
   XOR2_X1 i_30 (.A(p_1[27]), .B(n_39), .Z(p_0[27]));
   XOR2_X1 i_31 (.A(p_1[28]), .B(n_38), .Z(p_0[28]));
   XNOR2_X1 i_32 (.A(p_1[29]), .B(n_37), .ZN(p_0[29]));
   XNOR2_X1 i_33 (.A(p_1[30]), .B(n_36), .ZN(p_0[30]));
   XNOR2_X1 i_34 (.A(p_1[31]), .B(n_35), .ZN(p_0[31]));
   XOR2_X1 i_35 (.A(p_1[32]), .B(n_34), .Z(p_0[32]));
   XOR2_X1 i_36 (.A(p_1[33]), .B(n_33), .Z(p_0[33]));
   XNOR2_X1 i_37 (.A(p_1[34]), .B(n_32), .ZN(p_0[34]));
   XNOR2_X1 i_38 (.A(p_1[35]), .B(n_31), .ZN(p_0[35]));
   XNOR2_X1 i_39 (.A(p_1[36]), .B(n_30), .ZN(p_0[36]));
   XOR2_X1 i_40 (.A(p_1[37]), .B(n_29), .Z(p_0[37]));
   XOR2_X1 i_41 (.A(p_1[38]), .B(n_28), .Z(p_0[38]));
   XNOR2_X1 i_42 (.A(p_1[39]), .B(n_27), .ZN(p_0[39]));
   XNOR2_X1 i_43 (.A(p_1[40]), .B(n_26), .ZN(p_0[40]));
   XOR2_X1 i_44 (.A(p_1[41]), .B(n_25), .Z(p_0[41]));
   XNOR2_X1 i_45 (.A(p_1[42]), .B(n_24), .ZN(p_0[42]));
   XOR2_X1 i_46 (.A(p_1[43]), .B(n_23), .Z(p_0[43]));
   AND2_X1 i_47 (.A1(n_22), .A2(n_4), .ZN(p_0[44]));
   OAI21_X1 i_48 (.A(p_1[44]), .B1(n_23), .B2(p_1[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(p_1[45]), .B(n_22), .Z(p_0[45]));
   XOR2_X1 i_50 (.A(p_1[46]), .B(n_21), .Z(p_0[46]));
   XOR2_X1 i_51 (.A(p_1[47]), .B(n_20), .Z(p_0[47]));
   XOR2_X1 i_52 (.A(p_1[48]), .B(n_19), .Z(p_0[48]));
   XNOR2_X1 i_53 (.A(p_1[49]), .B(n_18), .ZN(p_0[49]));
   XNOR2_X1 i_54 (.A(p_1[50]), .B(n_17), .ZN(p_0[50]));
   XNOR2_X1 i_55 (.A(p_1[51]), .B(n_16), .ZN(p_0[51]));
   XOR2_X1 i_56 (.A(p_1[52]), .B(n_15), .Z(p_0[52]));
   XNOR2_X1 i_57 (.A(p_1[53]), .B(n_14), .ZN(p_0[53]));
   XNOR2_X1 i_58 (.A(p_1[54]), .B(n_13), .ZN(p_0[54]));
   XNOR2_X1 i_59 (.A(p_1[55]), .B(n_12), .ZN(p_0[55]));
   XOR2_X1 i_60 (.A(p_1[56]), .B(n_11), .Z(p_0[56]));
   AND2_X1 i_61 (.A1(n_10), .A2(n_5), .ZN(p_0[57]));
   OAI21_X1 i_62 (.A(p_1[57]), .B1(n_11), .B2(p_1[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(p_1[58]), .B(n_10), .Z(p_0[58]));
   XNOR2_X1 i_64 (.A(p_1[59]), .B(n_9), .ZN(p_0[59]));
   XNOR2_X1 i_65 (.A(p_1[60]), .B(n_8), .ZN(p_0[60]));
   XOR2_X1 i_66 (.A(p_1[61]), .B(n_7), .Z(p_0[61]));
   XNOR2_X1 i_67 (.A(p_1[62]), .B(n_6), .ZN(p_0[62]));
   NAND2_X1 i_68 (.A1(n_6), .A2(n_72), .ZN(p_0[63]));
   NOR2_X1 i_69 (.A1(n_7), .A2(p_1[61]), .ZN(n_6));
   NAND2_X1 i_70 (.A1(n_8), .A2(n_71), .ZN(n_7));
   NOR3_X1 i_71 (.A1(n_10), .A2(p_1[58]), .A3(p_1[59]), .ZN(n_8));
   NOR2_X1 i_72 (.A1(n_10), .A2(p_1[58]), .ZN(n_9));
   OR3_X1 i_73 (.A1(n_11), .A2(p_1[56]), .A3(p_1[57]), .ZN(n_10));
   NAND2_X1 i_74 (.A1(n_12), .A2(n_70), .ZN(n_11));
   NOR4_X1 i_75 (.A1(n_15), .A2(p_1[52]), .A3(p_1[53]), .A4(p_1[54]), .ZN(n_12));
   NOR3_X1 i_76 (.A1(n_15), .A2(p_1[52]), .A3(p_1[53]), .ZN(n_13));
   NOR2_X1 i_77 (.A1(n_15), .A2(p_1[52]), .ZN(n_14));
   NAND2_X1 i_78 (.A1(n_16), .A2(n_69), .ZN(n_15));
   NOR4_X1 i_79 (.A1(n_19), .A2(p_1[48]), .A3(p_1[49]), .A4(p_1[50]), .ZN(n_16));
   NOR3_X1 i_80 (.A1(n_19), .A2(p_1[48]), .A3(p_1[49]), .ZN(n_17));
   NOR2_X1 i_81 (.A1(n_19), .A2(p_1[48]), .ZN(n_18));
   OR2_X1 i_82 (.A1(n_20), .A2(p_1[47]), .ZN(n_19));
   OR2_X1 i_83 (.A1(n_21), .A2(p_1[46]), .ZN(n_20));
   OR2_X1 i_84 (.A1(n_22), .A2(p_1[45]), .ZN(n_21));
   OR3_X1 i_85 (.A1(n_23), .A2(p_1[43]), .A3(p_1[44]), .ZN(n_22));
   NAND2_X1 i_86 (.A1(n_24), .A2(n_68), .ZN(n_23));
   NOR2_X1 i_87 (.A1(n_25), .A2(p_1[41]), .ZN(n_24));
   NAND2_X1 i_88 (.A1(n_26), .A2(n_67), .ZN(n_25));
   NOR3_X1 i_89 (.A1(n_28), .A2(p_1[38]), .A3(p_1[39]), .ZN(n_26));
   NOR2_X1 i_90 (.A1(n_28), .A2(p_1[38]), .ZN(n_27));
   OR2_X1 i_91 (.A1(n_29), .A2(p_1[37]), .ZN(n_28));
   NAND2_X1 i_92 (.A1(n_30), .A2(n_66), .ZN(n_29));
   NOR4_X1 i_93 (.A1(n_33), .A2(p_1[33]), .A3(p_1[34]), .A4(p_1[35]), .ZN(n_30));
   NOR3_X1 i_94 (.A1(n_33), .A2(p_1[33]), .A3(p_1[34]), .ZN(n_31));
   NOR2_X1 i_95 (.A1(n_33), .A2(p_1[33]), .ZN(n_32));
   OR2_X1 i_96 (.A1(n_34), .A2(p_1[32]), .ZN(n_33));
   NAND2_X1 i_97 (.A1(n_35), .A2(n_65), .ZN(n_34));
   NOR4_X1 i_98 (.A1(n_38), .A2(p_1[28]), .A3(p_1[29]), .A4(p_1[30]), .ZN(n_35));
   NOR3_X1 i_99 (.A1(n_38), .A2(p_1[28]), .A3(p_1[29]), .ZN(n_36));
   NOR2_X1 i_100 (.A1(n_38), .A2(p_1[28]), .ZN(n_37));
   OR2_X1 i_101 (.A1(n_39), .A2(p_1[27]), .ZN(n_38));
   NAND2_X1 i_102 (.A1(n_40), .A2(n_64), .ZN(n_39));
   NOR4_X1 i_103 (.A1(n_43), .A2(p_1[23]), .A3(p_1[24]), .A4(p_1[25]), .ZN(n_40));
   NOR3_X1 i_104 (.A1(n_43), .A2(p_1[23]), .A3(p_1[24]), .ZN(n_41));
   NOR2_X1 i_105 (.A1(n_43), .A2(p_1[23]), .ZN(n_42));
   OR2_X1 i_106 (.A1(n_44), .A2(p_1[22]), .ZN(n_43));
   NAND2_X1 i_107 (.A1(n_45), .A2(n_63), .ZN(n_44));
   NOR4_X1 i_108 (.A1(n_48), .A2(p_1[18]), .A3(p_1[19]), .A4(p_1[20]), .ZN(n_45));
   NOR3_X1 i_109 (.A1(n_48), .A2(p_1[18]), .A3(p_1[19]), .ZN(n_46));
   NOR2_X1 i_110 (.A1(n_48), .A2(p_1[18]), .ZN(n_47));
   OR2_X1 i_111 (.A1(n_49), .A2(p_1[17]), .ZN(n_48));
   OR2_X1 i_112 (.A1(n_50), .A2(p_1[16]), .ZN(n_49));
   OR3_X1 i_113 (.A1(n_51), .A2(p_1[14]), .A3(p_1[15]), .ZN(n_50));
   NAND2_X1 i_114 (.A1(n_52), .A2(n_62), .ZN(n_51));
   NOR2_X1 i_115 (.A1(n_53), .A2(p_1[12]), .ZN(n_52));
   NAND2_X1 i_116 (.A1(n_54), .A2(n_61), .ZN(n_53));
   NOR2_X1 i_117 (.A1(n_55), .A2(p_1[10]), .ZN(n_54));
   OR3_X1 i_118 (.A1(n_56), .A2(p_1[8]), .A3(p_1[9]), .ZN(n_55));
   OR2_X1 i_119 (.A1(n_57), .A2(p_1[7]), .ZN(n_56));
   OR3_X1 i_120 (.A1(n_58), .A2(p_1[5]), .A3(p_1[6]), .ZN(n_57));
   OR2_X1 i_121 (.A1(n_59), .A2(p_1[4]), .ZN(n_58));
   OR2_X1 i_122 (.A1(n_60), .A2(p_1[3]), .ZN(n_59));
   OR3_X1 i_123 (.A1(p_1[2]), .A2(p_1[1]), .A3(p_1[0]), .ZN(n_60));
   INV_X1 i_124 (.A(p_1[11]), .ZN(n_61));
   INV_X1 i_125 (.A(p_1[13]), .ZN(n_62));
   INV_X1 i_126 (.A(p_1[21]), .ZN(n_63));
   INV_X1 i_127 (.A(p_1[26]), .ZN(n_64));
   INV_X1 i_128 (.A(p_1[31]), .ZN(n_65));
   INV_X1 i_129 (.A(p_1[36]), .ZN(n_66));
   INV_X1 i_130 (.A(p_1[40]), .ZN(n_67));
   INV_X1 i_131 (.A(p_1[42]), .ZN(n_68));
   INV_X1 i_132 (.A(p_1[51]), .ZN(n_69));
   INV_X1 i_133 (.A(p_1[55]), .ZN(n_70));
   INV_X1 i_134 (.A(p_1[60]), .ZN(n_71));
   INV_X1 i_135 (.A(p_1[62]), .ZN(n_72));
endmodule

module booth_multiplier(clk, rst, a, b, c);
   input clk;
   input rst;
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   wire n_0_0;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire [6:0]SC;
   wire [31:0]A;
   wire [31:0]multiplicand;
   wire [32:0]Q;
   wire out_sign;
   wire n_0_191;
   wire n_0_1;
   wire n_0_2_5;
   wire n_0_2_0;
   wire n_0_2_6;
   wire n_0_2_1;
   wire n_0_2_7;
   wire n_0_2_2;
   wire n_0_2_8;
   wire n_0_2_3;
   wire n_0_2_9;
   wire n_0_2_4;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_2_10;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_2_11;
   wire n_0_231;
   wire n_0_2_12;
   wire n_0_232;
   wire n_0_2_13;
   wire n_0_233;
   wire n_0_2_14;
   wire n_0_234;
   wire n_0_2_15;
   wire n_0_235;
   wire n_0_2_16;
   wire n_0_236;
   wire n_0_2_17;
   wire n_0_237;
   wire n_0_2_18;
   wire n_0_238;
   wire n_0_2_19;
   wire n_0_239;
   wire n_0_2_20;
   wire n_0_240;
   wire n_0_2_21;
   wire n_0_241;
   wire n_0_2_22;
   wire n_0_242;
   wire n_0_2_23;
   wire n_0_243;
   wire n_0_2_24;
   wire n_0_244;
   wire n_0_2_25;
   wire n_0_245;
   wire n_0_2_26;
   wire n_0_246;
   wire n_0_2_27;
   wire n_0_247;
   wire n_0_2_28;
   wire n_0_248;
   wire n_0_2_29;
   wire n_0_249;
   wire n_0_2_30;
   wire n_0_250;
   wire n_0_2_31;
   wire n_0_251;
   wire n_0_2_32;
   wire n_0_252;
   wire n_0_2_33;
   wire n_0_253;
   wire n_0_2_34;
   wire n_0_254;
   wire n_0_2_35;
   wire n_0_255;
   wire n_0_2_36;
   wire n_0_256;
   wire n_0_2_37;
   wire n_0_257;
   wire n_0_2_38;
   wire n_0_258;
   wire n_0_2_39;
   wire n_0_259;
   wire n_0_2_40;
   wire n_0_260;
   wire n_0_2_41;
   wire n_0_261;
   wire n_0_2_42;
   wire n_0_262;
   wire n_0_2_43;
   wire n_0_2_44;
   wire n_0_2_45;
   wire n_0_2_46;
   wire n_0_263;
   wire n_0_2_47;
   wire n_0_264;
   wire n_0_2_48;
   wire n_0_265;
   wire n_0_2_49;
   wire n_0_266;
   wire n_0_2_50;
   wire n_0_267;
   wire n_0_2_51;
   wire n_0_268;
   wire n_0_2_52;
   wire n_0_269;
   wire n_0_2_53;
   wire n_0_270;
   wire n_0_2_54;
   wire n_0_271;
   wire n_0_2_55;
   wire n_0_272;
   wire n_0_2_56;
   wire n_0_273;
   wire n_0_2_57;
   wire n_0_274;
   wire n_0_2_58;
   wire n_0_275;
   wire n_0_2_59;
   wire n_0_276;
   wire n_0_2_60;
   wire n_0_277;
   wire n_0_2_61;
   wire n_0_278;
   wire n_0_2_62;
   wire n_0_279;
   wire n_0_2_63;
   wire n_0_280;
   wire n_0_2_64;
   wire n_0_281;
   wire n_0_2_65;
   wire n_0_282;
   wire n_0_2_66;
   wire n_0_283;
   wire n_0_2_67;
   wire n_0_284;
   wire n_0_2_68;
   wire n_0_285;
   wire n_0_2_69;
   wire n_0_286;
   wire n_0_2_70;
   wire n_0_287;
   wire n_0_2_71;
   wire n_0_288;
   wire n_0_2_72;
   wire n_0_289;
   wire n_0_2_73;
   wire n_0_290;
   wire n_0_2_74;
   wire n_0_291;
   wire n_0_2_75;
   wire n_0_292;
   wire n_0_2_76;
   wire n_0_293;
   wire n_0_2_77;
   wire n_0_294;
   wire n_0_2_78;
   wire n_0_295;
   wire n_0_2_79;
   wire n_0_296;
   wire n_0_2_80;
   wire n_0_297;
   wire n_0_2_81;
   wire n_0_298;
   wire n_0_2_82;
   wire n_0_299;
   wire n_0_2_83;
   wire n_0_300;
   wire n_0_2_84;
   wire n_0_301;
   wire n_0_2_85;
   wire n_0_302;
   wire n_0_2_86;
   wire n_0_303;
   wire n_0_2_87;
   wire n_0_304;
   wire n_0_2_88;
   wire n_0_305;
   wire n_0_2_89;
   wire n_0_306;
   wire n_0_2_90;
   wire n_0_307;
   wire n_0_2_91;
   wire n_0_308;
   wire n_0_2_92;
   wire n_0_309;
   wire n_0_2_93;
   wire n_0_310;
   wire n_0_2_94;
   wire n_0_311;
   wire n_0_2_95;
   wire n_0_312;
   wire n_0_2_96;
   wire n_0_313;
   wire n_0_2_97;
   wire n_0_314;
   wire n_0_2_98;
   wire n_0_315;
   wire n_0_2_99;
   wire n_0_316;
   wire n_0_2_100;
   wire n_0_317;
   wire n_0_2_101;
   wire n_0_318;
   wire n_0_2_102;
   wire n_0_319;
   wire n_0_2_103;
   wire n_0_320;
   wire n_0_2_104;
   wire n_0_321;
   wire n_0_2_105;
   wire n_0_322;
   wire n_0_2_106;
   wire n_0_323;
   wire n_0_2_107;
   wire n_0_324;
   wire n_0_2_108;
   wire n_0_325;
   wire n_0_2_109;
   wire n_0_2_110;
   wire n_0_2_111;
   wire n_0_326;
   wire n_0_2_112;
   wire n_0_2_113;
   wire n_0_328;
   wire n_0_2_114;
   wire n_0_329;
   wire n_0_2_115;
   wire n_0_330;
   wire n_0_2_116;
   wire n_0_331;
   wire n_0_2_117;
   wire n_0_332;
   wire n_0_2_118;
   wire n_0_333;
   wire n_0_2_119;
   wire n_0_334;
   wire n_0_2_120;
   wire n_0_335;
   wire n_0_2_121;
   wire n_0_336;
   wire n_0_2_122;
   wire n_0_337;
   wire n_0_2_123;
   wire n_0_338;
   wire n_0_2_124;
   wire n_0_339;
   wire n_0_2_125;
   wire n_0_340;
   wire n_0_2_126;
   wire n_0_341;
   wire n_0_2_127;
   wire n_0_342;
   wire n_0_2_128;
   wire n_0_343;
   wire n_0_2_129;
   wire n_0_344;
   wire n_0_2_130;
   wire n_0_345;
   wire n_0_2_131;
   wire n_0_346;
   wire n_0_2_132;
   wire n_0_347;
   wire n_0_2_133;
   wire n_0_348;
   wire n_0_2_134;
   wire n_0_349;
   wire n_0_2_135;
   wire n_0_350;
   wire n_0_2_136;
   wire n_0_351;
   wire n_0_2_137;
   wire n_0_352;
   wire n_0_2_138;
   wire n_0_353;
   wire n_0_2_139;
   wire n_0_354;
   wire n_0_2_140;
   wire n_0_355;
   wire n_0_2_141;
   wire n_0_356;
   wire n_0_2_142;
   wire n_0_357;
   wire n_0_2_143;
   wire n_0_2_144;
   wire n_0_358;
   wire n_0_2_145;
   wire n_0_2_146;
   wire n_0_359;
   wire n_0_2_147;
   wire n_0_2_148;
   wire n_0_2_149;
   wire n_0_327;
   wire n_0_2_150;
   wire n_0_2_151;
   wire n_0_2_152;
   wire n_0_2_153;
   wire n_0_2_154;
   wire n_0_2_155;
   wire n_0_2_156;
   wire n_0_2_157;
   wire n_0_2_158;
   wire n_0_2_159;
   wire n_0_2_160;
   wire n_0_2_161;
   wire n_0_2_162;
   wire n_0_2_163;
   wire n_0_2_164;
   wire n_0_2_165;
   wire n_0_2_166;
   wire n_0_2_167;
   wire n_0_2_168;
   wire n_0_2_169;
   wire n_0_2_170;
   wire n_0_2_171;
   wire n_0_2_172;
   wire n_0_2_173;
   wire n_0_2_174;
   wire n_0_2_175;
   wire n_0_2_176;
   wire n_0_2_177;
   wire n_0_2_178;
   wire n_0_2_179;
   wire n_0_2_180;
   wire n_0_2_181;
   wire n_0_2_182;
   wire n_0_2_183;
   wire n_0_2_184;
   wire n_0_2_185;
   wire n_0_2_186;
   wire n_0_2_187;
   wire n_0_2_188;
   wire n_0_2_189;
   wire n_0_192;
   wire n_0_2_190;

   CLKGATETST_X1 clk_gate_c_reg (.CK(clk), .E(n_0_326), .SE(1'b0), .GCK(n_0_0));
   DFF_X1 \c_reg[63]  (.D(n_0_262), .CK(n_0_0), .Q(c[63]), .QN());
   DFF_X1 \c_reg[62]  (.D(n_0_261), .CK(n_0_0), .Q(c[62]), .QN());
   DFF_X1 \c_reg[61]  (.D(n_0_260), .CK(n_0_0), .Q(c[61]), .QN());
   DFF_X1 \c_reg[60]  (.D(n_0_259), .CK(n_0_0), .Q(c[60]), .QN());
   DFF_X1 \c_reg[59]  (.D(n_0_258), .CK(n_0_0), .Q(c[59]), .QN());
   DFF_X1 \c_reg[58]  (.D(n_0_257), .CK(n_0_0), .Q(c[58]), .QN());
   DFF_X1 \c_reg[57]  (.D(n_0_256), .CK(n_0_0), .Q(c[57]), .QN());
   DFF_X1 \c_reg[56]  (.D(n_0_255), .CK(n_0_0), .Q(c[56]), .QN());
   DFF_X1 \c_reg[55]  (.D(n_0_254), .CK(n_0_0), .Q(c[55]), .QN());
   DFF_X1 \c_reg[54]  (.D(n_0_253), .CK(n_0_0), .Q(c[54]), .QN());
   DFF_X1 \c_reg[53]  (.D(n_0_252), .CK(n_0_0), .Q(c[53]), .QN());
   DFF_X1 \c_reg[52]  (.D(n_0_251), .CK(n_0_0), .Q(c[52]), .QN());
   DFF_X1 \c_reg[51]  (.D(n_0_250), .CK(n_0_0), .Q(c[51]), .QN());
   DFF_X1 \c_reg[50]  (.D(n_0_249), .CK(n_0_0), .Q(c[50]), .QN());
   DFF_X1 \c_reg[49]  (.D(n_0_248), .CK(n_0_0), .Q(c[49]), .QN());
   DFF_X1 \c_reg[48]  (.D(n_0_247), .CK(n_0_0), .Q(c[48]), .QN());
   DFF_X1 \c_reg[47]  (.D(n_0_246), .CK(n_0_0), .Q(c[47]), .QN());
   DFF_X1 \c_reg[46]  (.D(n_0_245), .CK(n_0_0), .Q(c[46]), .QN());
   DFF_X1 \c_reg[45]  (.D(n_0_244), .CK(n_0_0), .Q(c[45]), .QN());
   DFF_X1 \c_reg[44]  (.D(n_0_243), .CK(n_0_0), .Q(c[44]), .QN());
   DFF_X1 \c_reg[43]  (.D(n_0_242), .CK(n_0_0), .Q(c[43]), .QN());
   DFF_X1 \c_reg[42]  (.D(n_0_241), .CK(n_0_0), .Q(c[42]), .QN());
   DFF_X1 \c_reg[41]  (.D(n_0_240), .CK(n_0_0), .Q(c[41]), .QN());
   DFF_X1 \c_reg[40]  (.D(n_0_239), .CK(n_0_0), .Q(c[40]), .QN());
   DFF_X1 \c_reg[39]  (.D(n_0_238), .CK(n_0_0), .Q(c[39]), .QN());
   DFF_X1 \c_reg[38]  (.D(n_0_237), .CK(n_0_0), .Q(c[38]), .QN());
   DFF_X1 \c_reg[37]  (.D(n_0_236), .CK(n_0_0), .Q(c[37]), .QN());
   DFF_X1 \c_reg[36]  (.D(n_0_235), .CK(n_0_0), .Q(c[36]), .QN());
   DFF_X1 \c_reg[35]  (.D(n_0_234), .CK(n_0_0), .Q(c[35]), .QN());
   DFF_X1 \c_reg[34]  (.D(n_0_233), .CK(n_0_0), .Q(c[34]), .QN());
   DFF_X1 \c_reg[33]  (.D(n_0_232), .CK(n_0_0), .Q(c[33]), .QN());
   DFF_X1 \c_reg[32]  (.D(n_0_231), .CK(n_0_0), .Q(c[32]), .QN());
   DFF_X1 \c_reg[31]  (.D(n_0_230), .CK(n_0_0), .Q(c[31]), .QN());
   DFF_X1 \c_reg[30]  (.D(n_0_229), .CK(n_0_0), .Q(c[30]), .QN());
   DFF_X1 \c_reg[29]  (.D(n_0_228), .CK(n_0_0), .Q(c[29]), .QN());
   DFF_X1 \c_reg[28]  (.D(n_0_227), .CK(n_0_0), .Q(c[28]), .QN());
   DFF_X1 \c_reg[27]  (.D(n_0_226), .CK(n_0_0), .Q(c[27]), .QN());
   DFF_X1 \c_reg[26]  (.D(n_0_225), .CK(n_0_0), .Q(c[26]), .QN());
   DFF_X1 \c_reg[25]  (.D(n_0_224), .CK(n_0_0), .Q(c[25]), .QN());
   DFF_X1 \c_reg[24]  (.D(n_0_223), .CK(n_0_0), .Q(c[24]), .QN());
   DFF_X1 \c_reg[23]  (.D(n_0_222), .CK(n_0_0), .Q(c[23]), .QN());
   DFF_X1 \c_reg[22]  (.D(n_0_221), .CK(n_0_0), .Q(c[22]), .QN());
   DFF_X1 \c_reg[21]  (.D(n_0_220), .CK(n_0_0), .Q(c[21]), .QN());
   DFF_X1 \c_reg[20]  (.D(n_0_219), .CK(n_0_0), .Q(c[20]), .QN());
   DFF_X1 \c_reg[19]  (.D(n_0_218), .CK(n_0_0), .Q(c[19]), .QN());
   DFF_X1 \c_reg[18]  (.D(n_0_217), .CK(n_0_0), .Q(c[18]), .QN());
   DFF_X1 \c_reg[17]  (.D(n_0_216), .CK(n_0_0), .Q(c[17]), .QN());
   DFF_X1 \c_reg[16]  (.D(n_0_215), .CK(n_0_0), .Q(c[16]), .QN());
   DFF_X1 \c_reg[15]  (.D(n_0_214), .CK(n_0_0), .Q(c[15]), .QN());
   DFF_X1 \c_reg[14]  (.D(n_0_213), .CK(n_0_0), .Q(c[14]), .QN());
   DFF_X1 \c_reg[13]  (.D(n_0_212), .CK(n_0_0), .Q(c[13]), .QN());
   DFF_X1 \c_reg[12]  (.D(n_0_211), .CK(n_0_0), .Q(c[12]), .QN());
   DFF_X1 \c_reg[11]  (.D(n_0_210), .CK(n_0_0), .Q(c[11]), .QN());
   DFF_X1 \c_reg[10]  (.D(n_0_209), .CK(n_0_0), .Q(c[10]), .QN());
   DFF_X1 \c_reg[9]  (.D(n_0_208), .CK(n_0_0), .Q(c[9]), .QN());
   DFF_X1 \c_reg[8]  (.D(n_0_207), .CK(n_0_0), .Q(c[8]), .QN());
   DFF_X1 \c_reg[7]  (.D(n_0_206), .CK(n_0_0), .Q(c[7]), .QN());
   DFF_X1 \c_reg[6]  (.D(n_0_205), .CK(n_0_0), .Q(c[6]), .QN());
   DFF_X1 \c_reg[5]  (.D(n_0_204), .CK(n_0_0), .Q(c[5]), .QN());
   DFF_X1 \c_reg[4]  (.D(n_0_203), .CK(n_0_0), .Q(c[4]), .QN());
   DFF_X1 \c_reg[3]  (.D(n_0_202), .CK(n_0_0), .Q(c[3]), .QN());
   DFF_X1 \c_reg[2]  (.D(n_0_201), .CK(n_0_0), .Q(c[2]), .QN());
   DFF_X1 \c_reg[1]  (.D(n_0_200), .CK(n_0_0), .Q(c[1]), .QN());
   DFF_X1 \c_reg[0]  (.D(n_0_328), .CK(n_0_0), .Q(c[0]), .QN());
   datapath i_0_1 (.p_0({n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
      n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, 
      n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, 
      n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, uc_0}), .b(b));
   datapath__0_1 i_0_3 (.p_0({n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, 
      n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, 
      n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, 
      n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, uc_1}), .a(a));
   datapath__0_3 i_0_5 (.A(A), .p_0({n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, 
      n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, 
      n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, 
      n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64}), 
      .multiplicand({n_0_325, n_0_324, n_0_323, n_0_322, n_0_321, n_0_320, 
      n_0_319, n_0_318, n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, n_0_312, 
      n_0_311, n_0_310, n_0_309, n_0_308, n_0_307, n_0_306, n_0_305, n_0_304, 
      n_0_303, n_0_302, n_0_301, n_0_300, n_0_299, n_0_298, n_0_297, n_0_296, 
      n_0_295, n_0_294}));
   datapath__0_4 i_0_6 (.multiplicand({n_0_325, n_0_324, n_0_323, n_0_322, 
      n_0_321, n_0_320, n_0_319, n_0_318, n_0_317, n_0_316, n_0_315, n_0_314, 
      n_0_313, n_0_312, n_0_311, n_0_310, n_0_309, n_0_308, n_0_307, n_0_306, 
      n_0_305, n_0_304, n_0_303, n_0_302, n_0_301, n_0_300, n_0_299, n_0_298, 
      n_0_297, n_0_296, n_0_295, n_0_294}), .A(A), .p_0({n_0_127, n_0_126, 
      n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, 
      n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, 
      n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, 
      n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96}));
   datapath__0_7 i_0_9 (.p_0({n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, 
      n_0_185, n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, 
      n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, 
      n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, 
      n_0_161, n_0_160, n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, 
      n_0_153, n_0_152, n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, 
      n_0_145, n_0_144, n_0_143, n_0_142, n_0_141, n_0_140, n_0_139, n_0_138, 
      n_0_137, n_0_136, n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, 
      n_0_129, n_0_128, uc_2}), .p_1({1'b0, n_0_293, n_0_292, n_0_291, n_0_290, 
      n_0_289, n_0_288, n_0_287, n_0_286, n_0_285, n_0_284, n_0_283, n_0_282, 
      n_0_281, n_0_280, n_0_279, n_0_278, n_0_277, n_0_276, n_0_275, n_0_274, 
      n_0_273, n_0_272, n_0_271, n_0_270, n_0_269, n_0_268, n_0_267, n_0_266, 
      n_0_265, n_0_264, n_0_263, n_0_359, n_0_358, n_0_357, n_0_356, n_0_355, 
      n_0_354, n_0_353, n_0_352, n_0_351, n_0_350, n_0_349, n_0_348, n_0_347, 
      n_0_346, n_0_345, n_0_344, n_0_343, n_0_342, n_0_341, n_0_340, n_0_339, 
      n_0_338, n_0_337, n_0_336, n_0_335, n_0_334, n_0_333, n_0_332, n_0_331, 
      n_0_330, n_0_329, n_0_328}));
   DFFR_X1 \SC_reg[6]  (.D(n_0_198), .RN(n_0_191), .CK(clk), .Q(SC[6]), .QN());
   DFFR_X1 \SC_reg[5]  (.D(n_0_197), .RN(n_0_191), .CK(clk), .Q(SC[5]), .QN());
   DFFR_X1 \SC_reg[4]  (.D(n_0_196), .RN(n_0_191), .CK(clk), .Q(SC[4]), .QN());
   DFFR_X1 \SC_reg[3]  (.D(n_0_195), .RN(n_0_191), .CK(clk), .Q(SC[3]), .QN());
   DFFR_X1 \SC_reg[2]  (.D(n_0_194), .RN(n_0_191), .CK(clk), .Q(SC[2]), .QN());
   DFFR_X1 \SC_reg[1]  (.D(n_0_193), .RN(n_0_191), .CK(clk), .Q(SC[1]), .QN());
   DFFR_X1 \SC_reg[0]  (.D(n_0_192), .RN(n_0_191), .CK(clk), .Q(SC[0]), .QN());
   DFFR_X1 \A_reg[31]  (.D(n_0_327), .RN(n_0_191), .CK(clk), .Q(A[31]), .QN());
   DFFR_X1 \A_reg[30]  (.D(n_0_293), .RN(n_0_191), .CK(clk), .Q(A[30]), .QN());
   DFFR_X1 \A_reg[29]  (.D(n_0_292), .RN(n_0_191), .CK(clk), .Q(A[29]), .QN());
   DFFR_X1 \A_reg[28]  (.D(n_0_291), .RN(n_0_191), .CK(clk), .Q(A[28]), .QN());
   DFFR_X1 \A_reg[27]  (.D(n_0_290), .RN(n_0_191), .CK(clk), .Q(A[27]), .QN());
   DFFR_X1 \A_reg[26]  (.D(n_0_289), .RN(n_0_191), .CK(clk), .Q(A[26]), .QN());
   DFFR_X1 \A_reg[25]  (.D(n_0_288), .RN(n_0_191), .CK(clk), .Q(A[25]), .QN());
   DFFR_X1 \A_reg[24]  (.D(n_0_287), .RN(n_0_191), .CK(clk), .Q(A[24]), .QN());
   DFFR_X1 \A_reg[23]  (.D(n_0_286), .RN(n_0_191), .CK(clk), .Q(A[23]), .QN());
   DFFR_X1 \A_reg[22]  (.D(n_0_285), .RN(n_0_191), .CK(clk), .Q(A[22]), .QN());
   DFFR_X1 \A_reg[21]  (.D(n_0_284), .RN(n_0_191), .CK(clk), .Q(A[21]), .QN());
   DFFR_X1 \A_reg[20]  (.D(n_0_283), .RN(n_0_191), .CK(clk), .Q(A[20]), .QN());
   DFFR_X1 \A_reg[19]  (.D(n_0_282), .RN(n_0_191), .CK(clk), .Q(A[19]), .QN());
   DFFR_X1 \A_reg[18]  (.D(n_0_281), .RN(n_0_191), .CK(clk), .Q(A[18]), .QN());
   DFFR_X1 \A_reg[17]  (.D(n_0_280), .RN(n_0_191), .CK(clk), .Q(A[17]), .QN());
   DFFR_X1 \A_reg[16]  (.D(n_0_279), .RN(n_0_191), .CK(clk), .Q(A[16]), .QN());
   DFFR_X1 \A_reg[15]  (.D(n_0_278), .RN(n_0_191), .CK(clk), .Q(A[15]), .QN());
   DFFR_X1 \A_reg[14]  (.D(n_0_277), .RN(n_0_191), .CK(clk), .Q(A[14]), .QN());
   DFFR_X1 \A_reg[13]  (.D(n_0_276), .RN(n_0_191), .CK(clk), .Q(A[13]), .QN());
   DFFR_X1 \A_reg[12]  (.D(n_0_275), .RN(n_0_191), .CK(clk), .Q(A[12]), .QN());
   DFFR_X1 \A_reg[11]  (.D(n_0_274), .RN(n_0_191), .CK(clk), .Q(A[11]), .QN());
   DFFR_X1 \A_reg[10]  (.D(n_0_273), .RN(n_0_191), .CK(clk), .Q(A[10]), .QN());
   DFFR_X1 \A_reg[9]  (.D(n_0_272), .RN(n_0_191), .CK(clk), .Q(A[9]), .QN());
   DFFR_X1 \A_reg[8]  (.D(n_0_271), .RN(n_0_191), .CK(clk), .Q(A[8]), .QN());
   DFFR_X1 \A_reg[7]  (.D(n_0_270), .RN(n_0_191), .CK(clk), .Q(A[7]), .QN());
   DFFR_X1 \A_reg[6]  (.D(n_0_269), .RN(n_0_191), .CK(clk), .Q(A[6]), .QN());
   DFFR_X1 \A_reg[5]  (.D(n_0_268), .RN(n_0_191), .CK(clk), .Q(A[5]), .QN());
   DFFR_X1 \A_reg[4]  (.D(n_0_267), .RN(n_0_191), .CK(clk), .Q(A[4]), .QN());
   DFFR_X1 \A_reg[3]  (.D(n_0_266), .RN(n_0_191), .CK(clk), .Q(A[3]), .QN());
   DFFR_X1 \A_reg[2]  (.D(n_0_265), .RN(n_0_191), .CK(clk), .Q(A[2]), .QN());
   DFFR_X1 \A_reg[1]  (.D(n_0_264), .RN(n_0_191), .CK(clk), .Q(A[1]), .QN());
   DFFR_X1 \A_reg[0]  (.D(n_0_263), .RN(n_0_191), .CK(clk), .Q(A[0]), .QN());
   DFF_X1 \multiplicand_reg[31]  (.D(n_0_325), .CK(n_0_1), .Q(multiplicand[31]), 
      .QN());
   DFF_X1 \multiplicand_reg[30]  (.D(n_0_324), .CK(n_0_1), .Q(multiplicand[30]), 
      .QN());
   DFF_X1 \multiplicand_reg[29]  (.D(n_0_323), .CK(n_0_1), .Q(multiplicand[29]), 
      .QN());
   DFF_X1 \multiplicand_reg[28]  (.D(n_0_322), .CK(n_0_1), .Q(multiplicand[28]), 
      .QN());
   DFF_X1 \multiplicand_reg[27]  (.D(n_0_321), .CK(n_0_1), .Q(multiplicand[27]), 
      .QN());
   DFF_X1 \multiplicand_reg[26]  (.D(n_0_320), .CK(n_0_1), .Q(multiplicand[26]), 
      .QN());
   DFF_X1 \multiplicand_reg[25]  (.D(n_0_319), .CK(n_0_1), .Q(multiplicand[25]), 
      .QN());
   DFF_X1 \multiplicand_reg[24]  (.D(n_0_318), .CK(n_0_1), .Q(multiplicand[24]), 
      .QN());
   DFF_X1 \multiplicand_reg[23]  (.D(n_0_317), .CK(n_0_1), .Q(multiplicand[23]), 
      .QN());
   DFF_X1 \multiplicand_reg[22]  (.D(n_0_316), .CK(n_0_1), .Q(multiplicand[22]), 
      .QN());
   DFF_X1 \multiplicand_reg[21]  (.D(n_0_315), .CK(n_0_1), .Q(multiplicand[21]), 
      .QN());
   DFF_X1 \multiplicand_reg[20]  (.D(n_0_314), .CK(n_0_1), .Q(multiplicand[20]), 
      .QN());
   DFF_X1 \multiplicand_reg[19]  (.D(n_0_313), .CK(n_0_1), .Q(multiplicand[19]), 
      .QN());
   DFF_X1 \multiplicand_reg[18]  (.D(n_0_312), .CK(n_0_1), .Q(multiplicand[18]), 
      .QN());
   DFF_X1 \multiplicand_reg[17]  (.D(n_0_311), .CK(n_0_1), .Q(multiplicand[17]), 
      .QN());
   DFF_X1 \multiplicand_reg[16]  (.D(n_0_310), .CK(n_0_1), .Q(multiplicand[16]), 
      .QN());
   DFF_X1 \multiplicand_reg[15]  (.D(n_0_309), .CK(n_0_1), .Q(multiplicand[15]), 
      .QN());
   DFF_X1 \multiplicand_reg[14]  (.D(n_0_308), .CK(n_0_1), .Q(multiplicand[14]), 
      .QN());
   DFF_X1 \multiplicand_reg[13]  (.D(n_0_307), .CK(n_0_1), .Q(multiplicand[13]), 
      .QN());
   DFF_X1 \multiplicand_reg[12]  (.D(n_0_306), .CK(n_0_1), .Q(multiplicand[12]), 
      .QN());
   DFF_X1 \multiplicand_reg[11]  (.D(n_0_305), .CK(n_0_1), .Q(multiplicand[11]), 
      .QN());
   DFF_X1 \multiplicand_reg[10]  (.D(n_0_304), .CK(n_0_1), .Q(multiplicand[10]), 
      .QN());
   DFF_X1 \multiplicand_reg[9]  (.D(n_0_303), .CK(n_0_1), .Q(multiplicand[9]), 
      .QN());
   DFF_X1 \multiplicand_reg[8]  (.D(n_0_302), .CK(n_0_1), .Q(multiplicand[8]), 
      .QN());
   DFF_X1 \multiplicand_reg[7]  (.D(n_0_301), .CK(n_0_1), .Q(multiplicand[7]), 
      .QN());
   DFF_X1 \multiplicand_reg[6]  (.D(n_0_300), .CK(n_0_1), .Q(multiplicand[6]), 
      .QN());
   DFF_X1 \multiplicand_reg[5]  (.D(n_0_299), .CK(n_0_1), .Q(multiplicand[5]), 
      .QN());
   DFF_X1 \multiplicand_reg[4]  (.D(n_0_298), .CK(n_0_1), .Q(multiplicand[4]), 
      .QN());
   DFF_X1 \multiplicand_reg[3]  (.D(n_0_297), .CK(n_0_1), .Q(multiplicand[3]), 
      .QN());
   DFF_X1 \multiplicand_reg[2]  (.D(n_0_296), .CK(n_0_1), .Q(multiplicand[2]), 
      .QN());
   DFF_X1 \multiplicand_reg[1]  (.D(n_0_295), .CK(n_0_1), .Q(multiplicand[1]), 
      .QN());
   DFF_X1 \multiplicand_reg[0]  (.D(n_0_294), .CK(n_0_1), .Q(multiplicand[0]), 
      .QN());
   DFF_X1 \Q_reg[32]  (.D(n_0_359), .CK(n_0_1), .Q(Q[32]), .QN());
   DFF_X1 \Q_reg[31]  (.D(n_0_358), .CK(n_0_1), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_0_357), .CK(n_0_1), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_0_356), .CK(n_0_1), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_0_355), .CK(n_0_1), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_0_354), .CK(n_0_1), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_0_353), .CK(n_0_1), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_0_352), .CK(n_0_1), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_0_351), .CK(n_0_1), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_0_350), .CK(n_0_1), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_0_349), .CK(n_0_1), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_0_348), .CK(n_0_1), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_0_347), .CK(n_0_1), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_0_346), .CK(n_0_1), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_0_345), .CK(n_0_1), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_0_344), .CK(n_0_1), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_0_343), .CK(n_0_1), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_0_342), .CK(n_0_1), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_0_341), .CK(n_0_1), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_0_340), .CK(n_0_1), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_0_339), .CK(n_0_1), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_0_338), .CK(n_0_1), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_0_337), .CK(n_0_1), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_0_336), .CK(n_0_1), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_0_335), .CK(n_0_1), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_0_334), .CK(n_0_1), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_0_333), .CK(n_0_1), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_0_332), .CK(n_0_1), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_0_331), .CK(n_0_1), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_0_330), .CK(n_0_1), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_0_329), .CK(n_0_1), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_0_328), .CK(n_0_1), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0_327), .CK(n_0_1), .Q(Q[0]), .QN());
   DFF_X1 out_sign_reg (.D(n_0_199), .CK(n_0_1), .Q(out_sign), .QN());
   INV_X1 i_0_0_0 (.A(rst), .ZN(n_0_191));
   CLKGATETST_X1 clk_gate_out_sign_reg (.CK(clk), .E(n_0_191), .SE(1'b0), 
      .GCK(n_0_1));
   HA_X1 i_0_2_0 (.A(SC[1]), .B(SC[0]), .CO(n_0_2_0), .S(n_0_2_5));
   HA_X1 i_0_2_1 (.A(SC[2]), .B(n_0_2_0), .CO(n_0_2_1), .S(n_0_2_6));
   HA_X1 i_0_2_2 (.A(SC[3]), .B(n_0_2_1), .CO(n_0_2_2), .S(n_0_2_7));
   HA_X1 i_0_2_3 (.A(SC[4]), .B(n_0_2_2), .CO(n_0_2_3), .S(n_0_2_8));
   HA_X1 i_0_2_4 (.A(SC[5]), .B(n_0_2_3), .CO(n_0_2_4), .S(n_0_2_9));
   AND2_X1 i_0_2_5 (.A1(n_0_2_5), .A2(n_0_2_112), .ZN(n_0_193));
   AND2_X1 i_0_2_6 (.A1(n_0_2_6), .A2(n_0_2_112), .ZN(n_0_194));
   AND2_X1 i_0_2_7 (.A1(n_0_2_7), .A2(n_0_2_112), .ZN(n_0_195));
   AND2_X1 i_0_2_8 (.A1(n_0_2_8), .A2(n_0_2_112), .ZN(n_0_196));
   AND2_X1 i_0_2_9 (.A1(n_0_2_9), .A2(n_0_2_112), .ZN(n_0_197));
   AOI221_X1 i_0_2_10 (.A(n_0_326), .B1(n_0_2_190), .B2(n_0_2_157), .C1(SC[6]), 
      .C2(n_0_2_4), .ZN(n_0_198));
   INV_X1 i_0_2_11 (.A(n_0_2_10), .ZN(n_0_199));
   AOI222_X1 i_0_2_12 (.A1(out_sign), .A2(n_0_2_153), .B1(n_0_2_188), .B2(
      n_0_2_146), .C1(a[31]), .C2(n_0_2_144), .ZN(n_0_2_10));
   AOI22_X1 i_0_2_13 (.A1(n_0_2_158), .A2(n_0_2_43), .B1(n_0_2_115), .B2(
      n_0_2_44), .ZN(n_0_200));
   AOI22_X1 i_0_2_14 (.A1(n_0_2_159), .A2(n_0_2_43), .B1(n_0_2_116), .B2(
      n_0_2_44), .ZN(n_0_201));
   AOI22_X1 i_0_2_15 (.A1(n_0_2_160), .A2(n_0_2_43), .B1(n_0_2_117), .B2(
      n_0_2_44), .ZN(n_0_202));
   AOI22_X1 i_0_2_16 (.A1(n_0_2_161), .A2(n_0_2_43), .B1(n_0_2_118), .B2(
      n_0_2_44), .ZN(n_0_203));
   AOI22_X1 i_0_2_17 (.A1(n_0_2_162), .A2(n_0_2_43), .B1(n_0_2_119), .B2(
      n_0_2_44), .ZN(n_0_204));
   AOI22_X1 i_0_2_18 (.A1(n_0_2_163), .A2(n_0_2_43), .B1(n_0_2_120), .B2(
      n_0_2_44), .ZN(n_0_205));
   AOI22_X1 i_0_2_19 (.A1(n_0_2_164), .A2(n_0_2_43), .B1(n_0_2_121), .B2(
      n_0_2_44), .ZN(n_0_206));
   AOI22_X1 i_0_2_20 (.A1(n_0_2_165), .A2(n_0_2_43), .B1(n_0_2_122), .B2(
      n_0_2_44), .ZN(n_0_207));
   AOI22_X1 i_0_2_21 (.A1(n_0_2_166), .A2(n_0_2_43), .B1(n_0_2_123), .B2(
      n_0_2_44), .ZN(n_0_208));
   AOI22_X1 i_0_2_22 (.A1(n_0_2_167), .A2(n_0_2_43), .B1(n_0_2_124), .B2(
      n_0_2_44), .ZN(n_0_209));
   AOI22_X1 i_0_2_23 (.A1(n_0_2_168), .A2(n_0_2_43), .B1(n_0_2_125), .B2(
      n_0_2_44), .ZN(n_0_210));
   AOI22_X1 i_0_2_24 (.A1(n_0_2_169), .A2(n_0_2_43), .B1(n_0_2_126), .B2(
      n_0_2_44), .ZN(n_0_211));
   AOI22_X1 i_0_2_25 (.A1(n_0_2_170), .A2(n_0_2_43), .B1(n_0_2_127), .B2(
      n_0_2_44), .ZN(n_0_212));
   AOI22_X1 i_0_2_26 (.A1(n_0_2_171), .A2(n_0_2_43), .B1(n_0_2_128), .B2(
      n_0_2_44), .ZN(n_0_213));
   AOI22_X1 i_0_2_27 (.A1(n_0_2_172), .A2(n_0_2_43), .B1(n_0_2_129), .B2(
      n_0_2_44), .ZN(n_0_214));
   AOI22_X1 i_0_2_28 (.A1(n_0_2_173), .A2(n_0_2_43), .B1(n_0_2_130), .B2(
      n_0_2_44), .ZN(n_0_215));
   AOI22_X1 i_0_2_29 (.A1(n_0_2_174), .A2(n_0_2_43), .B1(n_0_2_131), .B2(
      n_0_2_44), .ZN(n_0_216));
   AOI22_X1 i_0_2_30 (.A1(n_0_2_175), .A2(n_0_2_43), .B1(n_0_2_132), .B2(
      n_0_2_44), .ZN(n_0_217));
   AOI22_X1 i_0_2_31 (.A1(n_0_2_176), .A2(n_0_2_43), .B1(n_0_2_133), .B2(
      n_0_2_44), .ZN(n_0_218));
   AOI22_X1 i_0_2_32 (.A1(n_0_2_177), .A2(n_0_2_43), .B1(n_0_2_134), .B2(
      n_0_2_44), .ZN(n_0_219));
   AOI22_X1 i_0_2_33 (.A1(n_0_2_178), .A2(n_0_2_43), .B1(n_0_2_135), .B2(
      n_0_2_44), .ZN(n_0_220));
   AOI22_X1 i_0_2_34 (.A1(n_0_2_179), .A2(n_0_2_43), .B1(n_0_2_136), .B2(
      n_0_2_44), .ZN(n_0_221));
   AOI22_X1 i_0_2_35 (.A1(n_0_2_180), .A2(n_0_2_43), .B1(n_0_2_137), .B2(
      n_0_2_44), .ZN(n_0_222));
   AOI22_X1 i_0_2_36 (.A1(n_0_2_181), .A2(n_0_2_43), .B1(n_0_2_138), .B2(
      n_0_2_44), .ZN(n_0_223));
   AOI22_X1 i_0_2_37 (.A1(n_0_2_182), .A2(n_0_2_43), .B1(n_0_2_139), .B2(
      n_0_2_44), .ZN(n_0_224));
   AOI22_X1 i_0_2_38 (.A1(n_0_2_183), .A2(n_0_2_43), .B1(n_0_2_140), .B2(
      n_0_2_44), .ZN(n_0_225));
   AOI22_X1 i_0_2_39 (.A1(n_0_2_184), .A2(n_0_2_43), .B1(n_0_2_141), .B2(
      n_0_2_44), .ZN(n_0_226));
   AOI22_X1 i_0_2_40 (.A1(n_0_2_185), .A2(n_0_2_43), .B1(n_0_2_142), .B2(
      n_0_2_44), .ZN(n_0_227));
   AOI22_X1 i_0_2_41 (.A1(n_0_2_186), .A2(n_0_2_43), .B1(n_0_2_143), .B2(
      n_0_2_44), .ZN(n_0_228));
   AOI22_X1 i_0_2_42 (.A1(n_0_2_187), .A2(n_0_2_43), .B1(n_0_2_145), .B2(
      n_0_2_44), .ZN(n_0_229));
   OAI21_X1 i_0_2_43 (.A(n_0_2_11), .B1(n_0_2_147), .B2(n_0_2_43), .ZN(n_0_230));
   NAND2_X1 i_0_2_44 (.A1(n_0_158), .A2(n_0_2_43), .ZN(n_0_2_11));
   OAI21_X1 i_0_2_45 (.A(n_0_2_12), .B1(n_0_2_47), .B2(n_0_2_43), .ZN(n_0_231));
   NAND2_X1 i_0_2_46 (.A1(n_0_159), .A2(n_0_2_43), .ZN(n_0_2_12));
   OAI21_X1 i_0_2_47 (.A(n_0_2_13), .B1(n_0_2_48), .B2(n_0_2_43), .ZN(n_0_232));
   NAND2_X1 i_0_2_48 (.A1(n_0_160), .A2(n_0_2_43), .ZN(n_0_2_13));
   OAI21_X1 i_0_2_49 (.A(n_0_2_14), .B1(n_0_2_49), .B2(n_0_2_43), .ZN(n_0_233));
   NAND2_X1 i_0_2_50 (.A1(n_0_161), .A2(n_0_2_43), .ZN(n_0_2_14));
   OAI21_X1 i_0_2_51 (.A(n_0_2_15), .B1(n_0_2_50), .B2(n_0_2_43), .ZN(n_0_234));
   NAND2_X1 i_0_2_52 (.A1(n_0_162), .A2(n_0_2_43), .ZN(n_0_2_15));
   OAI21_X1 i_0_2_53 (.A(n_0_2_16), .B1(n_0_2_51), .B2(n_0_2_43), .ZN(n_0_235));
   NAND2_X1 i_0_2_54 (.A1(n_0_163), .A2(n_0_2_43), .ZN(n_0_2_16));
   OAI21_X1 i_0_2_55 (.A(n_0_2_17), .B1(n_0_2_52), .B2(n_0_2_43), .ZN(n_0_236));
   NAND2_X1 i_0_2_56 (.A1(n_0_164), .A2(n_0_2_43), .ZN(n_0_2_17));
   OAI21_X1 i_0_2_57 (.A(n_0_2_18), .B1(n_0_2_53), .B2(n_0_2_43), .ZN(n_0_237));
   NAND2_X1 i_0_2_58 (.A1(n_0_165), .A2(n_0_2_43), .ZN(n_0_2_18));
   OAI21_X1 i_0_2_59 (.A(n_0_2_19), .B1(n_0_2_54), .B2(n_0_2_43), .ZN(n_0_238));
   NAND2_X1 i_0_2_60 (.A1(n_0_166), .A2(n_0_2_43), .ZN(n_0_2_19));
   OAI21_X1 i_0_2_61 (.A(n_0_2_20), .B1(n_0_2_55), .B2(n_0_2_43), .ZN(n_0_239));
   NAND2_X1 i_0_2_62 (.A1(n_0_167), .A2(n_0_2_43), .ZN(n_0_2_20));
   OAI21_X1 i_0_2_63 (.A(n_0_2_21), .B1(n_0_2_56), .B2(n_0_2_43), .ZN(n_0_240));
   NAND2_X1 i_0_2_64 (.A1(n_0_168), .A2(n_0_2_43), .ZN(n_0_2_21));
   OAI21_X1 i_0_2_65 (.A(n_0_2_22), .B1(n_0_2_57), .B2(n_0_2_43), .ZN(n_0_241));
   NAND2_X1 i_0_2_66 (.A1(n_0_169), .A2(n_0_2_43), .ZN(n_0_2_22));
   OAI21_X1 i_0_2_67 (.A(n_0_2_23), .B1(n_0_2_58), .B2(n_0_2_43), .ZN(n_0_242));
   NAND2_X1 i_0_2_68 (.A1(n_0_170), .A2(n_0_2_43), .ZN(n_0_2_23));
   OAI21_X1 i_0_2_69 (.A(n_0_2_24), .B1(n_0_2_59), .B2(n_0_2_43), .ZN(n_0_243));
   NAND2_X1 i_0_2_70 (.A1(n_0_171), .A2(n_0_2_43), .ZN(n_0_2_24));
   OAI21_X1 i_0_2_71 (.A(n_0_2_25), .B1(n_0_2_60), .B2(n_0_2_43), .ZN(n_0_244));
   NAND2_X1 i_0_2_72 (.A1(n_0_172), .A2(n_0_2_43), .ZN(n_0_2_25));
   OAI21_X1 i_0_2_73 (.A(n_0_2_26), .B1(n_0_2_61), .B2(n_0_2_43), .ZN(n_0_245));
   NAND2_X1 i_0_2_74 (.A1(n_0_173), .A2(n_0_2_43), .ZN(n_0_2_26));
   OAI21_X1 i_0_2_75 (.A(n_0_2_27), .B1(n_0_2_62), .B2(n_0_2_43), .ZN(n_0_246));
   NAND2_X1 i_0_2_76 (.A1(n_0_174), .A2(n_0_2_43), .ZN(n_0_2_27));
   OAI21_X1 i_0_2_77 (.A(n_0_2_28), .B1(n_0_2_63), .B2(n_0_2_43), .ZN(n_0_247));
   NAND2_X1 i_0_2_78 (.A1(n_0_175), .A2(n_0_2_43), .ZN(n_0_2_28));
   OAI21_X1 i_0_2_79 (.A(n_0_2_29), .B1(n_0_2_64), .B2(n_0_2_43), .ZN(n_0_248));
   NAND2_X1 i_0_2_80 (.A1(n_0_176), .A2(n_0_2_43), .ZN(n_0_2_29));
   OAI21_X1 i_0_2_81 (.A(n_0_2_30), .B1(n_0_2_65), .B2(n_0_2_43), .ZN(n_0_249));
   NAND2_X1 i_0_2_82 (.A1(n_0_177), .A2(n_0_2_43), .ZN(n_0_2_30));
   OAI21_X1 i_0_2_83 (.A(n_0_2_31), .B1(n_0_2_66), .B2(n_0_2_43), .ZN(n_0_250));
   NAND2_X1 i_0_2_84 (.A1(n_0_178), .A2(n_0_2_43), .ZN(n_0_2_31));
   OAI21_X1 i_0_2_85 (.A(n_0_2_32), .B1(n_0_2_67), .B2(n_0_2_43), .ZN(n_0_251));
   NAND2_X1 i_0_2_86 (.A1(n_0_179), .A2(n_0_2_43), .ZN(n_0_2_32));
   OAI21_X1 i_0_2_87 (.A(n_0_2_33), .B1(n_0_2_68), .B2(n_0_2_43), .ZN(n_0_252));
   NAND2_X1 i_0_2_88 (.A1(n_0_180), .A2(n_0_2_43), .ZN(n_0_2_33));
   OAI21_X1 i_0_2_89 (.A(n_0_2_34), .B1(n_0_2_69), .B2(n_0_2_43), .ZN(n_0_253));
   NAND2_X1 i_0_2_90 (.A1(n_0_181), .A2(n_0_2_43), .ZN(n_0_2_34));
   OAI21_X1 i_0_2_91 (.A(n_0_2_35), .B1(n_0_2_70), .B2(n_0_2_43), .ZN(n_0_254));
   NAND2_X1 i_0_2_92 (.A1(n_0_182), .A2(n_0_2_43), .ZN(n_0_2_35));
   OAI21_X1 i_0_2_93 (.A(n_0_2_36), .B1(n_0_2_71), .B2(n_0_2_43), .ZN(n_0_255));
   NAND2_X1 i_0_2_94 (.A1(n_0_183), .A2(n_0_2_43), .ZN(n_0_2_36));
   OAI21_X1 i_0_2_95 (.A(n_0_2_37), .B1(n_0_2_72), .B2(n_0_2_43), .ZN(n_0_256));
   NAND2_X1 i_0_2_96 (.A1(n_0_184), .A2(n_0_2_43), .ZN(n_0_2_37));
   OAI21_X1 i_0_2_97 (.A(n_0_2_38), .B1(n_0_2_73), .B2(n_0_2_43), .ZN(n_0_257));
   NAND2_X1 i_0_2_98 (.A1(n_0_185), .A2(n_0_2_43), .ZN(n_0_2_38));
   OAI21_X1 i_0_2_99 (.A(n_0_2_39), .B1(n_0_2_74), .B2(n_0_2_43), .ZN(n_0_258));
   NAND2_X1 i_0_2_100 (.A1(n_0_186), .A2(n_0_2_43), .ZN(n_0_2_39));
   OAI21_X1 i_0_2_101 (.A(n_0_2_40), .B1(n_0_2_75), .B2(n_0_2_43), .ZN(n_0_259));
   NAND2_X1 i_0_2_102 (.A1(n_0_187), .A2(n_0_2_43), .ZN(n_0_2_40));
   OAI21_X1 i_0_2_103 (.A(n_0_2_41), .B1(n_0_2_76), .B2(n_0_2_43), .ZN(n_0_260));
   NAND2_X1 i_0_2_104 (.A1(n_0_188), .A2(n_0_2_43), .ZN(n_0_2_41));
   OAI21_X1 i_0_2_105 (.A(n_0_2_42), .B1(n_0_2_77), .B2(n_0_2_43), .ZN(n_0_261));
   NAND2_X1 i_0_2_106 (.A1(n_0_189), .A2(n_0_2_43), .ZN(n_0_2_42));
   AND2_X1 i_0_2_107 (.A1(n_0_190), .A2(n_0_2_43), .ZN(n_0_262));
   INV_X1 i_0_2_108 (.A(n_0_2_44), .ZN(n_0_2_43));
   NOR4_X1 i_0_2_109 (.A1(n_0_192), .A2(n_0_2_45), .A3(n_0_2_46), .A4(out_sign), 
      .ZN(n_0_2_44));
   NAND2_X1 i_0_2_110 (.A1(SC[4]), .A2(SC[1]), .ZN(n_0_2_45));
   NAND3_X1 i_0_2_111 (.A1(SC[3]), .A2(SC[2]), .A3(n_0_2_154), .ZN(n_0_2_46));
   INV_X1 i_0_2_112 (.A(n_0_2_47), .ZN(n_0_263));
   AOI222_X1 i_0_2_113 (.A1(n_0_97), .A2(n_0_2_151), .B1(n_0_65), .B2(n_0_2_149), 
      .C1(A[1]), .C2(n_0_2_148), .ZN(n_0_2_47));
   INV_X1 i_0_2_114 (.A(n_0_2_48), .ZN(n_0_264));
   AOI222_X1 i_0_2_115 (.A1(n_0_98), .A2(n_0_2_151), .B1(n_0_66), .B2(n_0_2_149), 
      .C1(A[2]), .C2(n_0_2_148), .ZN(n_0_2_48));
   INV_X1 i_0_2_116 (.A(n_0_2_49), .ZN(n_0_265));
   AOI222_X1 i_0_2_117 (.A1(n_0_99), .A2(n_0_2_151), .B1(n_0_67), .B2(n_0_2_149), 
      .C1(A[3]), .C2(n_0_2_148), .ZN(n_0_2_49));
   INV_X1 i_0_2_118 (.A(n_0_2_50), .ZN(n_0_266));
   AOI222_X1 i_0_2_119 (.A1(n_0_100), .A2(n_0_2_151), .B1(n_0_68), .B2(n_0_2_149), 
      .C1(A[4]), .C2(n_0_2_148), .ZN(n_0_2_50));
   INV_X1 i_0_2_120 (.A(n_0_2_51), .ZN(n_0_267));
   AOI222_X1 i_0_2_121 (.A1(n_0_101), .A2(n_0_2_151), .B1(n_0_69), .B2(n_0_2_149), 
      .C1(A[5]), .C2(n_0_2_148), .ZN(n_0_2_51));
   INV_X1 i_0_2_122 (.A(n_0_2_52), .ZN(n_0_268));
   AOI222_X1 i_0_2_123 (.A1(n_0_102), .A2(n_0_2_151), .B1(n_0_70), .B2(n_0_2_149), 
      .C1(A[6]), .C2(n_0_2_148), .ZN(n_0_2_52));
   INV_X1 i_0_2_124 (.A(n_0_2_53), .ZN(n_0_269));
   AOI222_X1 i_0_2_125 (.A1(n_0_103), .A2(n_0_2_151), .B1(n_0_71), .B2(n_0_2_149), 
      .C1(A[7]), .C2(n_0_2_148), .ZN(n_0_2_53));
   INV_X1 i_0_2_126 (.A(n_0_2_54), .ZN(n_0_270));
   AOI222_X1 i_0_2_127 (.A1(n_0_104), .A2(n_0_2_151), .B1(n_0_72), .B2(n_0_2_149), 
      .C1(A[8]), .C2(n_0_2_148), .ZN(n_0_2_54));
   INV_X1 i_0_2_128 (.A(n_0_2_55), .ZN(n_0_271));
   AOI222_X1 i_0_2_129 (.A1(n_0_105), .A2(n_0_2_151), .B1(n_0_73), .B2(n_0_2_149), 
      .C1(A[9]), .C2(n_0_2_148), .ZN(n_0_2_55));
   INV_X1 i_0_2_130 (.A(n_0_2_56), .ZN(n_0_272));
   AOI222_X1 i_0_2_131 (.A1(n_0_106), .A2(n_0_2_151), .B1(n_0_74), .B2(n_0_2_149), 
      .C1(A[10]), .C2(n_0_2_148), .ZN(n_0_2_56));
   INV_X1 i_0_2_132 (.A(n_0_2_57), .ZN(n_0_273));
   AOI222_X1 i_0_2_133 (.A1(n_0_107), .A2(n_0_2_151), .B1(n_0_75), .B2(n_0_2_149), 
      .C1(A[11]), .C2(n_0_2_148), .ZN(n_0_2_57));
   INV_X1 i_0_2_134 (.A(n_0_2_58), .ZN(n_0_274));
   AOI222_X1 i_0_2_135 (.A1(n_0_108), .A2(n_0_2_151), .B1(n_0_76), .B2(n_0_2_149), 
      .C1(A[12]), .C2(n_0_2_148), .ZN(n_0_2_58));
   INV_X1 i_0_2_136 (.A(n_0_2_59), .ZN(n_0_275));
   AOI222_X1 i_0_2_137 (.A1(n_0_109), .A2(n_0_2_151), .B1(n_0_77), .B2(n_0_2_149), 
      .C1(A[13]), .C2(n_0_2_148), .ZN(n_0_2_59));
   INV_X1 i_0_2_138 (.A(n_0_2_60), .ZN(n_0_276));
   AOI222_X1 i_0_2_139 (.A1(n_0_110), .A2(n_0_2_151), .B1(n_0_78), .B2(n_0_2_149), 
      .C1(A[14]), .C2(n_0_2_148), .ZN(n_0_2_60));
   INV_X1 i_0_2_140 (.A(n_0_2_61), .ZN(n_0_277));
   AOI222_X1 i_0_2_141 (.A1(n_0_111), .A2(n_0_2_151), .B1(n_0_79), .B2(n_0_2_149), 
      .C1(A[15]), .C2(n_0_2_148), .ZN(n_0_2_61));
   INV_X1 i_0_2_142 (.A(n_0_2_62), .ZN(n_0_278));
   AOI222_X1 i_0_2_143 (.A1(n_0_112), .A2(n_0_2_151), .B1(n_0_80), .B2(n_0_2_149), 
      .C1(A[16]), .C2(n_0_2_148), .ZN(n_0_2_62));
   INV_X1 i_0_2_144 (.A(n_0_2_63), .ZN(n_0_279));
   AOI222_X1 i_0_2_145 (.A1(n_0_113), .A2(n_0_2_151), .B1(n_0_81), .B2(n_0_2_149), 
      .C1(A[17]), .C2(n_0_2_148), .ZN(n_0_2_63));
   INV_X1 i_0_2_146 (.A(n_0_2_64), .ZN(n_0_280));
   AOI222_X1 i_0_2_147 (.A1(n_0_114), .A2(n_0_2_151), .B1(n_0_82), .B2(n_0_2_149), 
      .C1(A[18]), .C2(n_0_2_148), .ZN(n_0_2_64));
   INV_X1 i_0_2_148 (.A(n_0_2_65), .ZN(n_0_281));
   AOI222_X1 i_0_2_149 (.A1(n_0_115), .A2(n_0_2_151), .B1(n_0_83), .B2(n_0_2_149), 
      .C1(A[19]), .C2(n_0_2_148), .ZN(n_0_2_65));
   INV_X1 i_0_2_150 (.A(n_0_2_66), .ZN(n_0_282));
   AOI222_X1 i_0_2_151 (.A1(n_0_116), .A2(n_0_2_151), .B1(n_0_84), .B2(n_0_2_149), 
      .C1(A[20]), .C2(n_0_2_148), .ZN(n_0_2_66));
   INV_X1 i_0_2_152 (.A(n_0_2_67), .ZN(n_0_283));
   AOI222_X1 i_0_2_153 (.A1(n_0_117), .A2(n_0_2_151), .B1(n_0_85), .B2(n_0_2_149), 
      .C1(A[21]), .C2(n_0_2_148), .ZN(n_0_2_67));
   INV_X1 i_0_2_154 (.A(n_0_2_68), .ZN(n_0_284));
   AOI222_X1 i_0_2_155 (.A1(n_0_118), .A2(n_0_2_151), .B1(n_0_86), .B2(n_0_2_149), 
      .C1(A[22]), .C2(n_0_2_148), .ZN(n_0_2_68));
   INV_X1 i_0_2_156 (.A(n_0_2_69), .ZN(n_0_285));
   AOI222_X1 i_0_2_157 (.A1(n_0_119), .A2(n_0_2_151), .B1(n_0_87), .B2(n_0_2_149), 
      .C1(A[23]), .C2(n_0_2_148), .ZN(n_0_2_69));
   INV_X1 i_0_2_158 (.A(n_0_2_70), .ZN(n_0_286));
   AOI222_X1 i_0_2_159 (.A1(n_0_120), .A2(n_0_2_151), .B1(n_0_88), .B2(n_0_2_149), 
      .C1(A[24]), .C2(n_0_2_148), .ZN(n_0_2_70));
   INV_X1 i_0_2_160 (.A(n_0_2_71), .ZN(n_0_287));
   AOI222_X1 i_0_2_161 (.A1(n_0_121), .A2(n_0_2_151), .B1(n_0_89), .B2(n_0_2_149), 
      .C1(A[25]), .C2(n_0_2_148), .ZN(n_0_2_71));
   INV_X1 i_0_2_162 (.A(n_0_2_72), .ZN(n_0_288));
   AOI222_X1 i_0_2_163 (.A1(n_0_122), .A2(n_0_2_151), .B1(n_0_90), .B2(n_0_2_149), 
      .C1(A[26]), .C2(n_0_2_148), .ZN(n_0_2_72));
   INV_X1 i_0_2_164 (.A(n_0_2_73), .ZN(n_0_289));
   AOI222_X1 i_0_2_165 (.A1(n_0_123), .A2(n_0_2_151), .B1(n_0_91), .B2(n_0_2_149), 
      .C1(A[27]), .C2(n_0_2_148), .ZN(n_0_2_73));
   INV_X1 i_0_2_166 (.A(n_0_2_74), .ZN(n_0_290));
   AOI222_X1 i_0_2_167 (.A1(n_0_124), .A2(n_0_2_151), .B1(n_0_92), .B2(n_0_2_149), 
      .C1(A[28]), .C2(n_0_2_148), .ZN(n_0_2_74));
   INV_X1 i_0_2_168 (.A(n_0_2_75), .ZN(n_0_291));
   AOI222_X1 i_0_2_169 (.A1(n_0_125), .A2(n_0_2_151), .B1(n_0_93), .B2(n_0_2_149), 
      .C1(A[29]), .C2(n_0_2_148), .ZN(n_0_2_75));
   INV_X1 i_0_2_170 (.A(n_0_2_76), .ZN(n_0_292));
   AOI222_X1 i_0_2_171 (.A1(n_0_126), .A2(n_0_2_151), .B1(n_0_94), .B2(n_0_2_149), 
      .C1(A[30]), .C2(n_0_2_148), .ZN(n_0_2_76));
   INV_X1 i_0_2_172 (.A(n_0_2_77), .ZN(n_0_293));
   AOI222_X1 i_0_2_173 (.A1(n_0_127), .A2(n_0_2_151), .B1(n_0_95), .B2(n_0_2_149), 
      .C1(A[31]), .C2(n_0_2_148), .ZN(n_0_2_77));
   INV_X1 i_0_2_174 (.A(n_0_2_78), .ZN(n_0_294));
   AOI22_X1 i_0_2_175 (.A1(multiplicand[0]), .A2(n_0_2_153), .B1(a[0]), .B2(
      n_0_2_152), .ZN(n_0_2_78));
   INV_X1 i_0_2_176 (.A(n_0_2_79), .ZN(n_0_295));
   AOI222_X1 i_0_2_177 (.A1(multiplicand[1]), .A2(n_0_2_153), .B1(n_0_33), 
      .B2(n_0_2_111), .C1(a[1]), .C2(n_0_2_110), .ZN(n_0_2_79));
   INV_X1 i_0_2_178 (.A(n_0_2_80), .ZN(n_0_296));
   AOI222_X1 i_0_2_179 (.A1(multiplicand[2]), .A2(n_0_2_153), .B1(n_0_34), 
      .B2(n_0_2_111), .C1(a[2]), .C2(n_0_2_110), .ZN(n_0_2_80));
   INV_X1 i_0_2_180 (.A(n_0_2_81), .ZN(n_0_297));
   AOI222_X1 i_0_2_181 (.A1(multiplicand[3]), .A2(n_0_2_153), .B1(n_0_35), 
      .B2(n_0_2_111), .C1(a[3]), .C2(n_0_2_110), .ZN(n_0_2_81));
   INV_X1 i_0_2_182 (.A(n_0_2_82), .ZN(n_0_298));
   AOI222_X1 i_0_2_183 (.A1(multiplicand[4]), .A2(n_0_2_153), .B1(n_0_36), 
      .B2(n_0_2_111), .C1(a[4]), .C2(n_0_2_110), .ZN(n_0_2_82));
   INV_X1 i_0_2_184 (.A(n_0_2_83), .ZN(n_0_299));
   AOI222_X1 i_0_2_185 (.A1(multiplicand[5]), .A2(n_0_2_153), .B1(n_0_37), 
      .B2(n_0_2_111), .C1(a[5]), .C2(n_0_2_110), .ZN(n_0_2_83));
   INV_X1 i_0_2_186 (.A(n_0_2_84), .ZN(n_0_300));
   AOI222_X1 i_0_2_187 (.A1(multiplicand[6]), .A2(n_0_2_153), .B1(n_0_38), 
      .B2(n_0_2_111), .C1(a[6]), .C2(n_0_2_110), .ZN(n_0_2_84));
   INV_X1 i_0_2_188 (.A(n_0_2_85), .ZN(n_0_301));
   AOI222_X1 i_0_2_189 (.A1(multiplicand[7]), .A2(n_0_2_153), .B1(n_0_39), 
      .B2(n_0_2_111), .C1(a[7]), .C2(n_0_2_110), .ZN(n_0_2_85));
   INV_X1 i_0_2_190 (.A(n_0_2_86), .ZN(n_0_302));
   AOI222_X1 i_0_2_191 (.A1(multiplicand[8]), .A2(n_0_2_153), .B1(n_0_40), 
      .B2(n_0_2_111), .C1(a[8]), .C2(n_0_2_110), .ZN(n_0_2_86));
   INV_X1 i_0_2_192 (.A(n_0_2_87), .ZN(n_0_303));
   AOI222_X1 i_0_2_193 (.A1(multiplicand[9]), .A2(n_0_2_153), .B1(n_0_41), 
      .B2(n_0_2_111), .C1(a[9]), .C2(n_0_2_110), .ZN(n_0_2_87));
   INV_X1 i_0_2_194 (.A(n_0_2_88), .ZN(n_0_304));
   AOI222_X1 i_0_2_195 (.A1(multiplicand[10]), .A2(n_0_2_153), .B1(n_0_42), 
      .B2(n_0_2_111), .C1(a[10]), .C2(n_0_2_110), .ZN(n_0_2_88));
   INV_X1 i_0_2_196 (.A(n_0_2_89), .ZN(n_0_305));
   AOI222_X1 i_0_2_197 (.A1(multiplicand[11]), .A2(n_0_2_153), .B1(n_0_43), 
      .B2(n_0_2_111), .C1(a[11]), .C2(n_0_2_110), .ZN(n_0_2_89));
   INV_X1 i_0_2_198 (.A(n_0_2_90), .ZN(n_0_306));
   AOI222_X1 i_0_2_199 (.A1(multiplicand[12]), .A2(n_0_2_153), .B1(n_0_44), 
      .B2(n_0_2_111), .C1(a[12]), .C2(n_0_2_110), .ZN(n_0_2_90));
   INV_X1 i_0_2_200 (.A(n_0_2_91), .ZN(n_0_307));
   AOI222_X1 i_0_2_201 (.A1(multiplicand[13]), .A2(n_0_2_153), .B1(n_0_45), 
      .B2(n_0_2_111), .C1(a[13]), .C2(n_0_2_110), .ZN(n_0_2_91));
   INV_X1 i_0_2_202 (.A(n_0_2_92), .ZN(n_0_308));
   AOI222_X1 i_0_2_203 (.A1(multiplicand[14]), .A2(n_0_2_153), .B1(n_0_46), 
      .B2(n_0_2_111), .C1(a[14]), .C2(n_0_2_110), .ZN(n_0_2_92));
   INV_X1 i_0_2_204 (.A(n_0_2_93), .ZN(n_0_309));
   AOI222_X1 i_0_2_205 (.A1(multiplicand[15]), .A2(n_0_2_153), .B1(n_0_47), 
      .B2(n_0_2_111), .C1(a[15]), .C2(n_0_2_110), .ZN(n_0_2_93));
   INV_X1 i_0_2_206 (.A(n_0_2_94), .ZN(n_0_310));
   AOI222_X1 i_0_2_207 (.A1(multiplicand[16]), .A2(n_0_2_153), .B1(n_0_48), 
      .B2(n_0_2_111), .C1(a[16]), .C2(n_0_2_110), .ZN(n_0_2_94));
   INV_X1 i_0_2_208 (.A(n_0_2_95), .ZN(n_0_311));
   AOI222_X1 i_0_2_209 (.A1(multiplicand[17]), .A2(n_0_2_153), .B1(n_0_49), 
      .B2(n_0_2_111), .C1(a[17]), .C2(n_0_2_110), .ZN(n_0_2_95));
   INV_X1 i_0_2_210 (.A(n_0_2_96), .ZN(n_0_312));
   AOI222_X1 i_0_2_211 (.A1(multiplicand[18]), .A2(n_0_2_153), .B1(n_0_50), 
      .B2(n_0_2_111), .C1(a[18]), .C2(n_0_2_110), .ZN(n_0_2_96));
   INV_X1 i_0_2_212 (.A(n_0_2_97), .ZN(n_0_313));
   AOI222_X1 i_0_2_213 (.A1(multiplicand[19]), .A2(n_0_2_153), .B1(n_0_51), 
      .B2(n_0_2_111), .C1(a[19]), .C2(n_0_2_110), .ZN(n_0_2_97));
   INV_X1 i_0_2_214 (.A(n_0_2_98), .ZN(n_0_314));
   AOI222_X1 i_0_2_215 (.A1(multiplicand[20]), .A2(n_0_2_153), .B1(n_0_52), 
      .B2(n_0_2_111), .C1(a[20]), .C2(n_0_2_110), .ZN(n_0_2_98));
   INV_X1 i_0_2_216 (.A(n_0_2_99), .ZN(n_0_315));
   AOI222_X1 i_0_2_217 (.A1(multiplicand[21]), .A2(n_0_2_153), .B1(n_0_53), 
      .B2(n_0_2_111), .C1(a[21]), .C2(n_0_2_110), .ZN(n_0_2_99));
   INV_X1 i_0_2_218 (.A(n_0_2_100), .ZN(n_0_316));
   AOI222_X1 i_0_2_219 (.A1(multiplicand[22]), .A2(n_0_2_153), .B1(n_0_54), 
      .B2(n_0_2_111), .C1(a[22]), .C2(n_0_2_110), .ZN(n_0_2_100));
   INV_X1 i_0_2_220 (.A(n_0_2_101), .ZN(n_0_317));
   AOI222_X1 i_0_2_221 (.A1(multiplicand[23]), .A2(n_0_2_153), .B1(n_0_55), 
      .B2(n_0_2_111), .C1(a[23]), .C2(n_0_2_110), .ZN(n_0_2_101));
   INV_X1 i_0_2_222 (.A(n_0_2_102), .ZN(n_0_318));
   AOI222_X1 i_0_2_223 (.A1(multiplicand[24]), .A2(n_0_2_153), .B1(n_0_56), 
      .B2(n_0_2_111), .C1(a[24]), .C2(n_0_2_110), .ZN(n_0_2_102));
   INV_X1 i_0_2_224 (.A(n_0_2_103), .ZN(n_0_319));
   AOI222_X1 i_0_2_225 (.A1(multiplicand[25]), .A2(n_0_2_153), .B1(n_0_57), 
      .B2(n_0_2_111), .C1(a[25]), .C2(n_0_2_110), .ZN(n_0_2_103));
   INV_X1 i_0_2_226 (.A(n_0_2_104), .ZN(n_0_320));
   AOI222_X1 i_0_2_227 (.A1(multiplicand[26]), .A2(n_0_2_153), .B1(n_0_58), 
      .B2(n_0_2_111), .C1(a[26]), .C2(n_0_2_110), .ZN(n_0_2_104));
   INV_X1 i_0_2_228 (.A(n_0_2_105), .ZN(n_0_321));
   AOI222_X1 i_0_2_229 (.A1(multiplicand[27]), .A2(n_0_2_153), .B1(n_0_59), 
      .B2(n_0_2_111), .C1(a[27]), .C2(n_0_2_110), .ZN(n_0_2_105));
   INV_X1 i_0_2_230 (.A(n_0_2_106), .ZN(n_0_322));
   AOI222_X1 i_0_2_231 (.A1(multiplicand[28]), .A2(n_0_2_153), .B1(n_0_60), 
      .B2(n_0_2_111), .C1(a[28]), .C2(n_0_2_110), .ZN(n_0_2_106));
   INV_X1 i_0_2_232 (.A(n_0_2_107), .ZN(n_0_323));
   AOI222_X1 i_0_2_233 (.A1(multiplicand[29]), .A2(n_0_2_153), .B1(n_0_61), 
      .B2(n_0_2_111), .C1(a[29]), .C2(n_0_2_110), .ZN(n_0_2_107));
   INV_X1 i_0_2_234 (.A(n_0_2_108), .ZN(n_0_324));
   AOI222_X1 i_0_2_235 (.A1(multiplicand[30]), .A2(n_0_2_153), .B1(n_0_62), 
      .B2(n_0_2_111), .C1(a[30]), .C2(n_0_2_110), .ZN(n_0_2_108));
   INV_X1 i_0_2_236 (.A(n_0_2_109), .ZN(n_0_325));
   AOI22_X1 i_0_2_237 (.A1(multiplicand[31]), .A2(n_0_2_153), .B1(n_0_63), 
      .B2(n_0_2_111), .ZN(n_0_2_109));
   NOR2_X1 i_0_2_238 (.A1(a[31]), .A2(n_0_2_153), .ZN(n_0_2_110));
   NOR2_X1 i_0_2_239 (.A1(n_0_2_188), .A2(n_0_2_153), .ZN(n_0_2_111));
   INV_X1 i_0_2_240 (.A(n_0_2_112), .ZN(n_0_326));
   NAND4_X1 i_0_2_241 (.A1(SC[4]), .A2(SC[3]), .A3(n_0_2_154), .A4(n_0_2_113), 
      .ZN(n_0_2_112));
   AND3_X1 i_0_2_242 (.A1(SC[2]), .A2(SC[1]), .A3(SC[0]), .ZN(n_0_2_113));
   INV_X1 i_0_2_243 (.A(n_0_2_114), .ZN(n_0_328));
   AOI222_X1 i_0_2_244 (.A1(Q[2]), .A2(n_0_2_153), .B1(b[1]), .B2(n_0_2_144), 
      .C1(n_0_2), .C2(n_0_2_146), .ZN(n_0_2_114));
   INV_X1 i_0_2_245 (.A(n_0_2_115), .ZN(n_0_329));
   AOI222_X1 i_0_2_246 (.A1(Q[3]), .A2(n_0_2_153), .B1(b[2]), .B2(n_0_2_144), 
      .C1(n_0_3), .C2(n_0_2_146), .ZN(n_0_2_115));
   INV_X1 i_0_2_247 (.A(n_0_2_116), .ZN(n_0_330));
   AOI222_X1 i_0_2_248 (.A1(Q[4]), .A2(n_0_2_153), .B1(b[3]), .B2(n_0_2_144), 
      .C1(n_0_4), .C2(n_0_2_146), .ZN(n_0_2_116));
   INV_X1 i_0_2_249 (.A(n_0_2_117), .ZN(n_0_331));
   AOI222_X1 i_0_2_250 (.A1(Q[5]), .A2(n_0_2_153), .B1(b[4]), .B2(n_0_2_144), 
      .C1(n_0_5), .C2(n_0_2_146), .ZN(n_0_2_117));
   INV_X1 i_0_2_251 (.A(n_0_2_118), .ZN(n_0_332));
   AOI222_X1 i_0_2_252 (.A1(Q[6]), .A2(n_0_2_153), .B1(b[5]), .B2(n_0_2_144), 
      .C1(n_0_6), .C2(n_0_2_146), .ZN(n_0_2_118));
   INV_X1 i_0_2_253 (.A(n_0_2_119), .ZN(n_0_333));
   AOI222_X1 i_0_2_254 (.A1(Q[7]), .A2(n_0_2_153), .B1(b[6]), .B2(n_0_2_144), 
      .C1(n_0_7), .C2(n_0_2_146), .ZN(n_0_2_119));
   INV_X1 i_0_2_255 (.A(n_0_2_120), .ZN(n_0_334));
   AOI222_X1 i_0_2_256 (.A1(Q[8]), .A2(n_0_2_153), .B1(b[7]), .B2(n_0_2_144), 
      .C1(n_0_8), .C2(n_0_2_146), .ZN(n_0_2_120));
   INV_X1 i_0_2_257 (.A(n_0_2_121), .ZN(n_0_335));
   AOI222_X1 i_0_2_258 (.A1(Q[9]), .A2(n_0_2_153), .B1(b[8]), .B2(n_0_2_144), 
      .C1(n_0_9), .C2(n_0_2_146), .ZN(n_0_2_121));
   INV_X1 i_0_2_259 (.A(n_0_2_122), .ZN(n_0_336));
   AOI222_X1 i_0_2_260 (.A1(Q[10]), .A2(n_0_2_153), .B1(b[9]), .B2(n_0_2_144), 
      .C1(n_0_10), .C2(n_0_2_146), .ZN(n_0_2_122));
   INV_X1 i_0_2_261 (.A(n_0_2_123), .ZN(n_0_337));
   AOI222_X1 i_0_2_262 (.A1(Q[11]), .A2(n_0_2_153), .B1(b[10]), .B2(n_0_2_144), 
      .C1(n_0_11), .C2(n_0_2_146), .ZN(n_0_2_123));
   INV_X1 i_0_2_263 (.A(n_0_2_124), .ZN(n_0_338));
   AOI222_X1 i_0_2_264 (.A1(Q[12]), .A2(n_0_2_153), .B1(b[11]), .B2(n_0_2_144), 
      .C1(n_0_12), .C2(n_0_2_146), .ZN(n_0_2_124));
   INV_X1 i_0_2_265 (.A(n_0_2_125), .ZN(n_0_339));
   AOI222_X1 i_0_2_266 (.A1(Q[13]), .A2(n_0_2_153), .B1(b[12]), .B2(n_0_2_144), 
      .C1(n_0_13), .C2(n_0_2_146), .ZN(n_0_2_125));
   INV_X1 i_0_2_267 (.A(n_0_2_126), .ZN(n_0_340));
   AOI222_X1 i_0_2_268 (.A1(Q[14]), .A2(n_0_2_153), .B1(b[13]), .B2(n_0_2_144), 
      .C1(n_0_14), .C2(n_0_2_146), .ZN(n_0_2_126));
   INV_X1 i_0_2_269 (.A(n_0_2_127), .ZN(n_0_341));
   AOI222_X1 i_0_2_270 (.A1(Q[15]), .A2(n_0_2_153), .B1(b[14]), .B2(n_0_2_144), 
      .C1(n_0_15), .C2(n_0_2_146), .ZN(n_0_2_127));
   INV_X1 i_0_2_271 (.A(n_0_2_128), .ZN(n_0_342));
   AOI222_X1 i_0_2_272 (.A1(Q[16]), .A2(n_0_2_153), .B1(b[15]), .B2(n_0_2_144), 
      .C1(n_0_16), .C2(n_0_2_146), .ZN(n_0_2_128));
   INV_X1 i_0_2_273 (.A(n_0_2_129), .ZN(n_0_343));
   AOI222_X1 i_0_2_274 (.A1(Q[17]), .A2(n_0_2_153), .B1(b[16]), .B2(n_0_2_144), 
      .C1(n_0_17), .C2(n_0_2_146), .ZN(n_0_2_129));
   INV_X1 i_0_2_275 (.A(n_0_2_130), .ZN(n_0_344));
   AOI222_X1 i_0_2_276 (.A1(Q[18]), .A2(n_0_2_153), .B1(b[17]), .B2(n_0_2_144), 
      .C1(n_0_18), .C2(n_0_2_146), .ZN(n_0_2_130));
   INV_X1 i_0_2_277 (.A(n_0_2_131), .ZN(n_0_345));
   AOI222_X1 i_0_2_278 (.A1(Q[19]), .A2(n_0_2_153), .B1(b[18]), .B2(n_0_2_144), 
      .C1(n_0_19), .C2(n_0_2_146), .ZN(n_0_2_131));
   INV_X1 i_0_2_279 (.A(n_0_2_132), .ZN(n_0_346));
   AOI222_X1 i_0_2_280 (.A1(Q[20]), .A2(n_0_2_153), .B1(b[19]), .B2(n_0_2_144), 
      .C1(n_0_20), .C2(n_0_2_146), .ZN(n_0_2_132));
   INV_X1 i_0_2_281 (.A(n_0_2_133), .ZN(n_0_347));
   AOI222_X1 i_0_2_282 (.A1(Q[21]), .A2(n_0_2_153), .B1(b[20]), .B2(n_0_2_144), 
      .C1(n_0_21), .C2(n_0_2_146), .ZN(n_0_2_133));
   INV_X1 i_0_2_283 (.A(n_0_2_134), .ZN(n_0_348));
   AOI222_X1 i_0_2_284 (.A1(Q[22]), .A2(n_0_2_153), .B1(b[21]), .B2(n_0_2_144), 
      .C1(n_0_22), .C2(n_0_2_146), .ZN(n_0_2_134));
   INV_X1 i_0_2_285 (.A(n_0_2_135), .ZN(n_0_349));
   AOI222_X1 i_0_2_286 (.A1(Q[23]), .A2(n_0_2_153), .B1(b[22]), .B2(n_0_2_144), 
      .C1(n_0_23), .C2(n_0_2_146), .ZN(n_0_2_135));
   INV_X1 i_0_2_287 (.A(n_0_2_136), .ZN(n_0_350));
   AOI222_X1 i_0_2_288 (.A1(Q[24]), .A2(n_0_2_153), .B1(b[23]), .B2(n_0_2_144), 
      .C1(n_0_24), .C2(n_0_2_146), .ZN(n_0_2_136));
   INV_X1 i_0_2_289 (.A(n_0_2_137), .ZN(n_0_351));
   AOI222_X1 i_0_2_290 (.A1(Q[25]), .A2(n_0_2_153), .B1(b[24]), .B2(n_0_2_144), 
      .C1(n_0_25), .C2(n_0_2_146), .ZN(n_0_2_137));
   INV_X1 i_0_2_291 (.A(n_0_2_138), .ZN(n_0_352));
   AOI222_X1 i_0_2_292 (.A1(Q[26]), .A2(n_0_2_153), .B1(b[25]), .B2(n_0_2_144), 
      .C1(n_0_26), .C2(n_0_2_146), .ZN(n_0_2_138));
   INV_X1 i_0_2_293 (.A(n_0_2_139), .ZN(n_0_353));
   AOI222_X1 i_0_2_294 (.A1(Q[27]), .A2(n_0_2_153), .B1(b[26]), .B2(n_0_2_144), 
      .C1(n_0_27), .C2(n_0_2_146), .ZN(n_0_2_139));
   INV_X1 i_0_2_295 (.A(n_0_2_140), .ZN(n_0_354));
   AOI222_X1 i_0_2_296 (.A1(Q[28]), .A2(n_0_2_153), .B1(b[27]), .B2(n_0_2_144), 
      .C1(n_0_28), .C2(n_0_2_146), .ZN(n_0_2_140));
   INV_X1 i_0_2_297 (.A(n_0_2_141), .ZN(n_0_355));
   AOI222_X1 i_0_2_298 (.A1(Q[29]), .A2(n_0_2_153), .B1(b[28]), .B2(n_0_2_144), 
      .C1(n_0_29), .C2(n_0_2_146), .ZN(n_0_2_141));
   INV_X1 i_0_2_299 (.A(n_0_2_142), .ZN(n_0_356));
   AOI222_X1 i_0_2_300 (.A1(Q[30]), .A2(n_0_2_153), .B1(b[29]), .B2(n_0_2_144), 
      .C1(n_0_30), .C2(n_0_2_146), .ZN(n_0_2_142));
   INV_X1 i_0_2_301 (.A(n_0_2_143), .ZN(n_0_357));
   AOI222_X1 i_0_2_302 (.A1(Q[31]), .A2(n_0_2_153), .B1(b[30]), .B2(n_0_2_144), 
      .C1(n_0_31), .C2(n_0_2_146), .ZN(n_0_2_143));
   NOR2_X1 i_0_2_303 (.A1(b[31]), .A2(n_0_2_153), .ZN(n_0_2_144));
   INV_X1 i_0_2_304 (.A(n_0_2_145), .ZN(n_0_358));
   AOI22_X1 i_0_2_305 (.A1(n_0_32), .A2(n_0_2_146), .B1(Q[32]), .B2(n_0_2_153), 
      .ZN(n_0_2_145));
   AND2_X1 i_0_2_306 (.A1(b[31]), .A2(n_0_2_152), .ZN(n_0_2_146));
   INV_X1 i_0_2_307 (.A(n_0_2_147), .ZN(n_0_359));
   AOI222_X1 i_0_2_308 (.A1(n_0_96), .A2(n_0_2_151), .B1(n_0_64), .B2(n_0_2_149), 
      .C1(A[0]), .C2(n_0_2_148), .ZN(n_0_2_147));
   NOR2_X1 i_0_2_309 (.A1(n_0_2_151), .A2(n_0_2_149), .ZN(n_0_2_148));
   AOI21_X1 i_0_2_310 (.A(n_0_2_150), .B1(Q[0]), .B2(n_0_2_153), .ZN(n_0_2_149));
   INV_X1 i_0_2_311 (.A(n_0_2_150), .ZN(n_0_327));
   AOI22_X1 i_0_2_312 (.A1(Q[1]), .A2(n_0_2_153), .B1(b[0]), .B2(n_0_2_152), 
      .ZN(n_0_2_150));
   NOR3_X1 i_0_2_313 (.A1(Q[1]), .A2(n_0_2_152), .A3(n_0_2_189), .ZN(n_0_2_151));
   INV_X1 i_0_2_314 (.A(n_0_2_153), .ZN(n_0_2_152));
   NAND3_X1 i_0_2_315 (.A1(n_0_2_155), .A2(n_0_2_154), .A3(n_0_2_156), .ZN(
      n_0_2_153));
   NOR2_X1 i_0_2_316 (.A1(SC[6]), .A2(SC[5]), .ZN(n_0_2_154));
   NOR2_X1 i_0_2_317 (.A1(SC[4]), .A2(SC[3]), .ZN(n_0_2_155));
   NOR3_X1 i_0_2_318 (.A1(SC[2]), .A2(SC[1]), .A3(SC[0]), .ZN(n_0_2_156));
   INV_X1 i_0_2_319 (.A(n_0_2_4), .ZN(n_0_2_157));
   INV_X1 i_0_2_320 (.A(n_0_128), .ZN(n_0_2_158));
   INV_X1 i_0_2_321 (.A(n_0_129), .ZN(n_0_2_159));
   INV_X1 i_0_2_322 (.A(n_0_130), .ZN(n_0_2_160));
   INV_X1 i_0_2_323 (.A(n_0_131), .ZN(n_0_2_161));
   INV_X1 i_0_2_324 (.A(n_0_132), .ZN(n_0_2_162));
   INV_X1 i_0_2_325 (.A(n_0_133), .ZN(n_0_2_163));
   INV_X1 i_0_2_326 (.A(n_0_134), .ZN(n_0_2_164));
   INV_X1 i_0_2_327 (.A(n_0_135), .ZN(n_0_2_165));
   INV_X1 i_0_2_328 (.A(n_0_136), .ZN(n_0_2_166));
   INV_X1 i_0_2_329 (.A(n_0_137), .ZN(n_0_2_167));
   INV_X1 i_0_2_330 (.A(n_0_138), .ZN(n_0_2_168));
   INV_X1 i_0_2_331 (.A(n_0_139), .ZN(n_0_2_169));
   INV_X1 i_0_2_332 (.A(n_0_140), .ZN(n_0_2_170));
   INV_X1 i_0_2_333 (.A(n_0_141), .ZN(n_0_2_171));
   INV_X1 i_0_2_334 (.A(n_0_142), .ZN(n_0_2_172));
   INV_X1 i_0_2_335 (.A(n_0_143), .ZN(n_0_2_173));
   INV_X1 i_0_2_336 (.A(n_0_144), .ZN(n_0_2_174));
   INV_X1 i_0_2_337 (.A(n_0_145), .ZN(n_0_2_175));
   INV_X1 i_0_2_338 (.A(n_0_146), .ZN(n_0_2_176));
   INV_X1 i_0_2_339 (.A(n_0_147), .ZN(n_0_2_177));
   INV_X1 i_0_2_340 (.A(n_0_148), .ZN(n_0_2_178));
   INV_X1 i_0_2_341 (.A(n_0_149), .ZN(n_0_2_179));
   INV_X1 i_0_2_342 (.A(n_0_150), .ZN(n_0_2_180));
   INV_X1 i_0_2_343 (.A(n_0_151), .ZN(n_0_2_181));
   INV_X1 i_0_2_344 (.A(n_0_152), .ZN(n_0_2_182));
   INV_X1 i_0_2_345 (.A(n_0_153), .ZN(n_0_2_183));
   INV_X1 i_0_2_346 (.A(n_0_154), .ZN(n_0_2_184));
   INV_X1 i_0_2_347 (.A(n_0_155), .ZN(n_0_2_185));
   INV_X1 i_0_2_348 (.A(n_0_156), .ZN(n_0_2_186));
   INV_X1 i_0_2_349 (.A(n_0_157), .ZN(n_0_2_187));
   INV_X1 i_0_2_350 (.A(a[31]), .ZN(n_0_2_188));
   INV_X1 i_0_2_351 (.A(Q[0]), .ZN(n_0_2_189));
   INV_X1 i_0_2_352 (.A(SC[0]), .ZN(n_0_192));
   INV_X1 i_0_2_353 (.A(SC[6]), .ZN(n_0_2_190));
endmodule
