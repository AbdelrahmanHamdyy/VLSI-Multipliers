/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu Dec 22 18:59:11 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 380499138 */

module datapath(firstInputComplement, inputOne);
   output [31:0]firstInputComplement;
   input [31:0]inputOne;

   AOI21_X1 i_0 (.A(n_3), .B1(inputOne[1]), .B2(inputOne[0]), .ZN(
      firstInputComplement[1]));
   AOI21_X1 i_1 (.A(n_12), .B1(inputOne[4]), .B2(n_5), .ZN(
      firstInputComplement[4]));
   AOI21_X1 i_2 (.A(n_10), .B1(inputOne[5]), .B2(n_11), .ZN(
      firstInputComplement[5]));
   AOI21_X1 i_3 (.A(n_22), .B1(inputOne[7]), .B2(n_0), .ZN(
      firstInputComplement[7]));
   INV_X1 i_4 (.A(n_8), .ZN(n_0));
   AOI21_X1 i_5 (.A(n_20), .B1(inputOne[8]), .B2(n_21), .ZN(
      firstInputComplement[8]));
   AOI21_X1 i_6 (.A(n_18), .B1(inputOne[9]), .B2(n_19), .ZN(
      firstInputComplement[9]));
   AOI21_X1 i_23 (.A(n_38), .B1(inputOne[12]), .B2(n_30), .ZN(
      firstInputComplement[12]));
   AOI21_X1 i_24 (.A(n_36), .B1(inputOne[13]), .B2(n_37), .ZN(
      firstInputComplement[13]));
   AOI21_X1 i_33 (.A(n_51), .B1(inputOne[16]), .B2(n_44), .ZN(
      firstInputComplement[16]));
   AOI21_X1 i_34 (.A(n_49), .B1(inputOne[17]), .B2(n_50), .ZN(
      firstInputComplement[17]));
   AOI21_X1 i_43 (.A(n_61), .B1(inputOne[20]), .B2(n_56), .ZN(
      firstInputComplement[20]));
   AOI21_X1 i_7 (.A(n_77), .B1(inputOne[23]), .B2(n_63), .ZN(
      firstInputComplement[23]));
   AOI21_X1 i_8 (.A(n_68), .B1(inputOne[24]), .B2(n_69), .ZN(
      firstInputComplement[24]));
   AOI22_X1 i_9 (.A1(n_80), .A2(inputOne[29]), .B1(n_74), .B2(n_83), .ZN(
      firstInputComplement[29]));
   INV_X1 i_10 (.A(n_1), .ZN(firstInputComplement[2]));
   OAI21_X1 i_11 (.A(n_2), .B1(n_4), .B2(n_3), .ZN(n_1));
   NAND2_X1 i_12 (.A1(n_4), .A2(n_3), .ZN(n_2));
   NOR2_X1 i_13 (.A1(inputOne[1]), .A2(inputOne[0]), .ZN(n_3));
   INV_X1 i_14 (.A(inputOne[2]), .ZN(n_4));
   AOI21_X1 i_15 (.A(n_6), .B1(inputOne[3]), .B2(n_2), .ZN(
      firstInputComplement[3]));
   INV_X1 i_16 (.A(n_6), .ZN(n_5));
   NOR4_X1 i_17 (.A1(inputOne[3]), .A2(inputOne[0]), .A3(n_7), .A4(inputOne[1]), 
      .ZN(n_6));
   INV_X1 i_18 (.A(n_4), .ZN(n_7));
   AOI21_X1 i_19 (.A(n_8), .B1(inputOne[6]), .B2(n_9), .ZN(
      firstInputComplement[6]));
   NOR2_X1 i_20 (.A1(inputOne[6]), .A2(n_9), .ZN(n_8));
   INV_X1 i_21 (.A(n_10), .ZN(n_9));
   NOR2_X1 i_22 (.A1(inputOne[5]), .A2(n_11), .ZN(n_10));
   INV_X1 i_25 (.A(n_12), .ZN(n_11));
   NOR2_X1 i_26 (.A1(inputOne[4]), .A2(n_5), .ZN(n_12));
   INV_X1 i_27 (.A(inputOne[4]), .ZN(n_13));
   INV_X1 i_28 (.A(inputOne[5]), .ZN(n_14));
   INV_X1 i_29 (.A(inputOne[6]), .ZN(n_15));
   AOI21_X1 i_30 (.A(n_16), .B1(inputOne[10]), .B2(n_17), .ZN(
      firstInputComplement[10]));
   NOR2_X1 i_31 (.A1(inputOne[10]), .A2(n_17), .ZN(n_16));
   INV_X1 i_32 (.A(n_18), .ZN(n_17));
   NOR2_X1 i_35 (.A1(inputOne[9]), .A2(n_19), .ZN(n_18));
   INV_X1 i_36 (.A(n_20), .ZN(n_19));
   NOR2_X1 i_37 (.A1(inputOne[8]), .A2(n_21), .ZN(n_20));
   INV_X1 i_38 (.A(n_22), .ZN(n_21));
   NOR2_X1 i_39 (.A1(n_5), .A2(n_23), .ZN(n_22));
   NAND4_X1 i_40 (.A1(n_14), .A2(n_13), .A3(n_24), .A4(n_15), .ZN(n_23));
   INV_X1 i_41 (.A(inputOne[7]), .ZN(n_24));
   INV_X1 i_42 (.A(inputOne[8]), .ZN(n_25));
   INV_X1 i_44 (.A(inputOne[9]), .ZN(n_26));
   INV_X1 i_45 (.A(inputOne[10]), .ZN(n_27));
   INV_X1 i_46 (.A(n_28), .ZN(firstInputComplement[11]));
   OAI21_X1 i_47 (.A(n_30), .B1(n_32), .B2(n_16), .ZN(n_28));
   INV_X1 i_48 (.A(n_30), .ZN(n_29));
   NAND3_X1 i_49 (.A1(n_33), .A2(n_6), .A3(n_31), .ZN(n_30));
   AND4_X1 i_50 (.A1(n_26), .A2(n_25), .A3(n_32), .A4(n_27), .ZN(n_31));
   INV_X1 i_51 (.A(inputOne[11]), .ZN(n_32));
   INV_X1 i_52 (.A(n_23), .ZN(n_33));
   AOI21_X1 i_53 (.A(n_34), .B1(inputOne[14]), .B2(n_35), .ZN(
      firstInputComplement[14]));
   NOR2_X1 i_54 (.A1(inputOne[14]), .A2(n_35), .ZN(n_34));
   INV_X1 i_55 (.A(n_36), .ZN(n_35));
   NOR2_X1 i_56 (.A1(inputOne[13]), .A2(n_37), .ZN(n_36));
   INV_X1 i_57 (.A(n_38), .ZN(n_37));
   NOR2_X1 i_58 (.A1(inputOne[12]), .A2(n_30), .ZN(n_38));
   INV_X1 i_59 (.A(inputOne[12]), .ZN(n_39));
   INV_X1 i_60 (.A(inputOne[13]), .ZN(n_40));
   INV_X1 i_61 (.A(inputOne[14]), .ZN(n_41));
   INV_X1 i_62 (.A(n_42), .ZN(firstInputComplement[15]));
   OAI21_X1 i_63 (.A(n_44), .B1(n_46), .B2(n_34), .ZN(n_42));
   INV_X1 i_64 (.A(n_44), .ZN(n_43));
   NAND4_X1 i_65 (.A1(n_6), .A2(n_31), .A3(n_45), .A4(n_33), .ZN(n_44));
   AND4_X1 i_66 (.A1(n_40), .A2(n_39), .A3(n_46), .A4(n_41), .ZN(n_45));
   INV_X1 i_67 (.A(inputOne[15]), .ZN(n_46));
   AOI21_X1 i_68 (.A(n_47), .B1(inputOne[18]), .B2(n_48), .ZN(
      firstInputComplement[18]));
   NOR2_X1 i_69 (.A1(inputOne[18]), .A2(n_48), .ZN(n_47));
   INV_X1 i_70 (.A(n_49), .ZN(n_48));
   NOR2_X1 i_71 (.A1(inputOne[17]), .A2(n_50), .ZN(n_49));
   INV_X1 i_72 (.A(n_51), .ZN(n_50));
   NOR2_X1 i_73 (.A1(inputOne[16]), .A2(n_44), .ZN(n_51));
   INV_X1 i_74 (.A(inputOne[16]), .ZN(n_52));
   INV_X1 i_75 (.A(inputOne[17]), .ZN(n_53));
   INV_X1 i_76 (.A(inputOne[18]), .ZN(n_54));
   INV_X1 i_77 (.A(n_55), .ZN(firstInputComplement[19]));
   OAI21_X1 i_78 (.A(n_56), .B1(n_58), .B2(n_47), .ZN(n_55));
   NAND2_X1 i_79 (.A1(n_43), .A2(n_57), .ZN(n_56));
   AND4_X1 i_80 (.A1(n_53), .A2(n_52), .A3(n_58), .A4(n_54), .ZN(n_57));
   INV_X1 i_81 (.A(inputOne[19]), .ZN(n_58));
   AOI21_X1 i_82 (.A(n_59), .B1(inputOne[21]), .B2(n_60), .ZN(
      firstInputComplement[21]));
   NOR2_X1 i_83 (.A1(inputOne[21]), .A2(n_60), .ZN(n_59));
   INV_X1 i_84 (.A(n_61), .ZN(n_60));
   NOR2_X1 i_85 (.A1(inputOne[20]), .A2(n_56), .ZN(n_61));
   AOI21_X1 i_86 (.A(n_62), .B1(inputOne[22]), .B2(n_65), .ZN(
      firstInputComplement[22]));
   INV_X1 i_87 (.A(n_63), .ZN(n_62));
   NAND4_X1 i_88 (.A1(n_29), .A2(n_45), .A3(n_57), .A4(n_64), .ZN(n_63));
   NOR3_X1 i_89 (.A1(inputOne[22]), .A2(inputOne[20]), .A3(inputOne[21]), 
      .ZN(n_64));
   INV_X1 i_90 (.A(n_59), .ZN(n_65));
   INV_X1 i_91 (.A(n_66), .ZN(firstInputComplement[25]));
   OAI21_X1 i_92 (.A(n_67), .B1(n_71), .B2(n_68), .ZN(n_66));
   NAND2_X1 i_93 (.A1(n_71), .A2(n_68), .ZN(n_67));
   NOR2_X1 i_94 (.A1(inputOne[24]), .A2(n_69), .ZN(n_68));
   NAND4_X1 i_95 (.A1(n_70), .A2(n_43), .A3(n_57), .A4(n_64), .ZN(n_69));
   INV_X1 i_96 (.A(inputOne[23]), .ZN(n_70));
   INV_X1 i_97 (.A(inputOne[25]), .ZN(n_71));
   AOI21_X1 i_98 (.A(n_72), .B1(inputOne[26]), .B2(n_67), .ZN(
      firstInputComplement[26]));
   NOR2_X1 i_99 (.A1(n_69), .A2(n_73), .ZN(n_72));
   OR3_X1 i_100 (.A1(inputOne[26]), .A2(inputOne[24]), .A3(inputOne[25]), 
      .ZN(n_73));
   AOI21_X1 i_101 (.A(n_74), .B1(inputOne[27]), .B2(n_76), .ZN(
      firstInputComplement[27]));
   NOR3_X1 i_102 (.A1(n_73), .A2(inputOne[27]), .A3(n_69), .ZN(n_74));
   NOR2_X1 i_103 (.A1(n_73), .A2(inputOne[27]), .ZN(n_75));
   INV_X1 i_104 (.A(n_72), .ZN(n_76));
   INV_X1 i_105 (.A(n_69), .ZN(n_77));
   NAND2_X1 i_106 (.A1(n_77), .A2(n_75), .ZN(n_78));
   NOR2_X1 i_107 (.A1(n_78), .A2(inputOne[28]), .ZN(n_79));
   AOI21_X1 i_108 (.A(n_79), .B1(inputOne[28]), .B2(n_78), .ZN(
      firstInputComplement[28]));
   INV_X1 i_109 (.A(n_79), .ZN(n_80));
   AOI22_X1 i_110 (.A1(n_74), .A2(n_82), .B1(inputOne[30]), .B2(n_81), .ZN(
      firstInputComplement[30]));
   NAND3_X1 i_111 (.A1(n_77), .A2(n_75), .A3(n_83), .ZN(n_81));
   NOR3_X1 i_112 (.A1(inputOne[29]), .A2(inputOne[28]), .A3(inputOne[30]), 
      .ZN(n_82));
   NOR2_X1 i_113 (.A1(inputOne[29]), .A2(inputOne[28]), .ZN(n_83));
   AOI21_X1 i_114 (.A(n_84), .B1(inputOne[31]), .B2(n_85), .ZN(
      firstInputComplement[31]));
   AND4_X1 i_115 (.A1(n_86), .A2(n_77), .A3(n_75), .A4(n_82), .ZN(n_84));
   NAND4_X1 i_116 (.A1(n_62), .A2(n_70), .A3(n_75), .A4(n_82), .ZN(n_85));
   INV_X1 i_117 (.A(inputOne[31]), .ZN(n_86));
endmodule

module datapath__0_10(p_0, finalResult, p_1);
   input [63:0]p_0;
   input [63:0]finalResult;
   output [63:0]p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1[0]));
   OAI21_X1 i_1 (.A(n_366), .B1(p_0[0]), .B2(finalResult[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_366), .B(n_1), .Z(p_1[1]));
   OAI21_X1 i_3 (.A(n_365), .B1(p_0[1]), .B2(finalResult[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_364), .B(n_2), .ZN(p_1[2]));
   OAI21_X1 i_5 (.A(n_369), .B1(p_0[2]), .B2(finalResult[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_363), .B(n_3), .Z(p_1[3]));
   OAI21_X1 i_7 (.A(n_370), .B1(n_376), .B2(n_372), .ZN(n_3));
   XOR2_X1 i_8 (.A(n_361), .B(n_10), .Z(p_1[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_1[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_1[6]));
   NOR2_X1 i_11 (.A1(n_358), .A2(n_349), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_1[7]));
   OAI22_X1 i_13 (.A1(p_0[6]), .A2(finalResult[6]), .B1(n_349), .B2(n_7), 
      .ZN(n_5));
   AOI21_X1 i_14 (.A(n_359), .B1(p_0[5]), .B2(finalResult[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_359), .B1(n_353), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_356), .B1(n_361), .B2(n_354), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_354), .B1(p_0[4]), .B2(finalResult[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_360), .A2(n_351), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_347), .B(n_18), .ZN(p_1[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_1[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_1[10]));
   NOR2_X1 i_23 (.A1(n_344), .A2(n_335), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_1[11]));
   OAI22_X1 i_25 (.A1(p_0[10]), .A2(finalResult[10]), .B1(n_335), .B2(n_15), 
      .ZN(n_13));
   AOI21_X1 i_26 (.A(n_345), .B1(p_0[9]), .B2(finalResult[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_345), .B1(n_339), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_342), .B1(n_347), .B2(n_340), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_342), .B1(p_0[8]), .B2(finalResult[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_346), .A2(n_337), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_333), .B(n_26), .Z(p_1[12]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(p_1[13]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(p_1[14]));
   NOR2_X1 i_35 (.A1(n_330), .A2(n_321), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(p_1[15]));
   OAI22_X1 i_37 (.A1(p_0[14]), .A2(finalResult[14]), .B1(n_321), .B2(n_23), 
      .ZN(n_21));
   AOI21_X1 i_38 (.A(n_331), .B1(p_0[13]), .B2(finalResult[13]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_331), .B1(n_325), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_328), .B1(n_333), .B2(n_326), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_326), .B1(p_0[12]), .B2(finalResult[12]), .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_332), .A2(n_323), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_319), .B(n_34), .Z(p_1[16]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(p_1[17]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(p_1[18]));
   NOR2_X1 i_47 (.A1(n_285), .A2(n_275), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(p_1[19]));
   OAI21_X1 i_49 (.A(n_284), .B1(n_275), .B2(n_31), .ZN(n_29));
   NOR2_X1 i_50 (.A1(n_287), .A2(n_277), .ZN(n_30));
   INV_X1 i_51 (.A(n_32), .ZN(n_31));
   OAI21_X1 i_52 (.A(n_286), .B1(n_277), .B2(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_282), .B1(n_319), .B2(n_279), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_279), .B1(p_0[16]), .B2(finalResult[16]), .ZN(n_34));
   AOI21_X1 i_55 (.A(n_289), .B1(p_0[19]), .B2(finalResult[19]), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_63), .B(n_42), .Z(p_1[20]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(p_1[21]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(p_1[22]));
   NOR2_X1 i_59 (.A1(n_313), .A2(n_257), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(p_1[23]));
   OAI21_X1 i_61 (.A(n_312), .B1(n_257), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_315), .A2(n_259), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_314), .B1(n_259), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_318), .B1(n_261), .B2(n_63), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_261), .B1(p_0[20]), .B2(finalResult[20]), .ZN(n_42));
   AOI21_X1 i_67 (.A(n_317), .B1(p_0[23]), .B2(finalResult[23]), .ZN(n_43));
   XOR2_X1 i_68 (.A(n_61), .B(n_50), .Z(p_1[24]));
   XOR2_X1 i_69 (.A(n_49), .B(n_46), .Z(p_1[25]));
   XOR2_X1 i_70 (.A(n_47), .B(n_44), .Z(p_1[26]));
   NOR2_X1 i_71 (.A1(n_296), .A2(n_269), .ZN(n_44));
   XNOR2_X1 i_72 (.A(n_51), .B(n_45), .ZN(p_1[27]));
   OAI21_X1 i_73 (.A(n_295), .B1(n_269), .B2(n_47), .ZN(n_45));
   NOR2_X1 i_74 (.A1(n_298), .A2(n_271), .ZN(n_46));
   INV_X1 i_75 (.A(n_48), .ZN(n_47));
   OAI21_X1 i_76 (.A(n_297), .B1(n_271), .B2(n_49), .ZN(n_48));
   AOI21_X1 i_77 (.A(n_293), .B1(n_273), .B2(n_61), .ZN(n_49));
   OAI21_X1 i_78 (.A(n_273), .B1(p_0[24]), .B2(finalResult[24]), .ZN(n_50));
   AOI21_X1 i_79 (.A(n_300), .B1(p_0[27]), .B2(finalResult[27]), .ZN(n_51));
   XOR2_X1 i_80 (.A(n_59), .B(n_58), .Z(p_1[28]));
   XOR2_X1 i_81 (.A(n_57), .B(n_54), .Z(p_1[29]));
   XOR2_X1 i_82 (.A(n_55), .B(n_52), .Z(p_1[30]));
   NOR2_X1 i_83 (.A1(n_305), .A2(n_263), .ZN(n_52));
   XOR2_X1 i_84 (.A(n_65), .B(n_53), .Z(p_1[31]));
   OAI21_X1 i_85 (.A(n_304), .B1(n_263), .B2(n_55), .ZN(n_53));
   NOR2_X1 i_86 (.A1(n_307), .A2(n_266), .ZN(n_54));
   INV_X1 i_87 (.A(n_56), .ZN(n_55));
   OAI21_X1 i_88 (.A(n_306), .B1(n_266), .B2(n_57), .ZN(n_56));
   AOI21_X1 i_89 (.A(n_302), .B1(n_267), .B2(n_59), .ZN(n_57));
   OAI21_X1 i_90 (.A(n_267), .B1(p_0[28]), .B2(finalResult[28]), .ZN(n_58));
   INV_X1 i_91 (.A(n_60), .ZN(n_59));
   OAI21_X1 i_92 (.A(n_268), .B1(n_292), .B2(n_61), .ZN(n_60));
   INV_X1 i_93 (.A(n_62), .ZN(n_61));
   OAI21_X1 i_94 (.A(n_256), .B1(n_310), .B2(n_63), .ZN(n_62));
   INV_X1 i_95 (.A(n_64), .ZN(n_63));
   OAI21_X1 i_96 (.A(n_274), .B1(n_319), .B2(n_281), .ZN(n_64));
   OAI21_X1 i_97 (.A(n_308), .B1(n_377), .B2(n_373), .ZN(n_65));
   XOR2_X1 i_98 (.A(n_254), .B(n_72), .Z(p_1[32]));
   XOR2_X1 i_99 (.A(n_71), .B(n_68), .Z(p_1[33]));
   XOR2_X1 i_100 (.A(n_69), .B(n_66), .Z(p_1[34]));
   NOR2_X1 i_101 (.A1(n_223), .A2(n_213), .ZN(n_66));
   XNOR2_X1 i_102 (.A(n_73), .B(n_67), .ZN(p_1[35]));
   OAI21_X1 i_103 (.A(n_222), .B1(n_213), .B2(n_69), .ZN(n_67));
   NOR2_X1 i_104 (.A1(n_225), .A2(n_215), .ZN(n_68));
   INV_X1 i_105 (.A(n_70), .ZN(n_69));
   OAI21_X1 i_106 (.A(n_224), .B1(n_215), .B2(n_71), .ZN(n_70));
   AOI21_X1 i_107 (.A(n_220), .B1(n_254), .B2(n_217), .ZN(n_71));
   OAI21_X1 i_108 (.A(n_217), .B1(p_0[32]), .B2(finalResult[32]), .ZN(n_72));
   AOI21_X1 i_109 (.A(n_227), .B1(p_0[35]), .B2(finalResult[35]), .ZN(n_73));
   XOR2_X1 i_110 (.A(n_101), .B(n_80), .Z(p_1[36]));
   XOR2_X1 i_111 (.A(n_79), .B(n_76), .Z(p_1[37]));
   XOR2_X1 i_112 (.A(n_77), .B(n_74), .Z(p_1[38]));
   NOR2_X1 i_113 (.A1(n_248), .A2(n_206), .ZN(n_74));
   XNOR2_X1 i_114 (.A(n_81), .B(n_75), .ZN(p_1[39]));
   OAI21_X1 i_115 (.A(n_247), .B1(n_206), .B2(n_77), .ZN(n_75));
   NOR2_X1 i_116 (.A1(n_250), .A2(n_208), .ZN(n_76));
   INV_X1 i_117 (.A(n_78), .ZN(n_77));
   OAI21_X1 i_118 (.A(n_249), .B1(n_208), .B2(n_79), .ZN(n_78));
   AOI21_X1 i_119 (.A(n_253), .B1(n_210), .B2(n_101), .ZN(n_79));
   OAI21_X1 i_120 (.A(n_210), .B1(p_0[36]), .B2(finalResult[36]), .ZN(n_80));
   AOI21_X1 i_121 (.A(n_252), .B1(p_0[39]), .B2(finalResult[39]), .ZN(n_81));
   XOR2_X1 i_122 (.A(n_99), .B(n_88), .Z(p_1[40]));
   XOR2_X1 i_123 (.A(n_87), .B(n_84), .Z(p_1[41]));
   XOR2_X1 i_124 (.A(n_85), .B(n_82), .Z(p_1[42]));
   NOR2_X1 i_125 (.A1(n_234), .A2(n_192), .ZN(n_82));
   XNOR2_X1 i_126 (.A(n_89), .B(n_83), .ZN(p_1[43]));
   OAI21_X1 i_127 (.A(n_233), .B1(n_192), .B2(n_85), .ZN(n_83));
   NOR2_X1 i_128 (.A1(n_236), .A2(n_194), .ZN(n_84));
   INV_X1 i_129 (.A(n_86), .ZN(n_85));
   OAI21_X1 i_130 (.A(n_235), .B1(n_194), .B2(n_87), .ZN(n_86));
   AOI21_X1 i_131 (.A(n_231), .B1(n_196), .B2(n_99), .ZN(n_87));
   OAI21_X1 i_132 (.A(n_196), .B1(p_0[40]), .B2(finalResult[40]), .ZN(n_88));
   AOI21_X1 i_133 (.A(n_238), .B1(p_0[43]), .B2(finalResult[43]), .ZN(n_89));
   XNOR2_X1 i_134 (.A(n_98), .B(n_97), .ZN(p_1[44]));
   XOR2_X1 i_135 (.A(n_95), .B(n_94), .Z(p_1[45]));
   XNOR2_X1 i_136 (.A(n_91), .B(n_90), .ZN(p_1[46]));
   OAI22_X1 i_137 (.A1(p_0[45]), .A2(finalResult[45]), .B1(n_202), .B2(n_95), 
      .ZN(n_90));
   NOR2_X1 i_138 (.A1(n_242), .A2(n_199), .ZN(n_91));
   XNOR2_X1 i_139 (.A(n_103), .B(n_92), .ZN(p_1[47]));
   OAI21_X1 i_140 (.A(n_93), .B1(n_241), .B2(n_199), .ZN(n_92));
   NAND3_X1 i_141 (.A1(n_200), .A2(n_94), .A3(n_96), .ZN(n_93));
   NOR2_X1 i_142 (.A1(n_243), .A2(n_202), .ZN(n_94));
   INV_X1 i_143 (.A(n_96), .ZN(n_95));
   OAI22_X1 i_144 (.A1(p_0[44]), .A2(finalResult[44]), .B1(n_203), .B2(n_98), 
      .ZN(n_96));
   OAI21_X1 i_145 (.A(n_204), .B1(p_0[44]), .B2(finalResult[44]), .ZN(n_97));
   OAI21_X1 i_146 (.A(n_191), .B1(n_230), .B2(n_99), .ZN(n_98));
   INV_X1 i_147 (.A(n_100), .ZN(n_99));
   OAI21_X1 i_148 (.A(n_205), .B1(n_245), .B2(n_101), .ZN(n_100));
   INV_X1 i_149 (.A(n_102), .ZN(n_101));
   OAI21_X1 i_150 (.A(n_212), .B1(n_254), .B2(n_219), .ZN(n_102));
   AOI21_X1 i_151 (.A(n_244), .B1(p_0[47]), .B2(finalResult[47]), .ZN(n_103));
   XOR2_X1 i_152 (.A(n_189), .B(n_110), .Z(p_1[48]));
   XOR2_X1 i_153 (.A(n_109), .B(n_106), .Z(p_1[49]));
   XOR2_X1 i_154 (.A(n_107), .B(n_104), .Z(p_1[50]));
   NOR2_X1 i_155 (.A1(n_186), .A2(n_177), .ZN(n_104));
   XNOR2_X1 i_156 (.A(n_111), .B(n_105), .ZN(p_1[51]));
   OAI22_X1 i_157 (.A1(p_0[50]), .A2(finalResult[50]), .B1(n_177), .B2(n_107), 
      .ZN(n_105));
   AOI21_X1 i_158 (.A(n_187), .B1(p_0[49]), .B2(finalResult[49]), .ZN(n_106));
   AOI21_X1 i_159 (.A(n_187), .B1(n_181), .B2(n_108), .ZN(n_107));
   INV_X1 i_160 (.A(n_109), .ZN(n_108));
   AOI21_X1 i_161 (.A(n_184), .B1(n_189), .B2(n_182), .ZN(n_109));
   OAI21_X1 i_162 (.A(n_182), .B1(p_0[48]), .B2(finalResult[48]), .ZN(n_110));
   NOR2_X1 i_163 (.A1(n_188), .A2(n_179), .ZN(n_111));
   XOR2_X1 i_164 (.A(n_175), .B(n_118), .Z(p_1[52]));
   XOR2_X1 i_165 (.A(n_117), .B(n_114), .Z(p_1[53]));
   XOR2_X1 i_166 (.A(n_115), .B(n_112), .Z(p_1[54]));
   NOR2_X1 i_167 (.A1(n_164), .A2(n_154), .ZN(n_112));
   XNOR2_X1 i_168 (.A(n_119), .B(n_113), .ZN(p_1[55]));
   OAI21_X1 i_169 (.A(n_163), .B1(n_154), .B2(n_115), .ZN(n_113));
   NOR2_X1 i_170 (.A1(n_166), .A2(n_156), .ZN(n_114));
   INV_X1 i_171 (.A(n_116), .ZN(n_115));
   OAI21_X1 i_172 (.A(n_165), .B1(n_156), .B2(n_117), .ZN(n_116));
   AOI21_X1 i_173 (.A(n_161), .B1(n_175), .B2(n_158), .ZN(n_117));
   OAI21_X1 i_174 (.A(n_158), .B1(p_0[52]), .B2(finalResult[52]), .ZN(n_118));
   AOI21_X1 i_175 (.A(n_168), .B1(p_0[55]), .B2(finalResult[55]), .ZN(n_119));
   XNOR2_X1 i_176 (.A(n_128), .B(n_127), .ZN(p_1[56]));
   XOR2_X1 i_177 (.A(n_125), .B(n_124), .Z(p_1[57]));
   XNOR2_X1 i_178 (.A(n_121), .B(n_120), .ZN(p_1[58]));
   OAI22_X1 i_179 (.A1(p_0[57]), .A2(finalResult[57]), .B1(n_149), .B2(n_125), 
      .ZN(n_120));
   NOR2_X1 i_180 (.A1(n_172), .A2(n_145), .ZN(n_121));
   XNOR2_X1 i_181 (.A(n_129), .B(n_122), .ZN(p_1[59]));
   OAI21_X1 i_182 (.A(n_123), .B1(n_171), .B2(n_145), .ZN(n_122));
   NAND3_X1 i_183 (.A1(n_146), .A2(n_124), .A3(n_126), .ZN(n_123));
   NOR2_X1 i_184 (.A1(n_173), .A2(n_149), .ZN(n_124));
   INV_X1 i_185 (.A(n_126), .ZN(n_125));
   OAI22_X1 i_186 (.A1(p_0[56]), .A2(finalResult[56]), .B1(n_150), .B2(n_128), 
      .ZN(n_126));
   OAI21_X1 i_187 (.A(n_151), .B1(p_0[56]), .B2(finalResult[56]), .ZN(n_127));
   OAI21_X1 i_188 (.A(n_153), .B1(n_175), .B2(n_160), .ZN(n_128));
   AOI21_X1 i_189 (.A(n_174), .B1(p_0[59]), .B2(finalResult[59]), .ZN(n_129));
   XNOR2_X1 i_190 (.A(n_143), .B(n_142), .ZN(p_1[60]));
   AOI22_X1 i_191 (.A1(n_140), .A2(n_136), .B1(n_141), .B2(n_135), .ZN(p_1[61]));
   OAI21_X1 i_200 (.A(n_137), .B1(n_379), .B2(n_375), .ZN(n_136));
   INV_X1 i_209 (.A(n_146), .ZN(n_145));
   NAND2_X1 i_210 (.A1(p_0[58]), .A2(finalResult[58]), .ZN(n_146));
   OAI21_X1 i_212 (.A(n_170), .B1(n_150), .B2(n_149), .ZN(n_148));
   AND2_X1 i_213 (.A1(p_0[57]), .A2(finalResult[57]), .ZN(n_149));
   INV_X1 i_214 (.A(n_151), .ZN(n_150));
   NAND2_X1 i_215 (.A1(p_0[56]), .A2(finalResult[56]), .ZN(n_151));
   AOI221_X1 i_217 (.A(n_155), .B1(p_0[55]), .B2(finalResult[55]), .C1(n_167), 
      .C2(n_154), .ZN(n_153));
   AND2_X1 i_218 (.A1(p_0[54]), .A2(finalResult[54]), .ZN(n_154));
   AOI21_X1 i_219 (.A(n_162), .B1(n_158), .B2(n_157), .ZN(n_155));
   INV_X1 i_220 (.A(n_157), .ZN(n_156));
   NAND2_X1 i_221 (.A1(p_0[53]), .A2(finalResult[53]), .ZN(n_157));
   NAND2_X1 i_222 (.A1(p_0[52]), .A2(finalResult[52]), .ZN(n_158));
   NOR2_X1 i_225 (.A1(p_0[52]), .A2(finalResult[52]), .ZN(n_161));
   NAND3_X1 i_226 (.A1(n_167), .A2(n_163), .A3(n_165), .ZN(n_162));
   INV_X1 i_227 (.A(n_164), .ZN(n_163));
   NOR2_X1 i_228 (.A1(p_0[54]), .A2(finalResult[54]), .ZN(n_164));
   INV_X1 i_229 (.A(n_166), .ZN(n_165));
   NOR2_X1 i_230 (.A1(p_0[53]), .A2(finalResult[53]), .ZN(n_166));
   INV_X1 i_231 (.A(n_168), .ZN(n_167));
   NOR2_X1 i_232 (.A1(p_0[55]), .A2(finalResult[55]), .ZN(n_168));
   NOR3_X1 i_234 (.A1(n_174), .A2(n_172), .A3(n_173), .ZN(n_170));
   NOR2_X1 i_235 (.A1(n_173), .A2(n_172), .ZN(n_171));
   NOR2_X1 i_236 (.A1(p_0[58]), .A2(finalResult[58]), .ZN(n_172));
   NOR2_X1 i_237 (.A1(p_0[57]), .A2(finalResult[57]), .ZN(n_173));
   NOR2_X1 i_238 (.A1(p_0[59]), .A2(finalResult[59]), .ZN(n_174));
   INV_X1 i_241 (.A(n_178), .ZN(n_177));
   NAND2_X1 i_242 (.A1(p_0[50]), .A2(finalResult[50]), .ZN(n_178));
   NAND2_X1 i_245 (.A1(p_0[49]), .A2(finalResult[49]), .ZN(n_181));
   NAND2_X1 i_246 (.A1(p_0[48]), .A2(finalResult[48]), .ZN(n_182));
   NOR2_X1 i_250 (.A1(p_0[50]), .A2(finalResult[50]), .ZN(n_186));
   NOR2_X1 i_251 (.A1(p_0[49]), .A2(finalResult[49]), .ZN(n_187));
   NOR2_X1 i_252 (.A1(p_0[51]), .A2(finalResult[51]), .ZN(n_188));
   INV_X1 i_258 (.A(n_195), .ZN(n_194));
   INV_X1 i_263 (.A(n_200), .ZN(n_199));
   NAND2_X1 i_268 (.A1(p_0[44]), .A2(finalResult[44]), .ZN(n_204));
   INV_X1 i_272 (.A(n_209), .ZN(n_208));
   INV_X1 i_279 (.A(n_216), .ZN(n_215));
   NOR2_X1 i_284 (.A1(p_0[32]), .A2(finalResult[32]), .ZN(n_220));
   OR2_X1 i_294 (.A1(n_232), .A2(n_231), .ZN(n_230));
   NOR2_X1 i_295 (.A1(p_0[40]), .A2(finalResult[40]), .ZN(n_231));
   NOR2_X1 i_305 (.A1(n_243), .A2(n_242), .ZN(n_241));
   OR2_X1 i_309 (.A1(n_253), .A2(n_246), .ZN(n_245));
   NOR2_X1 i_317 (.A1(p_0[36]), .A2(finalResult[36]), .ZN(n_253));
   AND2_X1 i_321 (.A1(p_0[22]), .A2(finalResult[22]), .ZN(n_257));
   AOI21_X1 i_322 (.A(n_311), .B1(n_261), .B2(n_260), .ZN(n_258));
   INV_X1 i_323 (.A(n_260), .ZN(n_259));
   NAND2_X1 i_324 (.A1(p_0[21]), .A2(finalResult[21]), .ZN(n_260));
   NAND2_X1 i_325 (.A1(p_0[20]), .A2(finalResult[20]), .ZN(n_261));
   INV_X1 i_327 (.A(n_264), .ZN(n_263));
   NAND2_X1 i_328 (.A1(p_0[30]), .A2(finalResult[30]), .ZN(n_264));
   AOI21_X1 i_329 (.A(n_266), .B1(p_0[28]), .B2(finalResult[28]), .ZN(n_265));
   AND2_X1 i_330 (.A1(p_0[29]), .A2(finalResult[29]), .ZN(n_266));
   NAND2_X1 i_331 (.A1(p_0[28]), .A2(finalResult[28]), .ZN(n_267));
   AND2_X1 i_333 (.A1(p_0[26]), .A2(finalResult[26]), .ZN(n_269));
   AOI21_X1 i_334 (.A(n_294), .B1(n_273), .B2(n_272), .ZN(n_270));
   INV_X1 i_335 (.A(n_272), .ZN(n_271));
   NAND2_X1 i_336 (.A1(p_0[25]), .A2(finalResult[25]), .ZN(n_272));
   NAND2_X1 i_337 (.A1(p_0[24]), .A2(finalResult[24]), .ZN(n_273));
   AND2_X1 i_339 (.A1(p_0[18]), .A2(finalResult[18]), .ZN(n_275));
   AOI21_X1 i_340 (.A(n_283), .B1(n_279), .B2(n_278), .ZN(n_276));
   INV_X1 i_341 (.A(n_278), .ZN(n_277));
   NAND2_X1 i_342 (.A1(p_0[17]), .A2(finalResult[17]), .ZN(n_278));
   NAND2_X1 i_343 (.A1(p_0[16]), .A2(finalResult[16]), .ZN(n_279));
   NOR2_X1 i_346 (.A1(p_0[16]), .A2(finalResult[16]), .ZN(n_282));
   NAND3_X1 i_347 (.A1(n_288), .A2(n_284), .A3(n_286), .ZN(n_283));
   INV_X1 i_348 (.A(n_285), .ZN(n_284));
   NOR2_X1 i_349 (.A1(p_0[18]), .A2(finalResult[18]), .ZN(n_285));
   INV_X1 i_350 (.A(n_287), .ZN(n_286));
   NOR2_X1 i_351 (.A1(p_0[17]), .A2(finalResult[17]), .ZN(n_287));
   INV_X1 i_352 (.A(n_289), .ZN(n_288));
   NOR2_X1 i_353 (.A1(p_0[19]), .A2(finalResult[19]), .ZN(n_289));
   NOR2_X1 i_357 (.A1(p_0[24]), .A2(finalResult[24]), .ZN(n_293));
   NAND3_X1 i_358 (.A1(n_299), .A2(n_295), .A3(n_297), .ZN(n_294));
   INV_X1 i_359 (.A(n_296), .ZN(n_295));
   NOR2_X1 i_360 (.A1(p_0[26]), .A2(finalResult[26]), .ZN(n_296));
   INV_X1 i_361 (.A(n_298), .ZN(n_297));
   NOR2_X1 i_362 (.A1(p_0[25]), .A2(finalResult[25]), .ZN(n_298));
   INV_X1 i_363 (.A(n_300), .ZN(n_299));
   NOR2_X1 i_364 (.A1(p_0[27]), .A2(finalResult[27]), .ZN(n_300));
   NOR2_X1 i_369 (.A1(p_0[30]), .A2(finalResult[30]), .ZN(n_305));
   NOR2_X1 i_371 (.A1(p_0[29]), .A2(finalResult[29]), .ZN(n_307));
   NAND3_X1 i_375 (.A1(n_316), .A2(n_312), .A3(n_314), .ZN(n_311));
   INV_X1 i_376 (.A(n_313), .ZN(n_312));
   NOR2_X1 i_377 (.A1(p_0[22]), .A2(finalResult[22]), .ZN(n_313));
   INV_X1 i_378 (.A(n_315), .ZN(n_314));
   NOR2_X1 i_379 (.A1(p_0[21]), .A2(finalResult[21]), .ZN(n_315));
   INV_X1 i_380 (.A(n_317), .ZN(n_316));
   NOR2_X1 i_381 (.A1(p_0[23]), .A2(finalResult[23]), .ZN(n_317));
   NOR2_X1 i_382 (.A1(p_0[20]), .A2(finalResult[20]), .ZN(n_318));
   NOR2_X1 i_384 (.A1(n_332), .A2(n_322), .ZN(n_320));
   INV_X1 i_385 (.A(n_322), .ZN(n_321));
   NAND2_X1 i_386 (.A1(p_0[14]), .A2(finalResult[14]), .ZN(n_322));
   AND2_X1 i_387 (.A1(p_0[15]), .A2(finalResult[15]), .ZN(n_323));
   AOI21_X1 i_388 (.A(n_329), .B1(n_326), .B2(n_325), .ZN(n_324));
   NAND2_X1 i_389 (.A1(p_0[13]), .A2(finalResult[13]), .ZN(n_325));
   NAND2_X1 i_390 (.A1(p_0[12]), .A2(finalResult[12]), .ZN(n_326));
   NOR3_X1 i_391 (.A1(n_329), .A2(n_328), .A3(n_333), .ZN(n_327));
   NOR2_X1 i_392 (.A1(p_0[12]), .A2(finalResult[12]), .ZN(n_328));
   OR3_X1 i_393 (.A1(n_332), .A2(n_330), .A3(n_331), .ZN(n_329));
   NOR2_X1 i_394 (.A1(p_0[14]), .A2(finalResult[14]), .ZN(n_330));
   NOR2_X1 i_395 (.A1(p_0[13]), .A2(finalResult[13]), .ZN(n_331));
   NOR2_X1 i_396 (.A1(p_0[15]), .A2(finalResult[15]), .ZN(n_332));
   NOR4_X1 i_397 (.A1(n_337), .A2(n_334), .A3(n_338), .A4(n_341), .ZN(n_333));
   NOR2_X1 i_398 (.A1(n_346), .A2(n_336), .ZN(n_334));
   INV_X1 i_399 (.A(n_336), .ZN(n_335));
   NAND2_X1 i_400 (.A1(p_0[10]), .A2(finalResult[10]), .ZN(n_336));
   AND2_X1 i_401 (.A1(p_0[11]), .A2(finalResult[11]), .ZN(n_337));
   AOI21_X1 i_402 (.A(n_343), .B1(n_340), .B2(n_339), .ZN(n_338));
   NAND2_X1 i_403 (.A1(p_0[9]), .A2(finalResult[9]), .ZN(n_339));
   NAND2_X1 i_404 (.A1(p_0[8]), .A2(finalResult[8]), .ZN(n_340));
   NOR3_X1 i_405 (.A1(n_343), .A2(n_342), .A3(n_347), .ZN(n_341));
   NOR2_X1 i_406 (.A1(p_0[8]), .A2(finalResult[8]), .ZN(n_342));
   OR3_X1 i_407 (.A1(n_346), .A2(n_344), .A3(n_345), .ZN(n_343));
   NOR2_X1 i_408 (.A1(p_0[10]), .A2(finalResult[10]), .ZN(n_344));
   NOR2_X1 i_409 (.A1(p_0[9]), .A2(finalResult[9]), .ZN(n_345));
   NOR2_X1 i_410 (.A1(p_0[11]), .A2(finalResult[11]), .ZN(n_346));
   NOR4_X1 i_411 (.A1(n_351), .A2(n_348), .A3(n_352), .A4(n_355), .ZN(n_347));
   NOR2_X1 i_412 (.A1(n_360), .A2(n_350), .ZN(n_348));
   INV_X1 i_413 (.A(n_350), .ZN(n_349));
   NAND2_X1 i_414 (.A1(p_0[6]), .A2(finalResult[6]), .ZN(n_350));
   AND2_X1 i_415 (.A1(p_0[7]), .A2(finalResult[7]), .ZN(n_351));
   AOI21_X1 i_416 (.A(n_357), .B1(n_354), .B2(n_353), .ZN(n_352));
   NAND2_X1 i_417 (.A1(p_0[5]), .A2(finalResult[5]), .ZN(n_353));
   NAND2_X1 i_418 (.A1(p_0[4]), .A2(finalResult[4]), .ZN(n_354));
   NOR3_X1 i_419 (.A1(n_357), .A2(n_356), .A3(n_361), .ZN(n_355));
   NOR2_X1 i_420 (.A1(p_0[4]), .A2(finalResult[4]), .ZN(n_356));
   OR3_X1 i_421 (.A1(n_360), .A2(n_358), .A3(n_359), .ZN(n_357));
   NOR2_X1 i_422 (.A1(p_0[6]), .A2(finalResult[6]), .ZN(n_358));
   NOR2_X1 i_423 (.A1(p_0[5]), .A2(finalResult[5]), .ZN(n_359));
   NOR2_X1 i_424 (.A1(p_0[7]), .A2(finalResult[7]), .ZN(n_360));
   NAND2_X1 i_425 (.A1(n_370), .A2(n_362), .ZN(n_361));
   OAI21_X1 i_426 (.A(n_363), .B1(n_376), .B2(n_372), .ZN(n_362));
   OAI22_X1 i_427 (.A1(p_0[2]), .A2(finalResult[2]), .B1(n_368), .B2(n_364), 
      .ZN(n_363));
   AOI21_X1 i_428 (.A(n_367), .B1(n_366), .B2(n_365), .ZN(n_364));
   NAND2_X1 i_429 (.A1(p_0[1]), .A2(finalResult[1]), .ZN(n_365));
   NAND2_X1 i_430 (.A1(p_0[0]), .A2(finalResult[0]), .ZN(n_366));
   NOR2_X1 i_431 (.A1(p_0[1]), .A2(finalResult[1]), .ZN(n_367));
   INV_X1 i_432 (.A(n_369), .ZN(n_368));
   NAND2_X1 i_433 (.A1(p_0[2]), .A2(finalResult[2]), .ZN(n_369));
   NAND2_X1 i_434 (.A1(n_376), .A2(n_372), .ZN(n_370));
   INV_X1 i_436 (.A(finalResult[3]), .ZN(n_372));
   INV_X1 i_437 (.A(finalResult[31]), .ZN(n_373));
   INV_X1 i_438 (.A(finalResult[59]), .ZN(n_374));
   INV_X1 i_439 (.A(finalResult[61]), .ZN(n_375));
   INV_X1 i_440 (.A(p_0[3]), .ZN(n_376));
   INV_X1 i_441 (.A(p_0[31]), .ZN(n_377));
   INV_X1 i_442 (.A(p_0[59]), .ZN(n_378));
   INV_X1 i_443 (.A(p_0[61]), .ZN(n_379));
   NAND3_X1 i_192 (.A1(n_412), .A2(n_247), .A3(n_249), .ZN(n_246));
   INV_X1 i_193 (.A(n_136), .ZN(n_135));
   INV_X1 i_194 (.A(n_141), .ZN(n_140));
   NAND2_X1 i_195 (.A1(n_228), .A2(n_479), .ZN(n_141));
   INV_X1 i_196 (.A(n_130), .ZN(n_142));
   NAND2_X1 i_197 (.A1(n_478), .A2(n_479), .ZN(n_130));
   NOR2_X1 i_198 (.A1(n_229), .A2(n_240), .ZN(n_143));
   INV_X1 i_199 (.A(n_131), .ZN(n_175));
   NAND2_X1 i_201 (.A1(n_371), .A2(n_290), .ZN(n_131));
   INV_X1 i_202 (.A(n_301), .ZN(n_179));
   NOR2_X1 i_203 (.A1(p_0[48]), .A2(finalResult[48]), .ZN(n_184));
   INV_X1 i_204 (.A(n_132), .ZN(n_189));
   NAND3_X1 i_205 (.A1(n_415), .A2(n_405), .A3(n_385), .ZN(n_132));
   INV_X1 i_206 (.A(n_133), .ZN(n_212));
   NAND2_X1 i_207 (.A1(n_421), .A2(n_417), .ZN(n_133));
   INV_X1 i_208 (.A(n_406), .ZN(n_205));
   INV_X1 i_211 (.A(n_396), .ZN(n_191));
   INV_X1 i_216 (.A(n_204), .ZN(n_203));
   INV_X1 i_223 (.A(n_472), .ZN(n_243));
   NOR2_X1 i_224 (.A1(p_0[46]), .A2(finalResult[46]), .ZN(n_242));
   INV_X1 i_233 (.A(n_394), .ZN(n_202));
   INV_X1 i_239 (.A(n_235), .ZN(n_236));
   INV_X1 i_240 (.A(n_400), .ZN(n_192));
   INV_X1 i_243 (.A(n_410), .ZN(n_206));
   INV_X1 i_244 (.A(n_224), .ZN(n_225));
   INV_X1 i_247 (.A(n_420), .ZN(n_213));
   NAND2_X1 i_248 (.A1(n_431), .A2(n_432), .ZN(n_310));
   INV_X1 i_249 (.A(n_434), .ZN(n_256));
   INV_X1 i_253 (.A(n_440), .ZN(n_292));
   INV_X1 i_254 (.A(n_447), .ZN(n_268));
   NOR2_X1 i_255 (.A1(p_0[28]), .A2(finalResult[28]), .ZN(n_302));
   INV_X1 i_256 (.A(n_307), .ZN(n_306));
   INV_X1 i_257 (.A(n_305), .ZN(n_304));
   INV_X1 i_259 (.A(n_134), .ZN(p_1[62]));
   NAND2_X1 i_260 (.A1(n_144), .A2(n_138), .ZN(n_134));
   NAND3_X1 i_261 (.A1(n_139), .A2(n_180), .A3(n_169), .ZN(n_138));
   INV_X1 i_262 (.A(n_147), .ZN(n_139));
   OAI21_X1 i_264 (.A(n_176), .B1(n_147), .B2(n_159), .ZN(n_144));
   AOI21_X1 i_265 (.A(n_152), .B1(n_228), .B2(n_479), .ZN(n_147));
   INV_X1 i_266 (.A(n_137), .ZN(n_152));
   INV_X1 i_267 (.A(n_169), .ZN(n_159));
   NAND2_X1 i_269 (.A1(p_0[61]), .A2(finalResult[61]), .ZN(n_169));
   INV_X1 i_270 (.A(n_180), .ZN(n_176));
   NAND2_X1 i_271 (.A1(n_211), .A2(n_226), .ZN(n_180));
   NAND2_X1 i_273 (.A1(n_183), .A2(n_190), .ZN(p_1[63]));
   OAI21_X1 i_274 (.A(n_197), .B1(n_185), .B2(n_207), .ZN(n_183));
   INV_X1 i_275 (.A(n_214), .ZN(n_185));
   NAND3_X1 i_276 (.A1(n_214), .A2(n_201), .A3(n_193), .ZN(n_190));
   INV_X1 i_277 (.A(n_197), .ZN(n_193));
   XNOR2_X1 i_278 (.A(p_0[63]), .B(n_198), .ZN(n_197));
   INV_X1 i_280 (.A(finalResult[63]), .ZN(n_198));
   INV_X1 i_281 (.A(n_207), .ZN(n_201));
   OAI21_X1 i_282 (.A(n_211), .B1(n_137), .B2(n_221), .ZN(n_207));
   NAND2_X1 i_283 (.A1(n_379), .A2(n_375), .ZN(n_137));
   OR2_X1 i_285 (.A1(p_0[62]), .A2(finalResult[62]), .ZN(n_211));
   NAND3_X1 i_286 (.A1(n_228), .A2(n_479), .A3(n_218), .ZN(n_214));
   NOR2_X1 i_287 (.A1(n_136), .A2(n_221), .ZN(n_218));
   INV_X1 i_288 (.A(n_226), .ZN(n_221));
   NAND2_X1 i_289 (.A1(p_0[62]), .A2(finalResult[62]), .ZN(n_226));
   OAI21_X1 i_290 (.A(n_478), .B1(n_229), .B2(n_240), .ZN(n_228));
   OAI21_X1 i_291 (.A(n_237), .B1(n_153), .B2(n_280), .ZN(n_229));
   INV_X1 i_292 (.A(n_239), .ZN(n_237));
   OAI221_X1 i_293 (.A(n_148), .B1(n_146), .B2(n_174), .C1(n_378), .C2(n_374), 
      .ZN(n_239));
   AOI21_X1 i_296 (.A(n_251), .B1(n_371), .B2(n_290), .ZN(n_240));
   OR2_X1 i_297 (.A1(n_160), .A2(n_280), .ZN(n_251));
   NAND2_X1 i_298 (.A1(n_255), .A2(n_262), .ZN(n_160));
   INV_X1 i_299 (.A(n_162), .ZN(n_255));
   INV_X1 i_300 (.A(n_161), .ZN(n_262));
   OAI21_X1 i_301 (.A(n_170), .B1(p_0[56]), .B2(finalResult[56]), .ZN(n_280));
   INV_X1 i_302 (.A(n_291), .ZN(n_290));
   OAI211_X1 i_303 (.A(n_303), .B(n_301), .C1(n_188), .C2(n_178), .ZN(n_291));
   NAND2_X1 i_304 (.A1(p_0[51]), .A2(finalResult[51]), .ZN(n_301));
   NAND2_X1 i_306 (.A1(n_382), .A2(n_309), .ZN(n_303));
   NAND2_X1 i_307 (.A1(n_182), .A2(n_181), .ZN(n_309));
   OAI21_X1 i_308 (.A(n_380), .B1(n_384), .B2(n_414), .ZN(n_371));
   INV_X1 i_310 (.A(n_381), .ZN(n_380));
   OAI21_X1 i_311 (.A(n_382), .B1(p_0[48]), .B2(finalResult[48]), .ZN(n_381));
   INV_X1 i_312 (.A(n_383), .ZN(n_382));
   OR3_X1 i_313 (.A1(n_187), .A2(n_188), .A3(n_186), .ZN(n_383));
   NAND2_X1 i_314 (.A1(n_405), .A2(n_385), .ZN(n_384));
   INV_X1 i_315 (.A(n_386), .ZN(n_385));
   NAND2_X1 i_316 (.A1(n_395), .A2(n_387), .ZN(n_386));
   INV_X1 i_318 (.A(n_388), .ZN(n_387));
   OAI21_X1 i_319 (.A(n_389), .B1(n_468), .B2(n_392), .ZN(n_388));
   INV_X1 i_320 (.A(n_390), .ZN(n_389));
   OAI21_X1 i_326 (.A(n_391), .B1(n_244), .B2(n_200), .ZN(n_390));
   NAND2_X1 i_332 (.A1(p_0[47]), .A2(finalResult[47]), .ZN(n_391));
   NAND2_X1 i_338 (.A1(p_0[46]), .A2(finalResult[46]), .ZN(n_200));
   INV_X1 i_344 (.A(n_469), .ZN(n_244));
   INV_X1 i_345 (.A(n_393), .ZN(n_392));
   NAND2_X1 i_354 (.A1(n_204), .A2(n_394), .ZN(n_393));
   NAND2_X1 i_355 (.A1(p_0[45]), .A2(finalResult[45]), .ZN(n_394));
   NAND2_X1 i_356 (.A1(n_465), .A2(n_396), .ZN(n_395));
   OAI21_X1 i_365 (.A(n_397), .B1(n_232), .B2(n_403), .ZN(n_396));
   INV_X1 i_366 (.A(n_398), .ZN(n_397));
   OAI21_X1 i_367 (.A(n_399), .B1(n_238), .B2(n_400), .ZN(n_398));
   NAND2_X1 i_368 (.A1(p_0[43]), .A2(finalResult[43]), .ZN(n_399));
   NAND2_X1 i_370 (.A1(p_0[42]), .A2(finalResult[42]), .ZN(n_400));
   NOR2_X1 i_372 (.A1(p_0[43]), .A2(finalResult[43]), .ZN(n_238));
   OAI211_X1 i_373 (.A(n_233), .B(n_235), .C1(p_0[43]), .C2(finalResult[43]), 
      .ZN(n_232));
   INV_X1 i_374 (.A(n_234), .ZN(n_233));
   NOR2_X1 i_383 (.A1(p_0[42]), .A2(finalResult[42]), .ZN(n_234));
   NAND2_X1 i_435 (.A1(n_402), .A2(n_401), .ZN(n_235));
   INV_X1 i_444 (.A(finalResult[41]), .ZN(n_401));
   INV_X1 i_445 (.A(p_0[41]), .ZN(n_402));
   INV_X1 i_446 (.A(n_404), .ZN(n_403));
   NAND2_X1 i_447 (.A1(n_196), .A2(n_195), .ZN(n_404));
   NAND2_X1 i_448 (.A1(p_0[41]), .A2(finalResult[41]), .ZN(n_195));
   NAND2_X1 i_449 (.A1(p_0[40]), .A2(finalResult[40]), .ZN(n_196));
   NAND3_X1 i_450 (.A1(n_477), .A2(n_465), .A3(n_406), .ZN(n_405));
   NAND2_X1 i_451 (.A1(n_411), .A2(n_407), .ZN(n_406));
   INV_X1 i_452 (.A(n_408), .ZN(n_407));
   OAI21_X1 i_453 (.A(n_409), .B1(n_252), .B2(n_410), .ZN(n_408));
   NAND2_X1 i_454 (.A1(p_0[39]), .A2(finalResult[39]), .ZN(n_409));
   NAND2_X1 i_455 (.A1(p_0[38]), .A2(finalResult[38]), .ZN(n_410));
   NAND4_X1 i_456 (.A1(n_413), .A2(n_412), .A3(n_247), .A4(n_249), .ZN(n_411));
   INV_X1 i_457 (.A(n_248), .ZN(n_247));
   NOR2_X1 i_458 (.A1(p_0[38]), .A2(finalResult[38]), .ZN(n_248));
   INV_X1 i_459 (.A(n_250), .ZN(n_249));
   NOR2_X1 i_460 (.A1(p_0[37]), .A2(finalResult[37]), .ZN(n_250));
   INV_X1 i_461 (.A(n_252), .ZN(n_412));
   NOR2_X1 i_462 (.A1(p_0[39]), .A2(finalResult[39]), .ZN(n_252));
   NAND2_X1 i_463 (.A1(n_210), .A2(n_209), .ZN(n_413));
   NAND2_X1 i_464 (.A1(p_0[37]), .A2(finalResult[37]), .ZN(n_209));
   NAND2_X1 i_465 (.A1(p_0[36]), .A2(finalResult[36]), .ZN(n_210));
   INV_X1 i_466 (.A(n_415), .ZN(n_414));
   NAND4_X1 i_467 (.A1(n_476), .A2(n_477), .A3(n_465), .A4(n_416), .ZN(n_415));
   OAI211_X1 i_468 (.A(n_421), .B(n_417), .C1(n_219), .C2(n_254), .ZN(n_416));
   INV_X1 i_469 (.A(n_418), .ZN(n_417));
   OAI21_X1 i_470 (.A(n_419), .B1(n_227), .B2(n_420), .ZN(n_418));
   NAND2_X1 i_471 (.A1(p_0[35]), .A2(finalResult[35]), .ZN(n_419));
   NAND2_X1 i_472 (.A1(p_0[34]), .A2(finalResult[34]), .ZN(n_420));
   INV_X1 i_473 (.A(n_459), .ZN(n_227));
   NAND2_X1 i_474 (.A1(n_457), .A2(n_422), .ZN(n_421));
   NAND2_X1 i_475 (.A1(n_217), .A2(n_216), .ZN(n_422));
   NAND2_X1 i_476 (.A1(p_0[33]), .A2(finalResult[33]), .ZN(n_216));
   NAND2_X1 i_477 (.A1(p_0[32]), .A2(finalResult[32]), .ZN(n_217));
   INV_X1 i_478 (.A(n_423), .ZN(n_254));
   NAND4_X1 i_479 (.A1(n_441), .A2(n_433), .A3(n_424), .A4(n_446), .ZN(n_423));
   NAND4_X1 i_480 (.A1(n_453), .A2(n_308), .A3(n_440), .A4(n_425), .ZN(n_424));
   INV_X1 i_481 (.A(n_426), .ZN(n_425));
   NAND3_X1 i_482 (.A1(n_431), .A2(n_432), .A3(n_427), .ZN(n_426));
   OAI21_X1 i_483 (.A(n_274), .B1(n_319), .B2(n_281), .ZN(n_427));
   INV_X1 i_484 (.A(n_428), .ZN(n_274));
   NAND2_X1 i_485 (.A1(n_430), .A2(n_429), .ZN(n_428));
   AOI22_X1 i_486 (.A1(n_288), .A2(n_275), .B1(p_0[19]), .B2(finalResult[19]), 
      .ZN(n_429));
   INV_X1 i_487 (.A(n_276), .ZN(n_430));
   NOR4_X1 i_488 (.A1(n_327), .A2(n_323), .A3(n_320), .A4(n_324), .ZN(n_319));
   OR2_X1 i_489 (.A1(n_283), .A2(n_282), .ZN(n_281));
   INV_X1 i_490 (.A(n_311), .ZN(n_431));
   INV_X1 i_491 (.A(n_318), .ZN(n_432));
   NAND4_X1 i_492 (.A1(n_453), .A2(n_308), .A3(n_440), .A4(n_434), .ZN(n_433));
   OAI221_X1 i_493 (.A(n_436), .B1(n_439), .B2(n_438), .C1(n_437), .C2(n_435), 
      .ZN(n_434));
   INV_X1 i_494 (.A(n_316), .ZN(n_435));
   INV_X1 i_495 (.A(n_258), .ZN(n_436));
   INV_X1 i_496 (.A(n_257), .ZN(n_437));
   INV_X1 i_497 (.A(finalResult[23]), .ZN(n_438));
   INV_X1 i_498 (.A(p_0[23]), .ZN(n_439));
   NOR2_X1 i_499 (.A1(n_294), .A2(n_293), .ZN(n_440));
   INV_X1 i_500 (.A(n_442), .ZN(n_441));
   OAI22_X1 i_501 (.A1(n_443), .A2(n_456), .B1(n_377), .B2(n_373), .ZN(n_442));
   AOI21_X1 i_502 (.A(n_444), .B1(n_455), .B2(n_445), .ZN(n_443));
   INV_X1 i_503 (.A(n_264), .ZN(n_444));
   INV_X1 i_504 (.A(n_265), .ZN(n_445));
   NAND3_X1 i_505 (.A1(n_453), .A2(n_308), .A3(n_447), .ZN(n_446));
   OAI221_X1 i_506 (.A(n_449), .B1(n_452), .B2(n_451), .C1(n_450), .C2(n_448), 
      .ZN(n_447));
   INV_X1 i_507 (.A(n_299), .ZN(n_448));
   INV_X1 i_508 (.A(n_270), .ZN(n_449));
   INV_X1 i_509 (.A(n_269), .ZN(n_450));
   INV_X1 i_510 (.A(finalResult[27]), .ZN(n_451));
   INV_X1 i_511 (.A(p_0[27]), .ZN(n_452));
   INV_X1 i_512 (.A(n_454), .ZN(n_453));
   OAI21_X1 i_513 (.A(n_455), .B1(p_0[28]), .B2(finalResult[28]), .ZN(n_454));
   NOR2_X1 i_514 (.A1(n_305), .A2(n_307), .ZN(n_455));
   INV_X1 i_515 (.A(n_456), .ZN(n_308));
   NOR2_X1 i_516 (.A1(p_0[31]), .A2(finalResult[31]), .ZN(n_456));
   NAND2_X1 i_517 (.A1(n_457), .A2(n_464), .ZN(n_219));
   INV_X1 i_518 (.A(n_458), .ZN(n_457));
   NAND3_X1 i_519 (.A1(n_222), .A2(n_224), .A3(n_459), .ZN(n_458));
   INV_X1 i_520 (.A(n_223), .ZN(n_222));
   NOR2_X1 i_521 (.A1(p_0[34]), .A2(finalResult[34]), .ZN(n_223));
   NAND2_X1 i_522 (.A1(n_461), .A2(n_460), .ZN(n_459));
   INV_X1 i_523 (.A(finalResult[35]), .ZN(n_460));
   INV_X1 i_524 (.A(p_0[35]), .ZN(n_461));
   NAND2_X1 i_525 (.A1(n_463), .A2(n_462), .ZN(n_224));
   INV_X1 i_526 (.A(finalResult[33]), .ZN(n_462));
   INV_X1 i_527 (.A(p_0[33]), .ZN(n_463));
   INV_X1 i_528 (.A(n_220), .ZN(n_464));
   INV_X1 i_529 (.A(n_466), .ZN(n_465));
   NAND2_X1 i_530 (.A1(n_467), .A2(n_475), .ZN(n_466));
   INV_X1 i_531 (.A(n_468), .ZN(n_467));
   OAI211_X1 i_532 (.A(n_469), .B(n_472), .C1(p_0[46]), .C2(finalResult[46]), 
      .ZN(n_468));
   NAND2_X1 i_533 (.A1(n_471), .A2(n_470), .ZN(n_469));
   INV_X1 i_534 (.A(finalResult[47]), .ZN(n_470));
   INV_X1 i_535 (.A(p_0[47]), .ZN(n_471));
   NAND2_X1 i_536 (.A1(n_474), .A2(n_473), .ZN(n_472));
   INV_X1 i_537 (.A(finalResult[45]), .ZN(n_473));
   INV_X1 i_538 (.A(p_0[45]), .ZN(n_474));
   OR2_X1 i_539 (.A1(p_0[44]), .A2(finalResult[44]), .ZN(n_475));
   INV_X1 i_540 (.A(n_245), .ZN(n_476));
   INV_X1 i_541 (.A(n_230), .ZN(n_477));
   OR2_X1 i_542 (.A1(p_0[60]), .A2(finalResult[60]), .ZN(n_478));
   NAND2_X1 i_543 (.A1(p_0[60]), .A2(finalResult[60]), .ZN(n_479));
endmodule

module RadixNoaman(inputOne, inputTwo, finalResult, clk, reset, enable, 
      enableRegisterOutput);
   input [31:0]inputOne;
   input [31:0]inputTwo;
   output [63:0]finalResult;
   input clk;
   input reset;
   input enable;
   output enableRegisterOutput;

   wire [31:0]firstInputComplement;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_1_3;
   wire n_0_1_0;
   wire n_0_1_4;
   wire n_0_1_1;
   wire n_0_1_5;
   wire n_0_1_2;
   wire n_0_1_6;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_1_10;
   wire n_0_1_11;
   wire n_0_1_12;
   wire n_0_1_13;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_1_14;
   wire n_0_1_15;
   wire n_0_1_16;
   wire n_0_1_17;
   wire n_0_1_18;
   wire n_0_259;
   wire n_0_1_19;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_1_20;
   wire n_0_263;
   wire n_0_130;
   wire n_0_129;
   wire n_0_1_21;
   wire n_0_1_22;
   wire n_0_1_23;
   wire n_0_1_24;
   wire n_0_1_25;
   wire n_0_1_26;
   wire n_0_1_27;
   wire n_0_1_28;
   wire n_0_1_29;
   wire n_0_1_30;
   wire n_0_1_31;
   wire n_0_1_32;
   wire n_0_1_33;
   wire n_0_1_34;
   wire n_0_1_35;
   wire n_0_1_36;
   wire n_0_1_37;
   wire n_0_1_38;
   wire n_0_1_39;
   wire n_0_1_40;
   wire n_0_1_41;
   wire n_0_1_42;
   wire n_0_1_43;
   wire n_0_1_44;
   wire n_0_1_45;
   wire n_0_1_46;
   wire n_0_1_47;
   wire n_0_1_48;
   wire n_0_1_49;
   wire n_0_1_50;
   wire n_0_1_51;
   wire n_0_1_52;
   wire n_0_1_53;
   wire n_0_1_54;
   wire n_0_52;
   wire n_0_1_55;
   wire n_0_1_56;
   wire n_0_1_57;
   wire n_0_1_58;
   wire n_0_1_59;
   wire n_0_1_60;
   wire n_0_1_61;
   wire n_0_1_62;
   wire n_0_1_63;
   wire n_0_1_64;
   wire n_0_1_65;
   wire n_0_1_66;
   wire n_0_1_67;
   wire n_0_1_68;
   wire n_0_1_69;
   wire n_0_53;
   wire n_0_1_70;
   wire n_0_1_71;
   wire n_0_1_72;
   wire n_0_1_73;
   wire n_0_1_74;
   wire n_0_1_75;
   wire n_0_54;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_1_78;
   wire n_0_1_79;
   wire n_0_55;
   wire n_0_1_80;
   wire n_0_1_81;
   wire n_0_1_82;
   wire n_0_1_83;
   wire n_0_1_84;
   wire n_0_1_85;
   wire n_0_56;
   wire n_0_1_86;
   wire n_0_1_87;
   wire n_0_1_88;
   wire n_0_1_89;
   wire n_0_1_90;
   wire n_0_57;
   wire n_0_1_91;
   wire n_0_1_92;
   wire n_0_1_93;
   wire n_0_1_94;
   wire n_0_58;
   wire n_0_1_95;
   wire n_0_1_96;
   wire n_0_1_97;
   wire n_0_1_98;
   wire n_0_59;
   wire n_0_1_99;
   wire n_0_1_100;
   wire n_0_1_101;
   wire n_0_1_102;
   wire n_0_1_103;
   wire n_0_1_104;
   wire n_0_1_105;
   wire n_0_1_106;
   wire n_0_60;
   wire n_0_1_107;
   wire n_0_1_108;
   wire n_0_1_109;
   wire n_0_1_110;
   wire n_0_1_111;
   wire n_0_1_112;
   wire n_0_61;
   wire n_0_1_113;
   wire n_0_1_114;
   wire n_0_1_115;
   wire n_0_1_116;
   wire n_0_1_117;
   wire n_0_1_118;
   wire n_0_62;
   wire n_0_1_119;
   wire n_0_1_120;
   wire n_0_1_121;
   wire n_0_1_122;
   wire n_0_1_123;
   wire n_0_1_124;
   wire n_0_63;
   wire n_0_1_125;
   wire n_0_1_126;
   wire n_0_1_127;
   wire n_0_1_128;
   wire n_0_1_129;
   wire n_0_1_130;
   wire n_0_1_131;
   wire n_0_64;
   wire n_0_1_132;
   wire n_0_1_133;
   wire n_0_1_134;
   wire n_0_1_135;
   wire n_0_1_136;
   wire n_0_1_137;
   wire n_0_1_138;
   wire n_0_65;
   wire n_0_1_139;
   wire n_0_1_140;
   wire n_0_1_141;
   wire n_0_1_142;
   wire n_0_1_143;
   wire n_0_1_144;
   wire n_0_1_145;
   wire n_0_66;
   wire n_0_1_146;
   wire n_0_1_147;
   wire n_0_1_148;
   wire n_0_1_149;
   wire n_0_1_150;
   wire n_0_1_151;
   wire n_0_1_152;
   wire n_0_67;
   wire n_0_1_153;
   wire n_0_1_154;
   wire n_0_1_155;
   wire n_0_1_156;
   wire n_0_1_157;
   wire n_0_1_158;
   wire n_0_1_159;
   wire n_0_1_160;
   wire n_0_68;
   wire n_0_1_161;
   wire n_0_1_162;
   wire n_0_1_163;
   wire n_0_1_164;
   wire n_0_1_165;
   wire n_0_1_166;
   wire n_0_1_167;
   wire n_0_1_168;
   wire n_0_69;
   wire n_0_1_169;
   wire n_0_1_170;
   wire n_0_1_171;
   wire n_0_1_172;
   wire n_0_1_173;
   wire n_0_1_174;
   wire n_0_1_175;
   wire n_0_1_176;
   wire n_0_70;
   wire n_0_1_177;
   wire n_0_1_178;
   wire n_0_1_179;
   wire n_0_1_180;
   wire n_0_1_181;
   wire n_0_1_182;
   wire n_0_1_183;
   wire n_0_1_184;
   wire n_0_71;
   wire n_0_1_185;
   wire n_0_1_186;
   wire n_0_1_187;
   wire n_0_1_188;
   wire n_0_1_189;
   wire n_0_1_190;
   wire n_0_1_191;
   wire n_0_1_192;
   wire n_0_72;
   wire n_0_1_193;
   wire n_0_1_194;
   wire n_0_1_195;
   wire n_0_1_196;
   wire n_0_1_197;
   wire n_0_1_198;
   wire n_0_1_199;
   wire n_0_73;
   wire n_0_1_200;
   wire n_0_1_201;
   wire n_0_1_202;
   wire n_0_1_203;
   wire n_0_1_204;
   wire n_0_1_205;
   wire n_0_74;
   wire n_0_1_206;
   wire n_0_1_207;
   wire n_0_1_208;
   wire n_0_1_209;
   wire n_0_1_210;
   wire n_0_1_211;
   wire n_0_75;
   wire n_0_1_212;
   wire n_0_1_213;
   wire n_0_1_214;
   wire n_0_1_215;
   wire n_0_1_216;
   wire n_0_1_217;
   wire n_0_1_218;
   wire n_0_1_219;
   wire n_0_76;
   wire n_0_1_220;
   wire n_0_1_221;
   wire n_0_1_222;
   wire n_0_1_223;
   wire n_0_1_224;
   wire n_0_1_225;
   wire n_0_1_226;
   wire n_0_1_227;
   wire n_0_77;
   wire n_0_1_228;
   wire n_0_1_229;
   wire n_0_1_230;
   wire n_0_1_231;
   wire n_0_1_232;
   wire n_0_1_233;
   wire n_0_1_234;
   wire n_0_1_235;
   wire n_0_78;
   wire n_0_1_236;
   wire n_0_1_237;
   wire n_0_1_238;
   wire n_0_1_239;
   wire n_0_1_240;
   wire n_0_1_241;
   wire n_0_1_242;
   wire n_0_1_243;
   wire n_0_79;
   wire n_0_1_244;
   wire n_0_1_245;
   wire n_0_1_246;
   wire n_0_1_247;
   wire n_0_1_248;
   wire n_0_1_249;
   wire n_0_1_250;
   wire n_0_1_251;
   wire n_0_80;
   wire n_0_1_252;
   wire n_0_1_253;
   wire n_0_1_254;
   wire n_0_1_255;
   wire n_0_1_256;
   wire n_0_1_257;
   wire n_0_1_258;
   wire n_0_1_259;
   wire n_0_81;
   wire n_0_1_260;
   wire n_0_1_261;
   wire n_0_1_262;
   wire n_0_1_263;
   wire n_0_1_264;
   wire n_0_1_265;
   wire n_0_1_266;
   wire n_0_1_267;
   wire n_0_82;
   wire n_0_1_268;
   wire n_0_1_269;
   wire n_0_1_270;
   wire n_0_1_271;
   wire n_0_1_272;
   wire n_0_1_273;
   wire n_0_1_274;
   wire n_0_1_275;
   wire n_0_1_276;
   wire n_0_83;
   wire n_0_1_277;
   wire n_0_1_278;
   wire n_0_1_279;
   wire n_0_84;
   wire n_0_1_280;
   wire n_0_1_281;
   wire n_0_1_282;
   wire n_0_85;
   wire n_0_1_283;
   wire n_0_1_284;
   wire n_0_1_285;
   wire n_0_86;
   wire n_0_1_286;
   wire n_0_1_287;
   wire n_0_1_288;
   wire n_0_87;
   wire n_0_1_289;
   wire n_0_1_290;
   wire n_0_1_291;
   wire n_0_88;
   wire n_0_1_292;
   wire n_0_1_293;
   wire n_0_1_294;
   wire n_0_89;
   wire n_0_1_295;
   wire n_0_1_296;
   wire n_0_1_297;
   wire n_0_90;
   wire n_0_1_298;
   wire n_0_1_299;
   wire n_0_1_300;
   wire n_0_91;
   wire n_0_1_301;
   wire n_0_1_302;
   wire n_0_1_303;
   wire n_0_92;
   wire n_0_1_304;
   wire n_0_1_305;
   wire n_0_1_306;
   wire n_0_93;
   wire n_0_1_307;
   wire n_0_1_308;
   wire n_0_1_309;
   wire n_0_94;
   wire n_0_1_310;
   wire n_0_1_311;
   wire n_0_1_312;
   wire n_0_95;
   wire n_0_1_313;
   wire n_0_1_314;
   wire n_0_1_315;
   wire n_0_96;
   wire n_0_1_316;
   wire n_0_1_317;
   wire n_0_1_318;
   wire n_0_97;
   wire n_0_1_319;
   wire n_0_1_320;
   wire n_0_1_321;
   wire n_0_98;
   wire n_0_1_322;
   wire n_0_1_323;
   wire n_0_1_324;
   wire n_0_99;
   wire n_0_1_325;
   wire n_0_1_326;
   wire n_0_1_327;
   wire n_0_1_328;
   wire n_0_100;
   wire n_0_1_329;
   wire n_0_1_330;
   wire n_0_1_331;
   wire n_0_101;
   wire n_0_1_332;
   wire n_0_1_333;
   wire n_0_1_334;
   wire n_0_102;
   wire n_0_1_335;
   wire n_0_1_336;
   wire n_0_1_337;
   wire n_0_103;
   wire n_0_1_338;
   wire n_0_1_339;
   wire n_0_1_340;
   wire n_0_104;
   wire n_0_1_341;
   wire n_0_1_342;
   wire n_0_1_343;
   wire n_0_105;
   wire n_0_1_344;
   wire n_0_1_345;
   wire n_0_1_346;
   wire n_0_106;
   wire n_0_1_347;
   wire n_0_1_348;
   wire n_0_1_349;
   wire n_0_107;
   wire n_0_1_350;
   wire n_0_1_351;
   wire n_0_1_352;
   wire n_0_1_353;
   wire n_0_108;
   wire n_0_1_354;
   wire n_0_1_355;
   wire n_0_1_356;
   wire n_0_1_357;
   wire n_0_109;
   wire n_0_1_358;
   wire n_0_1_359;
   wire n_0_1_360;
   wire n_0_110;
   wire n_0_1_361;
   wire n_0_1_362;
   wire n_0_1_363;
   wire n_0_111;
   wire n_0_1_364;
   wire n_0_1_365;
   wire n_0_1_366;
   wire n_0_112;
   wire n_0_1_367;
   wire n_0_1_368;
   wire n_0_1_369;
   wire n_0_113;
   wire n_0_1_370;
   wire n_0_1_371;
   wire n_0_1_372;
   wire n_0_114;
   wire n_0_1_373;
   wire n_0_1_374;
   wire n_0_1_375;
   wire n_0_1_376;
   wire n_0_1_377;
   wire n_0_115;
   wire n_0_0;
   wire [4:0]counter;
   wire resetReg;
   wire n_0_264;

   TBUF_X1 i_1 (.A(n_64), .EN(n_0), .Z(finalResult[0]));
   TBUF_X1 i_3 (.A(n_63), .EN(n_0), .Z(finalResult[1]));
   TBUF_X1 i_5 (.A(n_62), .EN(n_0), .Z(finalResult[2]));
   TBUF_X1 i_7 (.A(n_61), .EN(n_0), .Z(finalResult[3]));
   TBUF_X1 i_9 (.A(n_60), .EN(n_0), .Z(finalResult[4]));
   TBUF_X1 i_11 (.A(n_59), .EN(n_0), .Z(finalResult[5]));
   TBUF_X1 i_13 (.A(n_58), .EN(n_0), .Z(finalResult[6]));
   TBUF_X1 i_15 (.A(n_57), .EN(n_0), .Z(finalResult[7]));
   TBUF_X1 i_17 (.A(n_56), .EN(n_0), .Z(finalResult[8]));
   TBUF_X1 i_19 (.A(n_55), .EN(n_0), .Z(finalResult[9]));
   TBUF_X1 i_21 (.A(n_54), .EN(n_0), .Z(finalResult[10]));
   TBUF_X1 i_23 (.A(n_53), .EN(n_0), .Z(finalResult[11]));
   TBUF_X1 i_25 (.A(n_52), .EN(n_0), .Z(finalResult[12]));
   TBUF_X1 i_27 (.A(n_51), .EN(n_0), .Z(finalResult[13]));
   TBUF_X1 i_29 (.A(n_50), .EN(n_0), .Z(finalResult[14]));
   TBUF_X1 i_31 (.A(n_49), .EN(n_0), .Z(finalResult[15]));
   TBUF_X1 i_33 (.A(n_48), .EN(n_0), .Z(finalResult[16]));
   TBUF_X1 i_35 (.A(n_47), .EN(n_0), .Z(finalResult[17]));
   TBUF_X1 i_37 (.A(n_46), .EN(n_0), .Z(finalResult[18]));
   TBUF_X1 i_39 (.A(n_45), .EN(n_0), .Z(finalResult[19]));
   TBUF_X1 i_41 (.A(n_44), .EN(n_0), .Z(finalResult[20]));
   TBUF_X1 i_43 (.A(n_43), .EN(n_0), .Z(finalResult[21]));
   TBUF_X1 i_45 (.A(n_42), .EN(n_0), .Z(finalResult[22]));
   TBUF_X1 i_47 (.A(n_41), .EN(n_0), .Z(finalResult[23]));
   TBUF_X1 i_49 (.A(n_40), .EN(n_0), .Z(finalResult[24]));
   TBUF_X1 i_51 (.A(n_39), .EN(n_0), .Z(finalResult[25]));
   TBUF_X1 i_53 (.A(n_38), .EN(n_0), .Z(finalResult[26]));
   TBUF_X1 i_55 (.A(n_37), .EN(n_0), .Z(finalResult[27]));
   TBUF_X1 i_57 (.A(n_36), .EN(n_0), .Z(finalResult[28]));
   TBUF_X1 i_59 (.A(n_35), .EN(n_0), .Z(finalResult[29]));
   TBUF_X1 i_61 (.A(n_34), .EN(n_0), .Z(finalResult[30]));
   TBUF_X1 i_63 (.A(n_33), .EN(n_0), .Z(finalResult[31]));
   TBUF_X1 i_65 (.A(n_32), .EN(n_0), .Z(finalResult[32]));
   TBUF_X1 i_67 (.A(n_31), .EN(n_0), .Z(finalResult[33]));
   TBUF_X1 i_69 (.A(n_30), .EN(n_0), .Z(finalResult[34]));
   TBUF_X1 i_71 (.A(n_29), .EN(n_0), .Z(finalResult[35]));
   TBUF_X1 i_73 (.A(n_28), .EN(n_0), .Z(finalResult[36]));
   TBUF_X1 i_75 (.A(n_27), .EN(n_0), .Z(finalResult[37]));
   TBUF_X1 i_77 (.A(n_26), .EN(n_0), .Z(finalResult[38]));
   TBUF_X1 i_79 (.A(n_25), .EN(n_0), .Z(finalResult[39]));
   TBUF_X1 i_81 (.A(n_24), .EN(n_0), .Z(finalResult[40]));
   TBUF_X1 i_83 (.A(n_23), .EN(n_0), .Z(finalResult[41]));
   TBUF_X1 i_85 (.A(n_22), .EN(n_0), .Z(finalResult[42]));
   TBUF_X1 i_87 (.A(n_21), .EN(n_0), .Z(finalResult[43]));
   TBUF_X1 i_89 (.A(n_20), .EN(n_0), .Z(finalResult[44]));
   TBUF_X1 i_91 (.A(n_19), .EN(n_0), .Z(finalResult[45]));
   TBUF_X1 i_93 (.A(n_18), .EN(n_0), .Z(finalResult[46]));
   TBUF_X1 i_95 (.A(n_17), .EN(n_0), .Z(finalResult[47]));
   TBUF_X1 i_97 (.A(n_16), .EN(n_0), .Z(finalResult[48]));
   TBUF_X1 i_99 (.A(n_15), .EN(n_0), .Z(finalResult[49]));
   TBUF_X1 i_101 (.A(n_14), .EN(n_0), .Z(finalResult[50]));
   TBUF_X1 i_103 (.A(n_13), .EN(n_0), .Z(finalResult[51]));
   TBUF_X1 i_105 (.A(n_12), .EN(n_0), .Z(finalResult[52]));
   TBUF_X1 i_107 (.A(n_11), .EN(n_0), .Z(finalResult[53]));
   TBUF_X1 i_109 (.A(n_10), .EN(n_0), .Z(finalResult[54]));
   TBUF_X1 i_111 (.A(n_9), .EN(n_0), .Z(finalResult[55]));
   TBUF_X1 i_113 (.A(n_8), .EN(n_0), .Z(finalResult[56]));
   TBUF_X1 i_115 (.A(n_7), .EN(n_0), .Z(finalResult[57]));
   TBUF_X1 i_117 (.A(n_6), .EN(n_0), .Z(finalResult[58]));
   TBUF_X1 i_119 (.A(n_5), .EN(n_0), .Z(finalResult[59]));
   TBUF_X1 i_121 (.A(n_4), .EN(n_0), .Z(finalResult[60]));
   TBUF_X1 i_123 (.A(n_3), .EN(n_0), .Z(finalResult[61]));
   TBUF_X1 i_125 (.A(n_2), .EN(n_0), .Z(finalResult[62]));
   TBUF_X1 i_127 (.A(n_1), .EN(n_0), .Z(finalResult[63]));
   datapath i_0_0 (.firstInputComplement({firstInputComplement[31], 
      firstInputComplement[30], firstInputComplement[29], 
      firstInputComplement[28], firstInputComplement[27], 
      firstInputComplement[26], firstInputComplement[25], 
      firstInputComplement[24], firstInputComplement[23], 
      firstInputComplement[22], firstInputComplement[21], 
      firstInputComplement[20], firstInputComplement[19], 
      firstInputComplement[18], firstInputComplement[17], 
      firstInputComplement[16], firstInputComplement[15], 
      firstInputComplement[14], firstInputComplement[13], 
      firstInputComplement[12], firstInputComplement[11], 
      firstInputComplement[10], firstInputComplement[9], firstInputComplement[8], 
      firstInputComplement[7], firstInputComplement[6], firstInputComplement[5], 
      firstInputComplement[4], firstInputComplement[3], firstInputComplement[2], 
      firstInputComplement[1], uc_0}), .inputOne(inputOne));
   DFF_X1 enableRegisterOutput_reg (.D(enable), .CK(clk), .Q(
      enableRegisterOutput), .QN());
   INV_X1 i_0_128 (.A(enableRegisterOutput), .ZN(n_0));
   DFF_X1 \finalResult_reg[63]  (.D(n_0_194), .CK(clk), .Q(n_1), .QN());
   DFF_X1 \finalResult_reg[62]  (.D(n_0_193), .CK(clk), .Q(n_2), .QN());
   DFF_X1 \finalResult_reg[61]  (.D(n_0_192), .CK(clk), .Q(n_3), .QN());
   DFF_X1 \finalResult_reg[60]  (.D(n_0_191), .CK(clk), .Q(n_4), .QN());
   DFF_X1 \finalResult_reg[59]  (.D(n_0_190), .CK(clk), .Q(n_5), .QN());
   DFF_X1 \finalResult_reg[58]  (.D(n_0_189), .CK(clk), .Q(n_6), .QN());
   DFF_X1 \finalResult_reg[57]  (.D(n_0_188), .CK(clk), .Q(n_7), .QN());
   DFF_X1 \finalResult_reg[56]  (.D(n_0_187), .CK(clk), .Q(n_8), .QN());
   DFF_X1 \finalResult_reg[55]  (.D(n_0_186), .CK(clk), .Q(n_9), .QN());
   DFF_X1 \finalResult_reg[54]  (.D(n_0_185), .CK(clk), .Q(n_10), .QN());
   DFF_X1 \finalResult_reg[53]  (.D(n_0_184), .CK(clk), .Q(n_11), .QN());
   DFF_X1 \finalResult_reg[52]  (.D(n_0_183), .CK(clk), .Q(n_12), .QN());
   DFF_X1 \finalResult_reg[51]  (.D(n_0_182), .CK(clk), .Q(n_13), .QN());
   DFF_X1 \finalResult_reg[50]  (.D(n_0_181), .CK(clk), .Q(n_14), .QN());
   DFF_X1 \finalResult_reg[49]  (.D(n_0_180), .CK(clk), .Q(n_15), .QN());
   DFF_X1 \finalResult_reg[48]  (.D(n_0_179), .CK(clk), .Q(n_16), .QN());
   DFF_X1 \finalResult_reg[47]  (.D(n_0_178), .CK(clk), .Q(n_17), .QN());
   DFF_X1 \finalResult_reg[46]  (.D(n_0_177), .CK(clk), .Q(n_18), .QN());
   DFF_X1 \finalResult_reg[45]  (.D(n_0_176), .CK(clk), .Q(n_19), .QN());
   DFF_X1 \finalResult_reg[44]  (.D(n_0_175), .CK(clk), .Q(n_20), .QN());
   DFF_X1 \finalResult_reg[43]  (.D(n_0_174), .CK(clk), .Q(n_21), .QN());
   DFF_X1 \finalResult_reg[42]  (.D(n_0_173), .CK(clk), .Q(n_22), .QN());
   DFF_X1 \finalResult_reg[41]  (.D(n_0_172), .CK(clk), .Q(n_23), .QN());
   DFF_X1 \finalResult_reg[40]  (.D(n_0_171), .CK(clk), .Q(n_24), .QN());
   DFF_X1 \finalResult_reg[39]  (.D(n_0_170), .CK(clk), .Q(n_25), .QN());
   DFF_X1 \finalResult_reg[38]  (.D(n_0_169), .CK(clk), .Q(n_26), .QN());
   DFF_X1 \finalResult_reg[37]  (.D(n_0_168), .CK(clk), .Q(n_27), .QN());
   DFF_X1 \finalResult_reg[36]  (.D(n_0_167), .CK(clk), .Q(n_28), .QN());
   DFF_X1 \finalResult_reg[35]  (.D(n_0_166), .CK(clk), .Q(n_29), .QN());
   DFF_X1 \finalResult_reg[34]  (.D(n_0_165), .CK(clk), .Q(n_30), .QN());
   DFF_X1 \finalResult_reg[33]  (.D(n_0_164), .CK(clk), .Q(n_31), .QN());
   DFF_X1 \finalResult_reg[32]  (.D(n_0_163), .CK(clk), .Q(n_32), .QN());
   DFF_X1 \finalResult_reg[31]  (.D(n_0_162), .CK(clk), .Q(n_33), .QN());
   DFF_X1 \finalResult_reg[30]  (.D(n_0_161), .CK(clk), .Q(n_34), .QN());
   DFF_X1 \finalResult_reg[29]  (.D(n_0_160), .CK(clk), .Q(n_35), .QN());
   DFF_X1 \finalResult_reg[28]  (.D(n_0_159), .CK(clk), .Q(n_36), .QN());
   DFF_X1 \finalResult_reg[27]  (.D(n_0_158), .CK(clk), .Q(n_37), .QN());
   DFF_X1 \finalResult_reg[26]  (.D(n_0_157), .CK(clk), .Q(n_38), .QN());
   DFF_X1 \finalResult_reg[25]  (.D(n_0_156), .CK(clk), .Q(n_39), .QN());
   DFF_X1 \finalResult_reg[24]  (.D(n_0_155), .CK(clk), .Q(n_40), .QN());
   DFF_X1 \finalResult_reg[23]  (.D(n_0_154), .CK(clk), .Q(n_41), .QN());
   DFF_X1 \finalResult_reg[22]  (.D(n_0_153), .CK(clk), .Q(n_42), .QN());
   DFF_X1 \finalResult_reg[21]  (.D(n_0_152), .CK(clk), .Q(n_43), .QN());
   DFF_X1 \finalResult_reg[20]  (.D(n_0_151), .CK(clk), .Q(n_44), .QN());
   DFF_X1 \finalResult_reg[19]  (.D(n_0_150), .CK(clk), .Q(n_45), .QN());
   DFF_X1 \finalResult_reg[18]  (.D(n_0_149), .CK(clk), .Q(n_46), .QN());
   DFF_X1 \finalResult_reg[17]  (.D(n_0_148), .CK(clk), .Q(n_47), .QN());
   DFF_X1 \finalResult_reg[16]  (.D(n_0_147), .CK(clk), .Q(n_48), .QN());
   DFF_X1 \finalResult_reg[15]  (.D(n_0_146), .CK(clk), .Q(n_49), .QN());
   DFF_X1 \finalResult_reg[14]  (.D(n_0_145), .CK(clk), .Q(n_50), .QN());
   DFF_X1 \finalResult_reg[13]  (.D(n_0_144), .CK(clk), .Q(n_51), .QN());
   DFF_X1 \finalResult_reg[12]  (.D(n_0_143), .CK(clk), .Q(n_52), .QN());
   DFF_X1 \finalResult_reg[11]  (.D(n_0_142), .CK(clk), .Q(n_53), .QN());
   DFF_X1 \finalResult_reg[10]  (.D(n_0_141), .CK(clk), .Q(n_54), .QN());
   DFF_X1 \finalResult_reg[9]  (.D(n_0_140), .CK(clk), .Q(n_55), .QN());
   DFF_X1 \finalResult_reg[8]  (.D(n_0_139), .CK(clk), .Q(n_56), .QN());
   DFF_X1 \finalResult_reg[7]  (.D(n_0_138), .CK(clk), .Q(n_57), .QN());
   DFF_X1 \finalResult_reg[6]  (.D(n_0_137), .CK(clk), .Q(n_58), .QN());
   DFF_X1 \finalResult_reg[5]  (.D(n_0_136), .CK(clk), .Q(n_59), .QN());
   DFF_X1 \finalResult_reg[4]  (.D(n_0_135), .CK(clk), .Q(n_60), .QN());
   DFF_X1 \finalResult_reg[3]  (.D(n_0_134), .CK(clk), .Q(n_61), .QN());
   DFF_X1 \finalResult_reg[2]  (.D(n_0_133), .CK(clk), .Q(n_62), .QN());
   DFF_X1 \finalResult_reg[1]  (.D(n_0_132), .CK(clk), .Q(n_63), .QN());
   DFF_X1 \finalResult_reg[0]  (.D(n_0_131), .CK(clk), .Q(n_64), .QN());
   datapath__0_10 i_0_200 (.p_0({n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, 
      n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, 
      n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, 
      n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, 
      n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, 
      n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, 
      n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, 
      n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52}), .finalResult({n_0_258, 
      n_0_257, n_0_256, n_0_255, n_0_254, n_0_253, n_0_252, n_0_251, n_0_250, 
      n_0_249, n_0_248, n_0_247, n_0_246, n_0_245, n_0_244, n_0_243, n_0_242, 
      n_0_241, n_0_240, n_0_239, n_0_238, n_0_237, n_0_236, n_0_235, n_0_234, 
      n_0_233, n_0_232, n_0_231, n_0_230, n_0_229, n_0_228, n_0_227, n_0_226, 
      n_0_225, n_0_224, n_0_223, n_0_222, n_0_221, n_0_220, n_0_219, n_0_218, 
      n_0_217, n_0_216, n_0_215, n_0_214, n_0_213, n_0_212, n_0_211, n_0_210, 
      n_0_209, n_0_208, n_0_207, n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, 
      n_0_201, n_0_200, n_0_199, n_0_198, n_0_197, n_0_196, n_0_195}), .p_1({
      n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, 
      n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_51, n_0_50, n_0_49, 
      n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, 
      n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, 
      n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, 
      n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, 
      n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, 
      n_0_2, n_0_1}));
   HA_X1 i_0_1_0 (.A(counter[1]), .B(counter[0]), .CO(n_0_1_0), .S(n_0_1_3));
   HA_X1 i_0_1_1 (.A(counter[2]), .B(n_0_1_0), .CO(n_0_1_1), .S(n_0_1_4));
   HA_X1 i_0_1_2 (.A(counter[3]), .B(n_0_1_1), .CO(n_0_1_2), .S(n_0_1_5));
   OAI21_X1 i_0_1_3 (.A(enable), .B1(resetReg), .B2(reset), .ZN(n_0_1_6));
   AND2_X1 i_0_1_4 (.A1(n_0_1_6), .A2(n_0_1), .ZN(n_0_131));
   AND2_X1 i_0_1_5 (.A1(n_0_1_6), .A2(n_0_2), .ZN(n_0_132));
   AND2_X1 i_0_1_6 (.A1(n_0_1_6), .A2(n_0_3), .ZN(n_0_133));
   AND2_X1 i_0_1_7 (.A1(n_0_1_6), .A2(n_0_4), .ZN(n_0_134));
   AND2_X1 i_0_1_8 (.A1(n_0_1_6), .A2(n_0_5), .ZN(n_0_135));
   AND2_X1 i_0_1_9 (.A1(n_0_1_6), .A2(n_0_6), .ZN(n_0_136));
   AND2_X1 i_0_1_10 (.A1(n_0_1_6), .A2(n_0_7), .ZN(n_0_137));
   AND2_X1 i_0_1_11 (.A1(n_0_1_6), .A2(n_0_8), .ZN(n_0_138));
   AND2_X1 i_0_1_12 (.A1(n_0_1_6), .A2(n_0_9), .ZN(n_0_139));
   AND2_X1 i_0_1_13 (.A1(n_0_1_6), .A2(n_0_10), .ZN(n_0_140));
   AND2_X1 i_0_1_14 (.A1(n_0_1_6), .A2(n_0_11), .ZN(n_0_141));
   AND2_X1 i_0_1_15 (.A1(n_0_1_6), .A2(n_0_12), .ZN(n_0_142));
   AND2_X1 i_0_1_16 (.A1(n_0_1_6), .A2(n_0_13), .ZN(n_0_143));
   AND2_X1 i_0_1_17 (.A1(n_0_1_6), .A2(n_0_14), .ZN(n_0_144));
   AND2_X1 i_0_1_18 (.A1(n_0_1_6), .A2(n_0_15), .ZN(n_0_145));
   AND2_X1 i_0_1_19 (.A1(n_0_1_6), .A2(n_0_16), .ZN(n_0_146));
   AND2_X1 i_0_1_20 (.A1(n_0_1_6), .A2(n_0_17), .ZN(n_0_147));
   AND2_X1 i_0_1_21 (.A1(n_0_1_6), .A2(n_0_18), .ZN(n_0_148));
   AND2_X1 i_0_1_22 (.A1(n_0_1_6), .A2(n_0_19), .ZN(n_0_149));
   AND2_X1 i_0_1_23 (.A1(n_0_1_6), .A2(n_0_20), .ZN(n_0_150));
   AND2_X1 i_0_1_24 (.A1(n_0_1_6), .A2(n_0_21), .ZN(n_0_151));
   AND2_X1 i_0_1_25 (.A1(n_0_1_6), .A2(n_0_22), .ZN(n_0_152));
   AND2_X1 i_0_1_26 (.A1(n_0_1_6), .A2(n_0_23), .ZN(n_0_153));
   AND2_X1 i_0_1_27 (.A1(n_0_1_6), .A2(n_0_24), .ZN(n_0_154));
   AND2_X1 i_0_1_28 (.A1(n_0_1_6), .A2(n_0_25), .ZN(n_0_155));
   AND2_X1 i_0_1_29 (.A1(n_0_1_6), .A2(n_0_26), .ZN(n_0_156));
   AND2_X1 i_0_1_30 (.A1(n_0_1_6), .A2(n_0_27), .ZN(n_0_157));
   AND2_X1 i_0_1_31 (.A1(n_0_1_6), .A2(n_0_28), .ZN(n_0_158));
   AND2_X1 i_0_1_32 (.A1(n_0_1_6), .A2(n_0_29), .ZN(n_0_159));
   AND2_X1 i_0_1_33 (.A1(n_0_1_6), .A2(n_0_30), .ZN(n_0_160));
   AND2_X1 i_0_1_34 (.A1(n_0_1_6), .A2(n_0_31), .ZN(n_0_161));
   AND2_X1 i_0_1_35 (.A1(n_0_1_6), .A2(n_0_32), .ZN(n_0_162));
   AND2_X1 i_0_1_36 (.A1(n_0_1_6), .A2(n_0_33), .ZN(n_0_163));
   AND2_X1 i_0_1_37 (.A1(n_0_1_6), .A2(n_0_34), .ZN(n_0_164));
   AND2_X1 i_0_1_38 (.A1(n_0_1_6), .A2(n_0_35), .ZN(n_0_165));
   AND2_X1 i_0_1_39 (.A1(n_0_1_6), .A2(n_0_36), .ZN(n_0_166));
   AND2_X1 i_0_1_40 (.A1(n_0_1_6), .A2(n_0_37), .ZN(n_0_167));
   AND2_X1 i_0_1_41 (.A1(n_0_1_6), .A2(n_0_38), .ZN(n_0_168));
   AND2_X1 i_0_1_42 (.A1(n_0_1_6), .A2(n_0_39), .ZN(n_0_169));
   AND2_X1 i_0_1_43 (.A1(n_0_1_6), .A2(n_0_40), .ZN(n_0_170));
   AND2_X1 i_0_1_44 (.A1(n_0_1_6), .A2(n_0_41), .ZN(n_0_171));
   AND2_X1 i_0_1_45 (.A1(n_0_1_6), .A2(n_0_42), .ZN(n_0_172));
   AND2_X1 i_0_1_46 (.A1(n_0_1_6), .A2(n_0_43), .ZN(n_0_173));
   AND2_X1 i_0_1_47 (.A1(n_0_1_6), .A2(n_0_44), .ZN(n_0_174));
   AND2_X1 i_0_1_48 (.A1(n_0_1_6), .A2(n_0_45), .ZN(n_0_175));
   AND2_X1 i_0_1_49 (.A1(n_0_1_6), .A2(n_0_46), .ZN(n_0_176));
   AND2_X1 i_0_1_50 (.A1(n_0_1_6), .A2(n_0_47), .ZN(n_0_177));
   AND2_X1 i_0_1_51 (.A1(n_0_1_6), .A2(n_0_48), .ZN(n_0_178));
   AND2_X1 i_0_1_52 (.A1(n_0_1_6), .A2(n_0_49), .ZN(n_0_179));
   AND2_X1 i_0_1_53 (.A1(n_0_1_6), .A2(n_0_50), .ZN(n_0_180));
   AND2_X1 i_0_1_54 (.A1(n_0_1_6), .A2(n_0_51), .ZN(n_0_181));
   AND2_X1 i_0_1_55 (.A1(n_0_1_6), .A2(n_0_116), .ZN(n_0_182));
   AND2_X1 i_0_1_56 (.A1(n_0_1_6), .A2(n_0_117), .ZN(n_0_183));
   AND2_X1 i_0_1_57 (.A1(n_0_1_6), .A2(n_0_118), .ZN(n_0_184));
   AND2_X1 i_0_1_58 (.A1(n_0_1_6), .A2(n_0_119), .ZN(n_0_185));
   AND2_X1 i_0_1_59 (.A1(n_0_1_6), .A2(n_0_120), .ZN(n_0_186));
   AND2_X1 i_0_1_60 (.A1(n_0_1_6), .A2(n_0_121), .ZN(n_0_187));
   AND2_X1 i_0_1_61 (.A1(n_0_1_6), .A2(n_0_122), .ZN(n_0_188));
   AND2_X1 i_0_1_62 (.A1(n_0_1_6), .A2(n_0_123), .ZN(n_0_189));
   AND2_X1 i_0_1_63 (.A1(n_0_1_6), .A2(n_0_124), .ZN(n_0_190));
   AND2_X1 i_0_1_64 (.A1(n_0_1_6), .A2(n_0_125), .ZN(n_0_191));
   AND2_X1 i_0_1_65 (.A1(n_0_1_6), .A2(n_0_126), .ZN(n_0_192));
   AND2_X1 i_0_1_66 (.A1(n_0_1_6), .A2(n_0_127), .ZN(n_0_193));
   AND2_X1 i_0_1_67 (.A1(n_0_1_6), .A2(n_0_128), .ZN(n_0_194));
   INV_X1 i_0_1_68 (.A(counter[2]), .ZN(n_0_1_7));
   INV_X1 i_0_1_69 (.A(counter[4]), .ZN(n_0_1_8));
   INV_X1 i_0_1_70 (.A(counter[3]), .ZN(n_0_1_9));
   NAND3_X1 i_0_1_71 (.A1(n_0_1_7), .A2(n_0_1_8), .A3(n_0_1_9), .ZN(n_0_1_10));
   NOR2_X1 i_0_1_72 (.A1(n_0_1_10), .A2(counter[1]), .ZN(n_0_1_11));
   INV_X1 i_0_1_73 (.A(counter[0]), .ZN(n_0_1_12));
   NAND2_X1 i_0_1_74 (.A1(n_0_1_11), .A2(n_0_1_12), .ZN(n_0_1_13));
   AND2_X1 i_0_1_75 (.A1(n_0_1_13), .A2(finalResult[0]), .ZN(n_0_195));
   AND2_X1 i_0_1_76 (.A1(n_0_1_13), .A2(finalResult[1]), .ZN(n_0_196));
   AND2_X1 i_0_1_77 (.A1(n_0_1_13), .A2(finalResult[2]), .ZN(n_0_197));
   AND2_X1 i_0_1_78 (.A1(n_0_1_13), .A2(finalResult[3]), .ZN(n_0_198));
   AND2_X1 i_0_1_79 (.A1(n_0_1_13), .A2(finalResult[4]), .ZN(n_0_199));
   AND2_X1 i_0_1_80 (.A1(n_0_1_13), .A2(finalResult[5]), .ZN(n_0_200));
   AND2_X1 i_0_1_81 (.A1(n_0_1_13), .A2(finalResult[6]), .ZN(n_0_201));
   AND2_X1 i_0_1_82 (.A1(n_0_1_13), .A2(finalResult[7]), .ZN(n_0_202));
   AND2_X1 i_0_1_83 (.A1(n_0_1_13), .A2(finalResult[8]), .ZN(n_0_203));
   AND2_X1 i_0_1_84 (.A1(n_0_1_13), .A2(finalResult[9]), .ZN(n_0_204));
   AND2_X1 i_0_1_85 (.A1(n_0_1_13), .A2(finalResult[10]), .ZN(n_0_205));
   AND2_X1 i_0_1_86 (.A1(n_0_1_13), .A2(finalResult[11]), .ZN(n_0_206));
   AND2_X1 i_0_1_87 (.A1(n_0_1_13), .A2(finalResult[12]), .ZN(n_0_207));
   AND2_X1 i_0_1_88 (.A1(n_0_1_13), .A2(finalResult[13]), .ZN(n_0_208));
   AND2_X1 i_0_1_89 (.A1(n_0_1_13), .A2(finalResult[14]), .ZN(n_0_209));
   AND2_X1 i_0_1_90 (.A1(n_0_1_13), .A2(finalResult[15]), .ZN(n_0_210));
   AND2_X1 i_0_1_91 (.A1(n_0_1_13), .A2(finalResult[16]), .ZN(n_0_211));
   AND2_X1 i_0_1_92 (.A1(n_0_1_13), .A2(finalResult[17]), .ZN(n_0_212));
   AND2_X1 i_0_1_93 (.A1(n_0_1_13), .A2(finalResult[18]), .ZN(n_0_213));
   AND2_X1 i_0_1_94 (.A1(n_0_1_13), .A2(finalResult[19]), .ZN(n_0_214));
   AND2_X1 i_0_1_95 (.A1(n_0_1_13), .A2(finalResult[20]), .ZN(n_0_215));
   AND2_X1 i_0_1_96 (.A1(n_0_1_13), .A2(finalResult[21]), .ZN(n_0_216));
   AND2_X1 i_0_1_97 (.A1(n_0_1_13), .A2(finalResult[22]), .ZN(n_0_217));
   AND2_X1 i_0_1_98 (.A1(n_0_1_13), .A2(finalResult[23]), .ZN(n_0_218));
   AND2_X1 i_0_1_99 (.A1(n_0_1_13), .A2(finalResult[24]), .ZN(n_0_219));
   AND2_X1 i_0_1_100 (.A1(n_0_1_13), .A2(finalResult[25]), .ZN(n_0_220));
   AND2_X1 i_0_1_101 (.A1(n_0_1_13), .A2(finalResult[26]), .ZN(n_0_221));
   AND2_X1 i_0_1_102 (.A1(n_0_1_13), .A2(finalResult[27]), .ZN(n_0_222));
   AND2_X1 i_0_1_103 (.A1(n_0_1_13), .A2(finalResult[28]), .ZN(n_0_223));
   AND2_X1 i_0_1_104 (.A1(n_0_1_13), .A2(finalResult[29]), .ZN(n_0_224));
   AND2_X1 i_0_1_105 (.A1(n_0_1_13), .A2(finalResult[30]), .ZN(n_0_225));
   AND2_X1 i_0_1_106 (.A1(n_0_1_13), .A2(finalResult[31]), .ZN(n_0_226));
   AND2_X1 i_0_1_107 (.A1(n_0_1_13), .A2(finalResult[32]), .ZN(n_0_227));
   AND2_X1 i_0_1_108 (.A1(n_0_1_13), .A2(finalResult[33]), .ZN(n_0_228));
   AND2_X1 i_0_1_109 (.A1(n_0_1_13), .A2(finalResult[34]), .ZN(n_0_229));
   AND2_X1 i_0_1_110 (.A1(n_0_1_13), .A2(finalResult[35]), .ZN(n_0_230));
   AND2_X1 i_0_1_111 (.A1(n_0_1_13), .A2(finalResult[36]), .ZN(n_0_231));
   AND2_X1 i_0_1_112 (.A1(n_0_1_13), .A2(finalResult[37]), .ZN(n_0_232));
   AND2_X1 i_0_1_113 (.A1(n_0_1_13), .A2(finalResult[38]), .ZN(n_0_233));
   AND2_X1 i_0_1_114 (.A1(n_0_1_13), .A2(finalResult[39]), .ZN(n_0_234));
   AND2_X1 i_0_1_115 (.A1(n_0_1_13), .A2(finalResult[40]), .ZN(n_0_235));
   AND2_X1 i_0_1_116 (.A1(n_0_1_13), .A2(finalResult[41]), .ZN(n_0_236));
   AND2_X1 i_0_1_117 (.A1(n_0_1_13), .A2(finalResult[42]), .ZN(n_0_237));
   AND2_X1 i_0_1_118 (.A1(n_0_1_13), .A2(finalResult[43]), .ZN(n_0_238));
   AND2_X1 i_0_1_119 (.A1(n_0_1_13), .A2(finalResult[44]), .ZN(n_0_239));
   AND2_X1 i_0_1_120 (.A1(n_0_1_13), .A2(finalResult[45]), .ZN(n_0_240));
   AND2_X1 i_0_1_121 (.A1(n_0_1_13), .A2(finalResult[46]), .ZN(n_0_241));
   AND2_X1 i_0_1_122 (.A1(n_0_1_13), .A2(finalResult[47]), .ZN(n_0_242));
   AND2_X1 i_0_1_123 (.A1(n_0_1_13), .A2(finalResult[48]), .ZN(n_0_243));
   AND2_X1 i_0_1_124 (.A1(n_0_1_13), .A2(finalResult[49]), .ZN(n_0_244));
   AND2_X1 i_0_1_125 (.A1(n_0_1_13), .A2(finalResult[50]), .ZN(n_0_245));
   AND2_X1 i_0_1_126 (.A1(n_0_1_13), .A2(finalResult[51]), .ZN(n_0_246));
   AND2_X1 i_0_1_127 (.A1(n_0_1_13), .A2(finalResult[52]), .ZN(n_0_247));
   AND2_X1 i_0_1_128 (.A1(n_0_1_13), .A2(finalResult[53]), .ZN(n_0_248));
   AND2_X1 i_0_1_129 (.A1(n_0_1_13), .A2(finalResult[54]), .ZN(n_0_249));
   AND2_X1 i_0_1_130 (.A1(n_0_1_13), .A2(finalResult[55]), .ZN(n_0_250));
   AND2_X1 i_0_1_131 (.A1(n_0_1_13), .A2(finalResult[56]), .ZN(n_0_251));
   AND2_X1 i_0_1_132 (.A1(n_0_1_13), .A2(finalResult[57]), .ZN(n_0_252));
   AND2_X1 i_0_1_133 (.A1(n_0_1_13), .A2(finalResult[58]), .ZN(n_0_253));
   AND2_X1 i_0_1_134 (.A1(n_0_1_13), .A2(finalResult[59]), .ZN(n_0_254));
   AND2_X1 i_0_1_135 (.A1(n_0_1_13), .A2(finalResult[60]), .ZN(n_0_255));
   AND2_X1 i_0_1_136 (.A1(n_0_1_13), .A2(finalResult[61]), .ZN(n_0_256));
   AND2_X1 i_0_1_137 (.A1(n_0_1_13), .A2(finalResult[62]), .ZN(n_0_257));
   AND2_X1 i_0_1_138 (.A1(n_0_1_13), .A2(finalResult[63]), .ZN(n_0_258));
   NOR2_X1 i_0_1_139 (.A1(n_0_1_8), .A2(counter[3]), .ZN(n_0_1_14));
   INV_X1 i_0_1_140 (.A(counter[1]), .ZN(n_0_1_15));
   NAND3_X1 i_0_1_141 (.A1(n_0_1_14), .A2(enable), .A3(n_0_1_15), .ZN(n_0_1_16));
   NAND2_X1 i_0_1_142 (.A1(n_0_1_7), .A2(n_0_1_12), .ZN(n_0_1_17));
   OAI21_X1 i_0_1_143 (.A(n_0_1_6), .B1(n_0_1_16), .B2(n_0_1_17), .ZN(n_0_1_18));
   NOR2_X1 i_0_1_144 (.A1(n_0_1_18), .A2(counter[0]), .ZN(n_0_259));
   INV_X1 i_0_1_145 (.A(n_0_1_18), .ZN(n_0_1_19));
   AND2_X1 i_0_1_146 (.A1(n_0_1_19), .A2(n_0_1_3), .ZN(n_0_260));
   AND2_X1 i_0_1_147 (.A1(n_0_1_19), .A2(n_0_1_4), .ZN(n_0_261));
   AND2_X1 i_0_1_148 (.A1(n_0_1_19), .A2(n_0_1_5), .ZN(n_0_262));
   INV_X1 i_0_1_149 (.A(n_0_1_2), .ZN(n_0_1_20));
   AOI221_X1 i_0_1_150 (.A(n_0_1_18), .B1(n_0_1_20), .B2(n_0_1_8), .C1(n_0_1_2), 
      .C2(counter[4]), .ZN(n_0_263));
   INV_X1 i_0_1_151 (.A(n_0_1_6), .ZN(n_0_130));
   AND2_X1 i_0_1_152 (.A1(enable), .A2(reset), .ZN(n_0_129));
   NOR2_X1 i_0_1_153 (.A1(counter[3]), .A2(counter[1]), .ZN(n_0_1_21));
   NOR2_X1 i_0_1_154 (.A1(n_0_1_15), .A2(counter[3]), .ZN(n_0_1_22));
   AOI221_X1 i_0_1_155 (.A(counter[0]), .B1(n_0_1_21), .B2(inputTwo[8]), 
      .C1(n_0_1_22), .C2(inputTwo[12]), .ZN(n_0_1_23));
   NOR2_X1 i_0_1_156 (.A1(n_0_1_9), .A2(n_0_1_15), .ZN(n_0_1_24));
   NOR2_X1 i_0_1_157 (.A1(n_0_1_9), .A2(counter[1]), .ZN(n_0_1_25));
   AOI22_X1 i_0_1_158 (.A1(inputTwo[28]), .A2(n_0_1_24), .B1(n_0_1_25), .B2(
      inputTwo[24]), .ZN(n_0_1_26));
   NAND2_X1 i_0_1_159 (.A1(n_0_1_23), .A2(n_0_1_26), .ZN(n_0_1_27));
   AOI22_X1 i_0_1_160 (.A1(inputTwo[30]), .A2(n_0_1_24), .B1(n_0_1_25), .B2(
      inputTwo[26]), .ZN(n_0_1_28));
   AOI22_X1 i_0_1_161 (.A1(n_0_1_22), .A2(inputTwo[14]), .B1(n_0_1_21), .B2(
      inputTwo[10]), .ZN(n_0_1_29));
   NAND3_X1 i_0_1_162 (.A1(n_0_1_28), .A2(n_0_1_29), .A3(counter[0]), .ZN(
      n_0_1_30));
   AOI21_X1 i_0_1_163 (.A(n_0_1_7), .B1(n_0_1_27), .B2(n_0_1_30), .ZN(n_0_1_31));
   AOI211_X1 i_0_1_164 (.A(counter[2]), .B(n_0_1_12), .C1(n_0_1_24), .C2(
      inputTwo[22]), .ZN(n_0_1_32));
   AOI222_X1 i_0_1_165 (.A1(n_0_1_25), .A2(inputTwo[18]), .B1(n_0_1_22), 
      .B2(inputTwo[6]), .C1(n_0_1_21), .C2(inputTwo[2]), .ZN(n_0_1_33));
   AOI21_X1 i_0_1_166 (.A(n_0_1_17), .B1(n_0_1_24), .B2(inputTwo[20]), .ZN(
      n_0_1_34));
   AOI222_X1 i_0_1_167 (.A1(n_0_1_25), .A2(inputTwo[16]), .B1(n_0_1_22), 
      .B2(inputTwo[4]), .C1(n_0_1_21), .C2(inputTwo[0]), .ZN(n_0_1_35));
   AOI221_X1 i_0_1_168 (.A(n_0_1_31), .B1(n_0_1_32), .B2(n_0_1_33), .C1(n_0_1_34), 
      .C2(n_0_1_35), .ZN(n_0_1_36));
   INV_X1 i_0_1_169 (.A(n_0_1_36), .ZN(n_0_1_37));
   AOI22_X1 i_0_1_170 (.A1(n_0_1_25), .A2(inputTwo[17]), .B1(n_0_1_22), .B2(
      inputTwo[5]), .ZN(n_0_1_38));
   AOI22_X1 i_0_1_171 (.A1(n_0_1_24), .A2(inputTwo[21]), .B1(n_0_1_21), .B2(
      inputTwo[1]), .ZN(n_0_1_39));
   NAND2_X1 i_0_1_172 (.A1(n_0_1_38), .A2(n_0_1_39), .ZN(n_0_1_40));
   NAND3_X1 i_0_1_173 (.A1(n_0_1_40), .A2(n_0_1_7), .A3(counter[0]), .ZN(
      n_0_1_41));
   AOI222_X1 i_0_1_174 (.A1(n_0_1_24), .A2(inputTwo[19]), .B1(n_0_1_22), 
      .B2(inputTwo[3]), .C1(n_0_1_25), .C2(inputTwo[15]), .ZN(n_0_1_42));
   AOI22_X1 i_0_1_175 (.A1(inputTwo[27]), .A2(n_0_1_24), .B1(n_0_1_25), .B2(
      inputTwo[23]), .ZN(n_0_1_43));
   AOI22_X1 i_0_1_176 (.A1(n_0_1_22), .A2(inputTwo[11]), .B1(n_0_1_21), .B2(
      inputTwo[7]), .ZN(n_0_1_44));
   AOI21_X1 i_0_1_177 (.A(counter[0]), .B1(n_0_1_43), .B2(n_0_1_44), .ZN(
      n_0_1_45));
   AOI22_X1 i_0_1_178 (.A1(n_0_1_24), .A2(inputTwo[29]), .B1(n_0_1_25), .B2(
      inputTwo[25]), .ZN(n_0_1_46));
   AOI22_X1 i_0_1_179 (.A1(inputTwo[13]), .A2(n_0_1_22), .B1(n_0_1_21), .B2(
      inputTwo[9]), .ZN(n_0_1_47));
   NAND2_X1 i_0_1_180 (.A1(n_0_1_46), .A2(n_0_1_47), .ZN(n_0_1_48));
   AOI21_X1 i_0_1_181 (.A(n_0_1_45), .B1(counter[0]), .B2(n_0_1_48), .ZN(
      n_0_1_49));
   OAI221_X1 i_0_1_182 (.A(n_0_1_41), .B1(n_0_1_42), .B2(n_0_1_17), .C1(n_0_1_49), 
      .C2(n_0_1_7), .ZN(n_0_1_50));
   INV_X1 i_0_1_183 (.A(n_0_1_50), .ZN(n_0_1_51));
   OAI22_X1 i_0_1_184 (.A1(n_0_1_37), .A2(n_0_1_51), .B1(n_0_1_36), .B2(n_0_1_50), 
      .ZN(n_0_1_52));
   INV_X1 i_0_1_185 (.A(inputOne[0]), .ZN(n_0_1_53));
   OR2_X1 i_0_1_186 (.A1(n_0_1_52), .A2(n_0_1_53), .ZN(n_0_1_54));
   NOR2_X1 i_0_1_187 (.A1(n_0_1_54), .A2(n_0_1_13), .ZN(n_0_52));
   AOI222_X1 i_0_1_188 (.A1(inputTwo[27]), .A2(n_0_1_25), .B1(n_0_1_22), 
      .B2(inputTwo[15]), .C1(n_0_1_21), .C2(inputTwo[11]), .ZN(n_0_1_55));
   AOI21_X1 i_0_1_189 (.A(n_0_1_7), .B1(n_0_1_24), .B2(inputTwo[31]), .ZN(
      n_0_1_56));
   AOI221_X1 i_0_1_190 (.A(counter[2]), .B1(n_0_1_21), .B2(inputTwo[3]), 
      .C1(inputTwo[23]), .C2(n_0_1_24), .ZN(n_0_1_57));
   AOI22_X1 i_0_1_191 (.A1(n_0_1_22), .A2(inputTwo[7]), .B1(n_0_1_25), .B2(
      inputTwo[19]), .ZN(n_0_1_58));
   AOI22_X1 i_0_1_192 (.A1(n_0_1_55), .A2(n_0_1_56), .B1(n_0_1_57), .B2(n_0_1_58), 
      .ZN(n_0_1_59));
   NAND2_X1 i_0_1_193 (.A1(n_0_1_12), .A2(counter[2]), .ZN(n_0_1_60));
   OAI222_X1 i_0_1_194 (.A1(n_0_1_59), .A2(n_0_1_12), .B1(n_0_1_48), .B2(
      n_0_1_60), .C1(n_0_1_17), .C2(n_0_1_40), .ZN(n_0_1_61));
   NOR3_X1 i_0_1_195 (.A1(n_0_1_36), .A2(n_0_1_50), .A3(n_0_1_61), .ZN(n_0_1_62));
   INV_X1 i_0_1_196 (.A(n_0_1_62), .ZN(n_0_1_63));
   NAND3_X1 i_0_1_197 (.A1(n_0_1_36), .A2(n_0_1_50), .A3(n_0_1_61), .ZN(n_0_1_64));
   AOI21_X1 i_0_1_198 (.A(n_0_1_53), .B1(n_0_1_63), .B2(n_0_1_64), .ZN(n_0_1_65));
   NOR2_X1 i_0_1_199 (.A1(n_0_1_52), .A2(n_0_1_61), .ZN(n_0_1_66));
   INV_X1 i_0_1_200 (.A(n_0_1_61), .ZN(n_0_1_67));
   NOR2_X1 i_0_1_201 (.A1(n_0_1_52), .A2(n_0_1_67), .ZN(n_0_1_68));
   AOI221_X1 i_0_1_202 (.A(n_0_1_65), .B1(n_0_1_66), .B2(firstInputComplement[1]), 
      .C1(inputOne[1]), .C2(n_0_1_68), .ZN(n_0_1_69));
   NOR2_X1 i_0_1_203 (.A1(n_0_1_69), .A2(n_0_1_13), .ZN(n_0_53));
   INV_X1 i_0_1_204 (.A(n_0_1_64), .ZN(n_0_1_70));
   AOI22_X1 i_0_1_205 (.A1(n_0_1_68), .A2(inputOne[2]), .B1(n_0_1_70), .B2(
      inputOne[1]), .ZN(n_0_1_71));
   AOI22_X1 i_0_1_206 (.A1(n_0_1_66), .A2(firstInputComplement[2]), .B1(
      firstInputComplement[1]), .B2(n_0_1_62), .ZN(n_0_1_72));
   NAND2_X1 i_0_1_207 (.A1(n_0_1_71), .A2(n_0_1_72), .ZN(n_0_1_73));
   INV_X1 i_0_1_208 (.A(n_0_1_73), .ZN(n_0_1_74));
   NAND2_X1 i_0_1_209 (.A1(n_0_1_11), .A2(counter[0]), .ZN(n_0_1_75));
   OAI22_X1 i_0_1_210 (.A1(n_0_1_74), .A2(n_0_1_13), .B1(n_0_1_54), .B2(n_0_1_75), 
      .ZN(n_0_54));
   AOI22_X1 i_0_1_211 (.A1(n_0_1_66), .A2(firstInputComplement[3]), .B1(n_0_1_68), 
      .B2(inputOne[3]), .ZN(n_0_1_76));
   AOI22_X1 i_0_1_212 (.A1(n_0_1_70), .A2(inputOne[2]), .B1(
      firstInputComplement[2]), .B2(n_0_1_62), .ZN(n_0_1_77));
   NAND2_X1 i_0_1_213 (.A1(n_0_1_76), .A2(n_0_1_77), .ZN(n_0_1_78));
   INV_X1 i_0_1_214 (.A(n_0_1_78), .ZN(n_0_1_79));
   OAI22_X1 i_0_1_215 (.A1(n_0_1_69), .A2(n_0_1_75), .B1(n_0_1_79), .B2(n_0_1_13), 
      .ZN(n_0_55));
   AOI22_X1 i_0_1_216 (.A1(n_0_1_66), .A2(firstInputComplement[4]), .B1(n_0_1_68), 
      .B2(inputOne[4]), .ZN(n_0_1_80));
   AOI22_X1 i_0_1_217 (.A1(n_0_1_70), .A2(inputOne[3]), .B1(
      firstInputComplement[3]), .B2(n_0_1_62), .ZN(n_0_1_81));
   NAND2_X1 i_0_1_218 (.A1(n_0_1_80), .A2(n_0_1_81), .ZN(n_0_1_82));
   INV_X1 i_0_1_219 (.A(n_0_1_54), .ZN(n_0_1_83));
   NOR2_X1 i_0_1_220 (.A1(n_0_1_10), .A2(n_0_1_15), .ZN(n_0_1_84));
   AOI22_X1 i_0_1_221 (.A1(n_0_1_82), .A2(n_0_1_11), .B1(n_0_1_83), .B2(n_0_1_84), 
      .ZN(n_0_1_85));
   OAI22_X1 i_0_1_222 (.A1(n_0_1_85), .A2(counter[0]), .B1(n_0_1_74), .B2(
      n_0_1_75), .ZN(n_0_56));
   INV_X1 i_0_1_223 (.A(n_0_1_69), .ZN(n_0_1_86));
   AOI22_X1 i_0_1_224 (.A1(n_0_1_66), .A2(firstInputComplement[5]), .B1(n_0_1_70), 
      .B2(inputOne[4]), .ZN(n_0_1_87));
   AOI22_X1 i_0_1_225 (.A1(n_0_1_68), .A2(inputOne[5]), .B1(
      firstInputComplement[4]), .B2(n_0_1_62), .ZN(n_0_1_88));
   NAND2_X1 i_0_1_226 (.A1(n_0_1_87), .A2(n_0_1_88), .ZN(n_0_1_89));
   AOI22_X1 i_0_1_227 (.A1(n_0_1_86), .A2(n_0_1_84), .B1(n_0_1_11), .B2(n_0_1_89), 
      .ZN(n_0_1_90));
   OAI22_X1 i_0_1_228 (.A1(n_0_1_90), .A2(counter[0]), .B1(n_0_1_79), .B2(
      n_0_1_75), .ZN(n_0_57));
   AOI22_X1 i_0_1_229 (.A1(n_0_1_68), .A2(inputOne[6]), .B1(n_0_1_70), .B2(
      inputOne[5]), .ZN(n_0_1_91));
   AOI22_X1 i_0_1_230 (.A1(n_0_1_66), .A2(firstInputComplement[6]), .B1(
      firstInputComplement[5]), .B2(n_0_1_62), .ZN(n_0_1_92));
   NAND2_X1 i_0_1_231 (.A1(n_0_1_91), .A2(n_0_1_92), .ZN(n_0_1_93));
   AOI22_X1 i_0_1_232 (.A1(n_0_1_93), .A2(n_0_1_11), .B1(n_0_1_73), .B2(n_0_1_84), 
      .ZN(n_0_1_94));
   OAI22_X1 i_0_1_233 (.A1(n_0_1_94), .A2(counter[0]), .B1(n_0_1_85), .B2(
      n_0_1_12), .ZN(n_0_58));
   AOI22_X1 i_0_1_234 (.A1(n_0_1_68), .A2(inputOne[7]), .B1(n_0_1_70), .B2(
      inputOne[6]), .ZN(n_0_1_95));
   AOI22_X1 i_0_1_235 (.A1(n_0_1_66), .A2(firstInputComplement[7]), .B1(
      firstInputComplement[6]), .B2(n_0_1_62), .ZN(n_0_1_96));
   NAND2_X1 i_0_1_236 (.A1(n_0_1_95), .A2(n_0_1_96), .ZN(n_0_1_97));
   AOI22_X1 i_0_1_237 (.A1(n_0_1_78), .A2(n_0_1_84), .B1(n_0_1_97), .B2(n_0_1_11), 
      .ZN(n_0_1_98));
   OAI22_X1 i_0_1_238 (.A1(n_0_1_90), .A2(n_0_1_12), .B1(n_0_1_98), .B2(
      counter[0]), .ZN(n_0_59));
   AOI22_X1 i_0_1_239 (.A1(n_0_1_68), .A2(inputOne[8]), .B1(n_0_1_70), .B2(
      inputOne[7]), .ZN(n_0_1_99));
   AOI22_X1 i_0_1_240 (.A1(n_0_1_66), .A2(firstInputComplement[8]), .B1(
      firstInputComplement[7]), .B2(n_0_1_62), .ZN(n_0_1_100));
   NAND2_X1 i_0_1_241 (.A1(n_0_1_99), .A2(n_0_1_100), .ZN(n_0_1_101));
   INV_X1 i_0_1_242 (.A(n_0_1_101), .ZN(n_0_1_102));
   NAND2_X1 i_0_1_243 (.A1(n_0_1_8), .A2(counter[2]), .ZN(n_0_1_103));
   OR2_X1 i_0_1_244 (.A1(n_0_1_103), .A2(counter[3]), .ZN(n_0_1_104));
   OAI22_X1 i_0_1_245 (.A1(n_0_1_102), .A2(n_0_1_10), .B1(n_0_1_54), .B2(
      n_0_1_104), .ZN(n_0_1_105));
   AOI22_X1 i_0_1_246 (.A1(n_0_1_105), .A2(n_0_1_15), .B1(n_0_1_82), .B2(
      n_0_1_84), .ZN(n_0_1_106));
   OAI22_X1 i_0_1_247 (.A1(n_0_1_106), .A2(counter[0]), .B1(n_0_1_12), .B2(
      n_0_1_94), .ZN(n_0_60));
   AOI22_X1 i_0_1_248 (.A1(n_0_1_66), .A2(firstInputComplement[9]), .B1(n_0_1_70), 
      .B2(inputOne[8]), .ZN(n_0_1_107));
   AOI22_X1 i_0_1_249 (.A1(n_0_1_68), .A2(inputOne[9]), .B1(
      firstInputComplement[8]), .B2(n_0_1_62), .ZN(n_0_1_108));
   NAND2_X1 i_0_1_250 (.A1(n_0_1_107), .A2(n_0_1_108), .ZN(n_0_1_109));
   INV_X1 i_0_1_251 (.A(n_0_1_109), .ZN(n_0_1_110));
   OAI22_X1 i_0_1_252 (.A1(n_0_1_69), .A2(n_0_1_104), .B1(n_0_1_110), .B2(
      n_0_1_10), .ZN(n_0_1_111));
   AOI22_X1 i_0_1_253 (.A1(n_0_1_111), .A2(n_0_1_15), .B1(n_0_1_89), .B2(
      n_0_1_84), .ZN(n_0_1_112));
   OAI22_X1 i_0_1_254 (.A1(n_0_1_112), .A2(counter[0]), .B1(n_0_1_12), .B2(
      n_0_1_98), .ZN(n_0_61));
   AOI22_X1 i_0_1_255 (.A1(n_0_1_68), .A2(inputOne[10]), .B1(n_0_1_70), .B2(
      inputOne[9]), .ZN(n_0_1_113));
   AOI22_X1 i_0_1_256 (.A1(n_0_1_66), .A2(firstInputComplement[10]), .B1(
      firstInputComplement[9]), .B2(n_0_1_62), .ZN(n_0_1_114));
   NAND2_X1 i_0_1_257 (.A1(n_0_1_113), .A2(n_0_1_114), .ZN(n_0_1_115));
   INV_X1 i_0_1_258 (.A(n_0_1_115), .ZN(n_0_1_116));
   OAI22_X1 i_0_1_259 (.A1(n_0_1_116), .A2(n_0_1_10), .B1(n_0_1_74), .B2(
      n_0_1_104), .ZN(n_0_1_117));
   AOI22_X1 i_0_1_260 (.A1(n_0_1_117), .A2(n_0_1_15), .B1(n_0_1_93), .B2(
      n_0_1_84), .ZN(n_0_1_118));
   OAI22_X1 i_0_1_261 (.A1(n_0_1_118), .A2(counter[0]), .B1(n_0_1_106), .B2(
      n_0_1_12), .ZN(n_0_62));
   AOI22_X1 i_0_1_262 (.A1(n_0_1_68), .A2(inputOne[11]), .B1(n_0_1_70), .B2(
      inputOne[10]), .ZN(n_0_1_119));
   AOI22_X1 i_0_1_263 (.A1(n_0_1_66), .A2(firstInputComplement[11]), .B1(
      firstInputComplement[10]), .B2(n_0_1_62), .ZN(n_0_1_120));
   NAND2_X1 i_0_1_264 (.A1(n_0_1_119), .A2(n_0_1_120), .ZN(n_0_1_121));
   INV_X1 i_0_1_265 (.A(n_0_1_121), .ZN(n_0_1_122));
   OAI22_X1 i_0_1_266 (.A1(n_0_1_79), .A2(n_0_1_104), .B1(n_0_1_122), .B2(
      n_0_1_10), .ZN(n_0_1_123));
   AOI22_X1 i_0_1_267 (.A1(n_0_1_123), .A2(n_0_1_15), .B1(n_0_1_97), .B2(
      n_0_1_84), .ZN(n_0_1_124));
   OAI22_X1 i_0_1_268 (.A1(n_0_1_112), .A2(n_0_1_12), .B1(n_0_1_124), .B2(
      counter[0]), .ZN(n_0_63));
   INV_X1 i_0_1_269 (.A(n_0_1_82), .ZN(n_0_1_125));
   AOI22_X1 i_0_1_270 (.A1(n_0_1_68), .A2(inputOne[12]), .B1(n_0_1_70), .B2(
      inputOne[11]), .ZN(n_0_1_126));
   AOI22_X1 i_0_1_271 (.A1(n_0_1_66), .A2(firstInputComplement[12]), .B1(
      firstInputComplement[11]), .B2(n_0_1_62), .ZN(n_0_1_127));
   NAND2_X1 i_0_1_272 (.A1(n_0_1_126), .A2(n_0_1_127), .ZN(n_0_1_128));
   INV_X1 i_0_1_273 (.A(n_0_1_128), .ZN(n_0_1_129));
   OAI22_X1 i_0_1_274 (.A1(n_0_1_125), .A2(n_0_1_104), .B1(n_0_1_129), .B2(
      n_0_1_10), .ZN(n_0_1_130));
   AOI22_X1 i_0_1_275 (.A1(n_0_1_130), .A2(n_0_1_15), .B1(n_0_1_105), .B2(
      counter[1]), .ZN(n_0_1_131));
   OAI22_X1 i_0_1_276 (.A1(n_0_1_131), .A2(counter[0]), .B1(n_0_1_118), .B2(
      n_0_1_12), .ZN(n_0_64));
   INV_X1 i_0_1_277 (.A(n_0_1_89), .ZN(n_0_1_132));
   AOI22_X1 i_0_1_278 (.A1(n_0_1_66), .A2(firstInputComplement[13]), .B1(
      n_0_1_70), .B2(inputOne[12]), .ZN(n_0_1_133));
   AOI22_X1 i_0_1_279 (.A1(n_0_1_68), .A2(inputOne[13]), .B1(
      firstInputComplement[12]), .B2(n_0_1_62), .ZN(n_0_1_134));
   NAND2_X1 i_0_1_280 (.A1(n_0_1_133), .A2(n_0_1_134), .ZN(n_0_1_135));
   INV_X1 i_0_1_281 (.A(n_0_1_135), .ZN(n_0_1_136));
   OAI22_X1 i_0_1_282 (.A1(n_0_1_132), .A2(n_0_1_104), .B1(n_0_1_136), .B2(
      n_0_1_10), .ZN(n_0_1_137));
   AOI22_X1 i_0_1_283 (.A1(n_0_1_111), .A2(counter[1]), .B1(n_0_1_137), .B2(
      n_0_1_15), .ZN(n_0_1_138));
   OAI22_X1 i_0_1_284 (.A1(n_0_1_138), .A2(counter[0]), .B1(n_0_1_124), .B2(
      n_0_1_12), .ZN(n_0_65));
   AOI22_X1 i_0_1_285 (.A1(n_0_1_68), .A2(inputOne[14]), .B1(n_0_1_70), .B2(
      inputOne[13]), .ZN(n_0_1_139));
   AOI22_X1 i_0_1_286 (.A1(n_0_1_66), .A2(firstInputComplement[14]), .B1(
      firstInputComplement[13]), .B2(n_0_1_62), .ZN(n_0_1_140));
   NAND2_X1 i_0_1_287 (.A1(n_0_1_139), .A2(n_0_1_140), .ZN(n_0_1_141));
   INV_X1 i_0_1_288 (.A(n_0_1_141), .ZN(n_0_1_142));
   INV_X1 i_0_1_289 (.A(n_0_1_93), .ZN(n_0_1_143));
   OAI22_X1 i_0_1_290 (.A1(n_0_1_142), .A2(n_0_1_10), .B1(n_0_1_143), .B2(
      n_0_1_104), .ZN(n_0_1_144));
   AOI22_X1 i_0_1_291 (.A1(n_0_1_144), .A2(n_0_1_15), .B1(n_0_1_117), .B2(
      counter[1]), .ZN(n_0_1_145));
   OAI22_X1 i_0_1_292 (.A1(n_0_1_145), .A2(counter[0]), .B1(n_0_1_131), .B2(
      n_0_1_12), .ZN(n_0_66));
   INV_X1 i_0_1_293 (.A(n_0_1_97), .ZN(n_0_1_146));
   AOI22_X1 i_0_1_294 (.A1(n_0_1_66), .A2(firstInputComplement[15]), .B1(
      n_0_1_70), .B2(inputOne[14]), .ZN(n_0_1_147));
   AOI22_X1 i_0_1_295 (.A1(n_0_1_68), .A2(inputOne[15]), .B1(n_0_1_62), .B2(
      firstInputComplement[14]), .ZN(n_0_1_148));
   NAND2_X1 i_0_1_296 (.A1(n_0_1_147), .A2(n_0_1_148), .ZN(n_0_1_149));
   INV_X1 i_0_1_297 (.A(n_0_1_149), .ZN(n_0_1_150));
   OAI22_X1 i_0_1_298 (.A1(n_0_1_146), .A2(n_0_1_104), .B1(n_0_1_150), .B2(
      n_0_1_10), .ZN(n_0_1_151));
   AOI22_X1 i_0_1_299 (.A1(n_0_1_151), .A2(n_0_1_15), .B1(n_0_1_123), .B2(
      counter[1]), .ZN(n_0_1_152));
   OAI22_X1 i_0_1_300 (.A1(n_0_1_138), .A2(n_0_1_12), .B1(n_0_1_152), .B2(
      counter[0]), .ZN(n_0_67));
   AOI22_X1 i_0_1_301 (.A1(n_0_1_66), .A2(firstInputComplement[16]), .B1(
      n_0_1_70), .B2(inputOne[15]), .ZN(n_0_1_153));
   AOI22_X1 i_0_1_302 (.A1(n_0_1_68), .A2(inputOne[16]), .B1(
      firstInputComplement[15]), .B2(n_0_1_62), .ZN(n_0_1_154));
   NAND2_X1 i_0_1_303 (.A1(n_0_1_153), .A2(n_0_1_154), .ZN(n_0_1_155));
   INV_X1 i_0_1_304 (.A(n_0_1_155), .ZN(n_0_1_156));
   OAI22_X1 i_0_1_305 (.A1(n_0_1_156), .A2(counter[3]), .B1(n_0_1_9), .B2(
      n_0_1_54), .ZN(n_0_1_157));
   NAND2_X1 i_0_1_306 (.A1(n_0_1_157), .A2(n_0_1_8), .ZN(n_0_1_158));
   OAI22_X1 i_0_1_307 (.A1(n_0_1_158), .A2(counter[2]), .B1(n_0_1_102), .B2(
      n_0_1_104), .ZN(n_0_1_159));
   AOI22_X1 i_0_1_308 (.A1(n_0_1_159), .A2(n_0_1_15), .B1(counter[1]), .B2(
      n_0_1_130), .ZN(n_0_1_160));
   OAI22_X1 i_0_1_309 (.A1(n_0_1_160), .A2(counter[0]), .B1(n_0_1_12), .B2(
      n_0_1_145), .ZN(n_0_68));
   AOI22_X1 i_0_1_310 (.A1(n_0_1_66), .A2(firstInputComplement[17]), .B1(
      n_0_1_70), .B2(inputOne[16]), .ZN(n_0_1_161));
   AOI22_X1 i_0_1_311 (.A1(n_0_1_68), .A2(inputOne[17]), .B1(
      firstInputComplement[16]), .B2(n_0_1_62), .ZN(n_0_1_162));
   NAND2_X1 i_0_1_312 (.A1(n_0_1_161), .A2(n_0_1_162), .ZN(n_0_1_163));
   OAI22_X1 i_0_1_313 (.A1(n_0_1_86), .A2(n_0_1_9), .B1(n_0_1_163), .B2(
      counter[3]), .ZN(n_0_1_164));
   NAND2_X1 i_0_1_314 (.A1(n_0_1_9), .A2(counter[2]), .ZN(n_0_1_165));
   OAI22_X1 i_0_1_315 (.A1(n_0_1_164), .A2(counter[2]), .B1(n_0_1_110), .B2(
      n_0_1_165), .ZN(n_0_1_166));
   NOR2_X1 i_0_1_316 (.A1(counter[4]), .A2(counter[1]), .ZN(n_0_1_167));
   AOI22_X1 i_0_1_317 (.A1(n_0_1_166), .A2(n_0_1_167), .B1(counter[1]), .B2(
      n_0_1_137), .ZN(n_0_1_168));
   OAI22_X1 i_0_1_318 (.A1(n_0_1_168), .A2(counter[0]), .B1(n_0_1_152), .B2(
      n_0_1_12), .ZN(n_0_69));
   AOI22_X1 i_0_1_319 (.A1(n_0_1_66), .A2(firstInputComplement[18]), .B1(
      n_0_1_70), .B2(inputOne[17]), .ZN(n_0_1_169));
   AOI22_X1 i_0_1_320 (.A1(n_0_1_68), .A2(inputOne[18]), .B1(
      firstInputComplement[17]), .B2(n_0_1_62), .ZN(n_0_1_170));
   NAND2_X1 i_0_1_321 (.A1(n_0_1_169), .A2(n_0_1_170), .ZN(n_0_1_171));
   INV_X1 i_0_1_322 (.A(n_0_1_171), .ZN(n_0_1_172));
   AOI22_X1 i_0_1_323 (.A1(n_0_1_172), .A2(n_0_1_9), .B1(n_0_1_74), .B2(
      counter[3]), .ZN(n_0_1_173));
   NAND2_X1 i_0_1_324 (.A1(n_0_1_173), .A2(n_0_1_8), .ZN(n_0_1_174));
   OAI22_X1 i_0_1_325 (.A1(n_0_1_174), .A2(counter[2]), .B1(n_0_1_116), .B2(
      n_0_1_104), .ZN(n_0_1_175));
   AOI22_X1 i_0_1_326 (.A1(n_0_1_175), .A2(n_0_1_15), .B1(counter[1]), .B2(
      n_0_1_144), .ZN(n_0_1_176));
   OAI22_X1 i_0_1_327 (.A1(n_0_1_176), .A2(counter[0]), .B1(n_0_1_160), .B2(
      n_0_1_12), .ZN(n_0_70));
   AOI22_X1 i_0_1_328 (.A1(n_0_1_68), .A2(inputOne[19]), .B1(n_0_1_66), .B2(
      firstInputComplement[19]), .ZN(n_0_1_177));
   AOI22_X1 i_0_1_329 (.A1(n_0_1_70), .A2(inputOne[18]), .B1(
      firstInputComplement[18]), .B2(n_0_1_62), .ZN(n_0_1_178));
   NAND2_X1 i_0_1_330 (.A1(n_0_1_177), .A2(n_0_1_178), .ZN(n_0_1_179));
   INV_X1 i_0_1_331 (.A(n_0_1_179), .ZN(n_0_1_180));
   AOI22_X1 i_0_1_332 (.A1(n_0_1_79), .A2(counter[3]), .B1(n_0_1_180), .B2(
      n_0_1_9), .ZN(n_0_1_181));
   NAND2_X1 i_0_1_333 (.A1(n_0_1_181), .A2(n_0_1_8), .ZN(n_0_1_182));
   OAI22_X1 i_0_1_334 (.A1(n_0_1_182), .A2(counter[2]), .B1(n_0_1_122), .B2(
      n_0_1_104), .ZN(n_0_1_183));
   AOI22_X1 i_0_1_335 (.A1(n_0_1_183), .A2(n_0_1_15), .B1(counter[1]), .B2(
      n_0_1_151), .ZN(n_0_1_184));
   OAI22_X1 i_0_1_336 (.A1(n_0_1_184), .A2(counter[0]), .B1(n_0_1_168), .B2(
      n_0_1_12), .ZN(n_0_71));
   AOI22_X1 i_0_1_337 (.A1(n_0_1_68), .A2(inputOne[20]), .B1(n_0_1_66), .B2(
      firstInputComplement[20]), .ZN(n_0_1_185));
   AOI22_X1 i_0_1_338 (.A1(n_0_1_70), .A2(inputOne[19]), .B1(
      firstInputComplement[19]), .B2(n_0_1_62), .ZN(n_0_1_186));
   NAND2_X1 i_0_1_339 (.A1(n_0_1_185), .A2(n_0_1_186), .ZN(n_0_1_187));
   INV_X1 i_0_1_340 (.A(n_0_1_187), .ZN(n_0_1_188));
   AOI22_X1 i_0_1_341 (.A1(n_0_1_125), .A2(counter[3]), .B1(n_0_1_188), .B2(
      n_0_1_9), .ZN(n_0_1_189));
   NAND2_X1 i_0_1_342 (.A1(n_0_1_189), .A2(n_0_1_8), .ZN(n_0_1_190));
   OAI22_X1 i_0_1_343 (.A1(n_0_1_190), .A2(counter[2]), .B1(n_0_1_104), .B2(
      n_0_1_129), .ZN(n_0_1_191));
   AOI22_X1 i_0_1_344 (.A1(n_0_1_191), .A2(n_0_1_15), .B1(n_0_1_159), .B2(
      counter[1]), .ZN(n_0_1_192));
   OAI22_X1 i_0_1_345 (.A1(n_0_1_192), .A2(counter[0]), .B1(n_0_1_176), .B2(
      n_0_1_12), .ZN(n_0_72));
   NOR2_X1 i_0_1_346 (.A1(n_0_1_15), .A2(counter[4]), .ZN(n_0_1_193));
   AOI22_X1 i_0_1_347 (.A1(n_0_1_66), .A2(firstInputComplement[21]), .B1(
      n_0_1_70), .B2(inputOne[20]), .ZN(n_0_1_194));
   AOI22_X1 i_0_1_348 (.A1(n_0_1_68), .A2(inputOne[21]), .B1(
      firstInputComplement[20]), .B2(n_0_1_62), .ZN(n_0_1_195));
   NAND2_X1 i_0_1_349 (.A1(n_0_1_194), .A2(n_0_1_195), .ZN(n_0_1_196));
   OAI22_X1 i_0_1_350 (.A1(n_0_1_196), .A2(counter[3]), .B1(n_0_1_89), .B2(
      n_0_1_9), .ZN(n_0_1_197));
   OAI22_X1 i_0_1_351 (.A1(n_0_1_197), .A2(counter[2]), .B1(n_0_1_136), .B2(
      n_0_1_165), .ZN(n_0_1_198));
   AOI22_X1 i_0_1_352 (.A1(n_0_1_166), .A2(n_0_1_193), .B1(n_0_1_167), .B2(
      n_0_1_198), .ZN(n_0_1_199));
   OAI22_X1 i_0_1_353 (.A1(n_0_1_184), .A2(n_0_1_12), .B1(n_0_1_199), .B2(
      counter[0]), .ZN(n_0_73));
   AOI22_X1 i_0_1_354 (.A1(n_0_1_66), .A2(firstInputComplement[22]), .B1(
      n_0_1_70), .B2(inputOne[21]), .ZN(n_0_1_200));
   AOI22_X1 i_0_1_355 (.A1(n_0_1_68), .A2(inputOne[22]), .B1(
      firstInputComplement[21]), .B2(n_0_1_62), .ZN(n_0_1_201));
   NAND2_X1 i_0_1_356 (.A1(n_0_1_200), .A2(n_0_1_201), .ZN(n_0_1_202));
   OAI22_X1 i_0_1_357 (.A1(n_0_1_202), .A2(counter[3]), .B1(n_0_1_93), .B2(
      n_0_1_9), .ZN(n_0_1_203));
   OAI22_X1 i_0_1_358 (.A1(n_0_1_203), .A2(counter[2]), .B1(n_0_1_142), .B2(
      n_0_1_165), .ZN(n_0_1_204));
   AOI22_X1 i_0_1_359 (.A1(n_0_1_175), .A2(counter[1]), .B1(n_0_1_204), .B2(
      n_0_1_167), .ZN(n_0_1_205));
   OAI22_X1 i_0_1_360 (.A1(n_0_1_192), .A2(n_0_1_12), .B1(n_0_1_205), .B2(
      counter[0]), .ZN(n_0_74));
   AOI22_X1 i_0_1_361 (.A1(n_0_1_66), .A2(firstInputComplement[23]), .B1(
      n_0_1_70), .B2(inputOne[22]), .ZN(n_0_1_206));
   AOI22_X1 i_0_1_362 (.A1(n_0_1_68), .A2(inputOne[23]), .B1(
      firstInputComplement[22]), .B2(n_0_1_62), .ZN(n_0_1_207));
   NAND2_X1 i_0_1_363 (.A1(n_0_1_206), .A2(n_0_1_207), .ZN(n_0_1_208));
   OAI22_X1 i_0_1_364 (.A1(n_0_1_208), .A2(counter[3]), .B1(n_0_1_97), .B2(
      n_0_1_9), .ZN(n_0_1_209));
   OAI22_X1 i_0_1_365 (.A1(n_0_1_209), .A2(counter[2]), .B1(n_0_1_150), .B2(
      n_0_1_165), .ZN(n_0_1_210));
   AOI22_X1 i_0_1_366 (.A1(n_0_1_183), .A2(counter[1]), .B1(n_0_1_210), .B2(
      n_0_1_167), .ZN(n_0_1_211));
   OAI22_X1 i_0_1_367 (.A1(n_0_1_211), .A2(counter[0]), .B1(n_0_1_199), .B2(
      n_0_1_12), .ZN(n_0_75));
   AOI22_X1 i_0_1_368 (.A1(n_0_1_68), .A2(inputOne[24]), .B1(n_0_1_70), .B2(
      inputOne[23]), .ZN(n_0_1_212));
   AOI22_X1 i_0_1_369 (.A1(n_0_1_66), .A2(firstInputComplement[24]), .B1(
      firstInputComplement[23]), .B2(n_0_1_62), .ZN(n_0_1_213));
   NAND2_X1 i_0_1_370 (.A1(n_0_1_212), .A2(n_0_1_213), .ZN(n_0_1_214));
   INV_X1 i_0_1_371 (.A(n_0_1_214), .ZN(n_0_1_215));
   AOI22_X1 i_0_1_372 (.A1(n_0_1_102), .A2(counter[3]), .B1(n_0_1_215), .B2(
      n_0_1_9), .ZN(n_0_1_216));
   NAND2_X1 i_0_1_373 (.A1(n_0_1_216), .A2(n_0_1_8), .ZN(n_0_1_217));
   OAI22_X1 i_0_1_374 (.A1(n_0_1_217), .A2(counter[2]), .B1(n_0_1_158), .B2(
      n_0_1_7), .ZN(n_0_1_218));
   AOI22_X1 i_0_1_375 (.A1(n_0_1_191), .A2(counter[1]), .B1(n_0_1_218), .B2(
      n_0_1_15), .ZN(n_0_1_219));
   OAI22_X1 i_0_1_376 (.A1(n_0_1_219), .A2(counter[0]), .B1(n_0_1_205), .B2(
      n_0_1_12), .ZN(n_0_76));
   AOI22_X1 i_0_1_377 (.A1(n_0_1_68), .A2(inputOne[25]), .B1(n_0_1_70), .B2(
      inputOne[24]), .ZN(n_0_1_220));
   AOI22_X1 i_0_1_378 (.A1(n_0_1_66), .A2(firstInputComplement[25]), .B1(
      firstInputComplement[24]), .B2(n_0_1_62), .ZN(n_0_1_221));
   NAND2_X1 i_0_1_379 (.A1(n_0_1_220), .A2(n_0_1_221), .ZN(n_0_1_222));
   INV_X1 i_0_1_380 (.A(n_0_1_222), .ZN(n_0_1_223));
   AOI22_X1 i_0_1_381 (.A1(n_0_1_110), .A2(counter[3]), .B1(n_0_1_223), .B2(
      n_0_1_9), .ZN(n_0_1_224));
   NAND2_X1 i_0_1_382 (.A1(n_0_1_224), .A2(n_0_1_8), .ZN(n_0_1_225));
   OAI22_X1 i_0_1_383 (.A1(n_0_1_225), .A2(counter[2]), .B1(n_0_1_164), .B2(
      n_0_1_103), .ZN(n_0_1_226));
   AOI22_X1 i_0_1_384 (.A1(n_0_1_226), .A2(n_0_1_15), .B1(n_0_1_193), .B2(
      n_0_1_198), .ZN(n_0_1_227));
   OAI22_X1 i_0_1_385 (.A1(n_0_1_227), .A2(counter[0]), .B1(n_0_1_211), .B2(
      n_0_1_12), .ZN(n_0_77));
   AOI22_X1 i_0_1_386 (.A1(n_0_1_66), .A2(firstInputComplement[26]), .B1(
      n_0_1_70), .B2(inputOne[25]), .ZN(n_0_1_228));
   AOI22_X1 i_0_1_387 (.A1(n_0_1_68), .A2(inputOne[26]), .B1(
      firstInputComplement[25]), .B2(n_0_1_62), .ZN(n_0_1_229));
   NAND2_X1 i_0_1_388 (.A1(n_0_1_228), .A2(n_0_1_229), .ZN(n_0_1_230));
   INV_X1 i_0_1_389 (.A(n_0_1_230), .ZN(n_0_1_231));
   AOI22_X1 i_0_1_390 (.A1(n_0_1_116), .A2(counter[3]), .B1(n_0_1_231), .B2(
      n_0_1_9), .ZN(n_0_1_232));
   NAND2_X1 i_0_1_391 (.A1(n_0_1_232), .A2(n_0_1_8), .ZN(n_0_1_233));
   AOI22_X1 i_0_1_392 (.A1(n_0_1_174), .A2(counter[2]), .B1(n_0_1_233), .B2(
      n_0_1_7), .ZN(n_0_1_234));
   AOI22_X1 i_0_1_393 (.A1(n_0_1_234), .A2(n_0_1_15), .B1(n_0_1_204), .B2(
      n_0_1_193), .ZN(n_0_1_235));
   OAI22_X1 i_0_1_394 (.A1(n_0_1_235), .A2(counter[0]), .B1(n_0_1_219), .B2(
      n_0_1_12), .ZN(n_0_78));
   AOI22_X1 i_0_1_395 (.A1(n_0_1_66), .A2(firstInputComplement[27]), .B1(
      n_0_1_70), .B2(inputOne[26]), .ZN(n_0_1_236));
   AOI22_X1 i_0_1_396 (.A1(n_0_1_68), .A2(inputOne[27]), .B1(
      firstInputComplement[26]), .B2(n_0_1_62), .ZN(n_0_1_237));
   NAND2_X1 i_0_1_397 (.A1(n_0_1_236), .A2(n_0_1_237), .ZN(n_0_1_238));
   INV_X1 i_0_1_398 (.A(n_0_1_238), .ZN(n_0_1_239));
   AOI22_X1 i_0_1_399 (.A1(n_0_1_122), .A2(counter[3]), .B1(n_0_1_239), .B2(
      n_0_1_9), .ZN(n_0_1_240));
   NAND2_X1 i_0_1_400 (.A1(n_0_1_240), .A2(n_0_1_8), .ZN(n_0_1_241));
   AOI22_X1 i_0_1_401 (.A1(n_0_1_182), .A2(counter[2]), .B1(n_0_1_241), .B2(
      n_0_1_7), .ZN(n_0_1_242));
   AOI22_X1 i_0_1_402 (.A1(n_0_1_242), .A2(n_0_1_15), .B1(n_0_1_210), .B2(
      n_0_1_193), .ZN(n_0_1_243));
   OAI22_X1 i_0_1_403 (.A1(n_0_1_243), .A2(counter[0]), .B1(n_0_1_227), .B2(
      n_0_1_12), .ZN(n_0_79));
   AOI22_X1 i_0_1_404 (.A1(n_0_1_66), .A2(firstInputComplement[28]), .B1(
      n_0_1_70), .B2(inputOne[27]), .ZN(n_0_1_244));
   AOI22_X1 i_0_1_405 (.A1(n_0_1_68), .A2(inputOne[28]), .B1(
      firstInputComplement[27]), .B2(n_0_1_62), .ZN(n_0_1_245));
   NAND2_X1 i_0_1_406 (.A1(n_0_1_244), .A2(n_0_1_245), .ZN(n_0_1_246));
   INV_X1 i_0_1_407 (.A(n_0_1_246), .ZN(n_0_1_247));
   AOI22_X1 i_0_1_408 (.A1(n_0_1_129), .A2(counter[3]), .B1(n_0_1_247), .B2(
      n_0_1_9), .ZN(n_0_1_248));
   NAND2_X1 i_0_1_409 (.A1(n_0_1_248), .A2(n_0_1_8), .ZN(n_0_1_249));
   OAI22_X1 i_0_1_410 (.A1(n_0_1_190), .A2(n_0_1_7), .B1(n_0_1_249), .B2(
      counter[2]), .ZN(n_0_1_250));
   AOI22_X1 i_0_1_411 (.A1(n_0_1_250), .A2(n_0_1_15), .B1(n_0_1_218), .B2(
      counter[1]), .ZN(n_0_1_251));
   OAI22_X1 i_0_1_412 (.A1(n_0_1_235), .A2(n_0_1_12), .B1(n_0_1_251), .B2(
      counter[0]), .ZN(n_0_80));
   AOI22_X1 i_0_1_413 (.A1(n_0_1_66), .A2(firstInputComplement[29]), .B1(
      n_0_1_70), .B2(inputOne[28]), .ZN(n_0_1_252));
   AOI22_X1 i_0_1_414 (.A1(n_0_1_68), .A2(inputOne[29]), .B1(
      firstInputComplement[28]), .B2(n_0_1_62), .ZN(n_0_1_253));
   NAND2_X1 i_0_1_415 (.A1(n_0_1_252), .A2(n_0_1_253), .ZN(n_0_1_254));
   INV_X1 i_0_1_416 (.A(n_0_1_254), .ZN(n_0_1_255));
   OAI22_X1 i_0_1_417 (.A1(n_0_1_255), .A2(counter[3]), .B1(n_0_1_136), .B2(
      n_0_1_9), .ZN(n_0_1_256));
   NAND2_X1 i_0_1_418 (.A1(n_0_1_256), .A2(n_0_1_8), .ZN(n_0_1_257));
   OAI22_X1 i_0_1_419 (.A1(n_0_1_257), .A2(counter[2]), .B1(n_0_1_197), .B2(
      n_0_1_103), .ZN(n_0_1_258));
   AOI22_X1 i_0_1_420 (.A1(n_0_1_226), .A2(counter[1]), .B1(n_0_1_258), .B2(
      n_0_1_15), .ZN(n_0_1_259));
   OAI22_X1 i_0_1_421 (.A1(n_0_1_243), .A2(n_0_1_12), .B1(n_0_1_259), .B2(
      counter[0]), .ZN(n_0_81));
   AOI22_X1 i_0_1_422 (.A1(n_0_1_68), .A2(inputOne[30]), .B1(n_0_1_70), .B2(
      inputOne[29]), .ZN(n_0_1_260));
   AOI22_X1 i_0_1_423 (.A1(n_0_1_66), .A2(firstInputComplement[30]), .B1(
      firstInputComplement[29]), .B2(n_0_1_62), .ZN(n_0_1_261));
   NAND2_X1 i_0_1_424 (.A1(n_0_1_260), .A2(n_0_1_261), .ZN(n_0_1_262));
   INV_X1 i_0_1_425 (.A(n_0_1_262), .ZN(n_0_1_263));
   AOI22_X1 i_0_1_426 (.A1(n_0_1_263), .A2(n_0_1_9), .B1(n_0_1_142), .B2(
      counter[3]), .ZN(n_0_1_264));
   NAND2_X1 i_0_1_427 (.A1(n_0_1_264), .A2(n_0_1_8), .ZN(n_0_1_265));
   OAI22_X1 i_0_1_428 (.A1(n_0_1_265), .A2(counter[2]), .B1(n_0_1_203), .B2(
      n_0_1_103), .ZN(n_0_1_266));
   AOI22_X1 i_0_1_429 (.A1(n_0_1_234), .A2(counter[1]), .B1(n_0_1_266), .B2(
      n_0_1_15), .ZN(n_0_1_267));
   OAI22_X1 i_0_1_430 (.A1(n_0_1_267), .A2(counter[0]), .B1(n_0_1_251), .B2(
      n_0_1_12), .ZN(n_0_82));
   AOI22_X1 i_0_1_431 (.A1(n_0_1_68), .A2(inputOne[31]), .B1(n_0_1_70), .B2(
      inputOne[30]), .ZN(n_0_1_268));
   AOI22_X1 i_0_1_432 (.A1(n_0_1_66), .A2(firstInputComplement[31]), .B1(
      firstInputComplement[30]), .B2(n_0_1_62), .ZN(n_0_1_269));
   NAND2_X1 i_0_1_433 (.A1(n_0_1_268), .A2(n_0_1_269), .ZN(n_0_1_270));
   AND2_X1 i_0_1_434 (.A1(n_0_1_270), .A2(n_0_1_8), .ZN(n_0_1_271));
   AND2_X1 i_0_1_435 (.A1(n_0_1_271), .A2(n_0_1_9), .ZN(n_0_1_272));
   NOR2_X1 i_0_1_436 (.A1(n_0_1_9), .A2(counter[4]), .ZN(n_0_1_273));
   AOI21_X1 i_0_1_437 (.A(n_0_1_272), .B1(n_0_1_149), .B2(n_0_1_273), .ZN(
      n_0_1_274));
   OAI22_X1 i_0_1_438 (.A1(n_0_1_274), .A2(counter[2]), .B1(n_0_1_103), .B2(
      n_0_1_209), .ZN(n_0_1_275));
   AOI22_X1 i_0_1_439 (.A1(n_0_1_275), .A2(n_0_1_15), .B1(n_0_1_242), .B2(
      counter[1]), .ZN(n_0_1_276));
   OAI22_X1 i_0_1_440 (.A1(n_0_1_276), .A2(counter[0]), .B1(n_0_1_259), .B2(
      n_0_1_12), .ZN(n_0_83));
   AOI221_X1 i_0_1_441 (.A(n_0_1_272), .B1(n_0_1_14), .B2(n_0_1_83), .C1(
      n_0_1_155), .C2(n_0_1_273), .ZN(n_0_1_277));
   OAI22_X1 i_0_1_442 (.A1(n_0_1_277), .A2(counter[2]), .B1(n_0_1_217), .B2(
      n_0_1_7), .ZN(n_0_1_278));
   AOI22_X1 i_0_1_443 (.A1(n_0_1_278), .A2(n_0_1_15), .B1(n_0_1_250), .B2(
      counter[1]), .ZN(n_0_1_279));
   OAI22_X1 i_0_1_444 (.A1(n_0_1_279), .A2(counter[0]), .B1(n_0_1_267), .B2(
      n_0_1_12), .ZN(n_0_84));
   AOI221_X1 i_0_1_445 (.A(n_0_1_272), .B1(n_0_1_163), .B2(n_0_1_273), .C1(
      n_0_1_86), .C2(n_0_1_14), .ZN(n_0_1_280));
   OAI22_X1 i_0_1_446 (.A1(n_0_1_280), .A2(counter[2]), .B1(n_0_1_225), .B2(
      n_0_1_7), .ZN(n_0_1_281));
   AOI22_X1 i_0_1_447 (.A1(n_0_1_281), .A2(n_0_1_15), .B1(counter[1]), .B2(
      n_0_1_258), .ZN(n_0_1_282));
   OAI22_X1 i_0_1_448 (.A1(n_0_1_282), .A2(counter[0]), .B1(n_0_1_276), .B2(
      n_0_1_12), .ZN(n_0_85));
   AOI221_X1 i_0_1_449 (.A(n_0_1_272), .B1(n_0_1_171), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_73), .ZN(n_0_1_283));
   OAI22_X1 i_0_1_450 (.A1(n_0_1_283), .A2(counter[2]), .B1(n_0_1_233), .B2(
      n_0_1_7), .ZN(n_0_1_284));
   AOI22_X1 i_0_1_451 (.A1(n_0_1_284), .A2(n_0_1_15), .B1(counter[1]), .B2(
      n_0_1_266), .ZN(n_0_1_285));
   OAI22_X1 i_0_1_452 (.A1(n_0_1_279), .A2(n_0_1_12), .B1(n_0_1_285), .B2(
      counter[0]), .ZN(n_0_86));
   AOI221_X1 i_0_1_453 (.A(n_0_1_272), .B1(n_0_1_179), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_78), .ZN(n_0_1_286));
   OAI22_X1 i_0_1_454 (.A1(n_0_1_286), .A2(counter[2]), .B1(n_0_1_241), .B2(
      n_0_1_7), .ZN(n_0_1_287));
   AOI22_X1 i_0_1_455 (.A1(n_0_1_287), .A2(n_0_1_15), .B1(n_0_1_275), .B2(
      counter[1]), .ZN(n_0_1_288));
   OAI22_X1 i_0_1_456 (.A1(n_0_1_282), .A2(n_0_1_12), .B1(n_0_1_288), .B2(
      counter[0]), .ZN(n_0_87));
   AOI221_X1 i_0_1_457 (.A(n_0_1_272), .B1(n_0_1_187), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_82), .ZN(n_0_1_289));
   OAI22_X1 i_0_1_458 (.A1(n_0_1_289), .A2(counter[2]), .B1(n_0_1_249), .B2(
      n_0_1_7), .ZN(n_0_1_290));
   AOI22_X1 i_0_1_459 (.A1(n_0_1_278), .A2(counter[1]), .B1(n_0_1_290), .B2(
      n_0_1_15), .ZN(n_0_1_291));
   OAI22_X1 i_0_1_460 (.A1(n_0_1_291), .A2(counter[0]), .B1(n_0_1_285), .B2(
      n_0_1_12), .ZN(n_0_88));
   AOI221_X1 i_0_1_461 (.A(n_0_1_272), .B1(n_0_1_196), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_89), .ZN(n_0_1_292));
   OAI22_X1 i_0_1_462 (.A1(n_0_1_292), .A2(counter[2]), .B1(n_0_1_257), .B2(
      n_0_1_7), .ZN(n_0_1_293));
   AOI22_X1 i_0_1_463 (.A1(n_0_1_281), .A2(counter[1]), .B1(n_0_1_293), .B2(
      n_0_1_15), .ZN(n_0_1_294));
   OAI22_X1 i_0_1_464 (.A1(n_0_1_294), .A2(counter[0]), .B1(n_0_1_288), .B2(
      n_0_1_12), .ZN(n_0_89));
   AOI221_X1 i_0_1_465 (.A(n_0_1_272), .B1(n_0_1_202), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_93), .ZN(n_0_1_295));
   OAI22_X1 i_0_1_466 (.A1(n_0_1_295), .A2(counter[2]), .B1(n_0_1_265), .B2(
      n_0_1_7), .ZN(n_0_1_296));
   AOI22_X1 i_0_1_467 (.A1(n_0_1_296), .A2(n_0_1_15), .B1(n_0_1_284), .B2(
      counter[1]), .ZN(n_0_1_297));
   OAI22_X1 i_0_1_468 (.A1(n_0_1_297), .A2(counter[0]), .B1(n_0_1_291), .B2(
      n_0_1_12), .ZN(n_0_90));
   AOI221_X1 i_0_1_469 (.A(n_0_1_272), .B1(n_0_1_208), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_97), .ZN(n_0_1_298));
   OAI22_X1 i_0_1_470 (.A1(n_0_1_298), .A2(counter[2]), .B1(n_0_1_7), .B2(
      n_0_1_274), .ZN(n_0_1_299));
   AOI22_X1 i_0_1_471 (.A1(n_0_1_287), .A2(counter[1]), .B1(n_0_1_299), .B2(
      n_0_1_15), .ZN(n_0_1_300));
   OAI22_X1 i_0_1_472 (.A1(n_0_1_294), .A2(n_0_1_12), .B1(n_0_1_300), .B2(
      counter[0]), .ZN(n_0_91));
   AOI221_X1 i_0_1_473 (.A(n_0_1_272), .B1(n_0_1_214), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_101), .ZN(n_0_1_301));
   OAI22_X1 i_0_1_474 (.A1(n_0_1_277), .A2(n_0_1_7), .B1(n_0_1_301), .B2(
      counter[2]), .ZN(n_0_1_302));
   AOI22_X1 i_0_1_475 (.A1(n_0_1_302), .A2(n_0_1_15), .B1(n_0_1_290), .B2(
      counter[1]), .ZN(n_0_1_303));
   OAI22_X1 i_0_1_476 (.A1(n_0_1_303), .A2(counter[0]), .B1(n_0_1_297), .B2(
      n_0_1_12), .ZN(n_0_92));
   AOI221_X1 i_0_1_477 (.A(n_0_1_272), .B1(n_0_1_222), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_109), .ZN(n_0_1_304));
   AOI22_X1 i_0_1_478 (.A1(n_0_1_280), .A2(counter[2]), .B1(n_0_1_304), .B2(
      n_0_1_7), .ZN(n_0_1_305));
   AOI22_X1 i_0_1_479 (.A1(n_0_1_305), .A2(n_0_1_15), .B1(n_0_1_293), .B2(
      counter[1]), .ZN(n_0_1_306));
   OAI22_X1 i_0_1_480 (.A1(n_0_1_306), .A2(counter[0]), .B1(n_0_1_300), .B2(
      n_0_1_12), .ZN(n_0_93));
   AOI221_X1 i_0_1_481 (.A(n_0_1_272), .B1(n_0_1_230), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_115), .ZN(n_0_1_307));
   OAI22_X1 i_0_1_482 (.A1(n_0_1_283), .A2(n_0_1_7), .B1(n_0_1_307), .B2(
      counter[2]), .ZN(n_0_1_308));
   AOI22_X1 i_0_1_483 (.A1(n_0_1_308), .A2(n_0_1_15), .B1(n_0_1_296), .B2(
      counter[1]), .ZN(n_0_1_309));
   OAI22_X1 i_0_1_484 (.A1(n_0_1_309), .A2(counter[0]), .B1(n_0_1_303), .B2(
      n_0_1_12), .ZN(n_0_94));
   AOI221_X1 i_0_1_485 (.A(n_0_1_272), .B1(n_0_1_238), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_121), .ZN(n_0_1_310));
   OAI22_X1 i_0_1_486 (.A1(n_0_1_286), .A2(n_0_1_7), .B1(n_0_1_310), .B2(
      counter[2]), .ZN(n_0_1_311));
   AOI22_X1 i_0_1_487 (.A1(n_0_1_311), .A2(n_0_1_15), .B1(n_0_1_299), .B2(
      counter[1]), .ZN(n_0_1_312));
   OAI22_X1 i_0_1_488 (.A1(n_0_1_306), .A2(n_0_1_12), .B1(n_0_1_312), .B2(
      counter[0]), .ZN(n_0_95));
   AOI221_X1 i_0_1_489 (.A(n_0_1_272), .B1(n_0_1_246), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_128), .ZN(n_0_1_313));
   OAI22_X1 i_0_1_490 (.A1(n_0_1_289), .A2(n_0_1_7), .B1(n_0_1_313), .B2(
      counter[2]), .ZN(n_0_1_314));
   AOI22_X1 i_0_1_491 (.A1(n_0_1_302), .A2(counter[1]), .B1(n_0_1_314), .B2(
      n_0_1_15), .ZN(n_0_1_315));
   OAI22_X1 i_0_1_492 (.A1(n_0_1_315), .A2(counter[0]), .B1(n_0_1_309), .B2(
      n_0_1_12), .ZN(n_0_96));
   AOI221_X1 i_0_1_493 (.A(n_0_1_272), .B1(n_0_1_254), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_135), .ZN(n_0_1_316));
   AOI22_X1 i_0_1_494 (.A1(n_0_1_292), .A2(counter[2]), .B1(n_0_1_316), .B2(
      n_0_1_7), .ZN(n_0_1_317));
   AOI22_X1 i_0_1_495 (.A1(n_0_1_305), .A2(counter[1]), .B1(n_0_1_317), .B2(
      n_0_1_15), .ZN(n_0_1_318));
   OAI22_X1 i_0_1_496 (.A1(n_0_1_318), .A2(counter[0]), .B1(n_0_1_312), .B2(
      n_0_1_12), .ZN(n_0_97));
   AOI221_X1 i_0_1_497 (.A(n_0_1_272), .B1(n_0_1_262), .B2(n_0_1_273), .C1(
      n_0_1_14), .C2(n_0_1_141), .ZN(n_0_1_319));
   AOI22_X1 i_0_1_498 (.A1(n_0_1_295), .A2(counter[2]), .B1(n_0_1_319), .B2(
      n_0_1_7), .ZN(n_0_1_320));
   AOI22_X1 i_0_1_499 (.A1(n_0_1_320), .A2(n_0_1_15), .B1(n_0_1_308), .B2(
      counter[1]), .ZN(n_0_1_321));
   OAI22_X1 i_0_1_500 (.A1(n_0_1_321), .A2(counter[0]), .B1(n_0_1_315), .B2(
      n_0_1_12), .ZN(n_0_98));
   AOI21_X1 i_0_1_501 (.A(n_0_1_271), .B1(n_0_1_14), .B2(n_0_1_149), .ZN(
      n_0_1_322));
   AOI22_X1 i_0_1_502 (.A1(n_0_1_298), .A2(counter[2]), .B1(n_0_1_7), .B2(
      n_0_1_322), .ZN(n_0_1_323));
   AOI22_X1 i_0_1_503 (.A1(n_0_1_311), .A2(counter[1]), .B1(n_0_1_323), .B2(
      n_0_1_15), .ZN(n_0_1_324));
   OAI22_X1 i_0_1_504 (.A1(n_0_1_318), .A2(n_0_1_12), .B1(n_0_1_324), .B2(
      counter[0]), .ZN(n_0_99));
   NAND2_X1 i_0_1_505 (.A1(n_0_1_157), .A2(counter[4]), .ZN(n_0_1_325));
   NOR2_X1 i_0_1_506 (.A1(n_0_1_271), .A2(counter[2]), .ZN(n_0_1_326));
   AOI22_X1 i_0_1_507 (.A1(n_0_1_301), .A2(counter[2]), .B1(n_0_1_325), .B2(
      n_0_1_326), .ZN(n_0_1_327));
   AOI22_X1 i_0_1_508 (.A1(n_0_1_314), .A2(counter[1]), .B1(n_0_1_327), .B2(
      n_0_1_15), .ZN(n_0_1_328));
   OAI22_X1 i_0_1_509 (.A1(n_0_1_321), .A2(n_0_1_12), .B1(n_0_1_328), .B2(
      counter[0]), .ZN(n_0_100));
   OR2_X1 i_0_1_510 (.A1(n_0_1_164), .A2(n_0_1_8), .ZN(n_0_1_329));
   AOI22_X1 i_0_1_511 (.A1(n_0_1_304), .A2(counter[2]), .B1(n_0_1_329), .B2(
      n_0_1_326), .ZN(n_0_1_330));
   AOI22_X1 i_0_1_512 (.A1(n_0_1_317), .A2(counter[1]), .B1(n_0_1_330), .B2(
      n_0_1_15), .ZN(n_0_1_331));
   OAI22_X1 i_0_1_513 (.A1(n_0_1_331), .A2(counter[0]), .B1(n_0_1_324), .B2(
      n_0_1_12), .ZN(n_0_101));
   NAND2_X1 i_0_1_514 (.A1(n_0_1_173), .A2(counter[4]), .ZN(n_0_1_332));
   AOI22_X1 i_0_1_515 (.A1(n_0_1_307), .A2(counter[2]), .B1(n_0_1_332), .B2(
      n_0_1_326), .ZN(n_0_1_333));
   AOI22_X1 i_0_1_516 (.A1(n_0_1_320), .A2(counter[1]), .B1(n_0_1_333), .B2(
      n_0_1_15), .ZN(n_0_1_334));
   OAI22_X1 i_0_1_517 (.A1(n_0_1_334), .A2(counter[0]), .B1(n_0_1_328), .B2(
      n_0_1_12), .ZN(n_0_102));
   NAND2_X1 i_0_1_518 (.A1(n_0_1_181), .A2(counter[4]), .ZN(n_0_1_335));
   AOI22_X1 i_0_1_519 (.A1(n_0_1_310), .A2(counter[2]), .B1(n_0_1_335), .B2(
      n_0_1_326), .ZN(n_0_1_336));
   AOI22_X1 i_0_1_520 (.A1(n_0_1_336), .A2(n_0_1_15), .B1(n_0_1_323), .B2(
      counter[1]), .ZN(n_0_1_337));
   OAI22_X1 i_0_1_521 (.A1(n_0_1_331), .A2(n_0_1_12), .B1(n_0_1_337), .B2(
      counter[0]), .ZN(n_0_103));
   NAND2_X1 i_0_1_522 (.A1(n_0_1_189), .A2(counter[4]), .ZN(n_0_1_338));
   AOI22_X1 i_0_1_523 (.A1(n_0_1_313), .A2(counter[2]), .B1(n_0_1_338), .B2(
      n_0_1_326), .ZN(n_0_1_339));
   AOI22_X1 i_0_1_524 (.A1(n_0_1_339), .A2(n_0_1_15), .B1(n_0_1_327), .B2(
      counter[1]), .ZN(n_0_1_340));
   OAI22_X1 i_0_1_525 (.A1(n_0_1_334), .A2(n_0_1_12), .B1(n_0_1_340), .B2(
      counter[0]), .ZN(n_0_104));
   OR2_X1 i_0_1_526 (.A1(n_0_1_197), .A2(n_0_1_8), .ZN(n_0_1_341));
   AOI22_X1 i_0_1_527 (.A1(n_0_1_316), .A2(counter[2]), .B1(n_0_1_341), .B2(
      n_0_1_326), .ZN(n_0_1_342));
   AOI22_X1 i_0_1_528 (.A1(n_0_1_330), .A2(counter[1]), .B1(n_0_1_342), .B2(
      n_0_1_15), .ZN(n_0_1_343));
   OAI22_X1 i_0_1_529 (.A1(n_0_1_337), .A2(n_0_1_12), .B1(n_0_1_343), .B2(
      counter[0]), .ZN(n_0_105));
   OR2_X1 i_0_1_530 (.A1(n_0_1_203), .A2(n_0_1_8), .ZN(n_0_1_344));
   AOI22_X1 i_0_1_531 (.A1(n_0_1_319), .A2(counter[2]), .B1(n_0_1_344), .B2(
      n_0_1_326), .ZN(n_0_1_345));
   AOI22_X1 i_0_1_532 (.A1(n_0_1_345), .A2(n_0_1_15), .B1(n_0_1_333), .B2(
      counter[1]), .ZN(n_0_1_346));
   OAI22_X1 i_0_1_533 (.A1(n_0_1_340), .A2(n_0_1_12), .B1(n_0_1_346), .B2(
      counter[0]), .ZN(n_0_106));
   OR2_X1 i_0_1_534 (.A1(n_0_1_209), .A2(n_0_1_8), .ZN(n_0_1_347));
   AOI22_X1 i_0_1_535 (.A1(n_0_1_347), .A2(n_0_1_326), .B1(n_0_1_322), .B2(
      counter[2]), .ZN(n_0_1_348));
   AOI22_X1 i_0_1_536 (.A1(n_0_1_336), .A2(counter[1]), .B1(n_0_1_15), .B2(
      n_0_1_348), .ZN(n_0_1_349));
   OAI22_X1 i_0_1_537 (.A1(n_0_1_343), .A2(n_0_1_12), .B1(n_0_1_349), .B2(
      counter[0]), .ZN(n_0_107));
   NAND2_X1 i_0_1_538 (.A1(n_0_1_216), .A2(counter[4]), .ZN(n_0_1_350));
   NOR2_X1 i_0_1_539 (.A1(n_0_1_271), .A2(n_0_1_7), .ZN(n_0_1_351));
   AOI22_X1 i_0_1_540 (.A1(n_0_1_350), .A2(n_0_1_326), .B1(n_0_1_325), .B2(
      n_0_1_351), .ZN(n_0_1_352));
   AOI22_X1 i_0_1_541 (.A1(n_0_1_339), .A2(counter[1]), .B1(n_0_1_15), .B2(
      n_0_1_352), .ZN(n_0_1_353));
   OAI22_X1 i_0_1_542 (.A1(n_0_1_346), .A2(n_0_1_12), .B1(n_0_1_353), .B2(
      counter[0]), .ZN(n_0_108));
   INV_X1 i_0_1_543 (.A(n_0_1_326), .ZN(n_0_1_354));
   AOI21_X1 i_0_1_544 (.A(n_0_1_354), .B1(n_0_1_224), .B2(counter[4]), .ZN(
      n_0_1_355));
   AOI21_X1 i_0_1_545 (.A(n_0_1_355), .B1(n_0_1_329), .B2(n_0_1_351), .ZN(
      n_0_1_356));
   AOI22_X1 i_0_1_546 (.A1(n_0_1_342), .A2(counter[1]), .B1(n_0_1_356), .B2(
      n_0_1_15), .ZN(n_0_1_357));
   OAI22_X1 i_0_1_547 (.A1(n_0_1_349), .A2(n_0_1_12), .B1(n_0_1_357), .B2(
      counter[0]), .ZN(n_0_109));
   NAND2_X1 i_0_1_548 (.A1(n_0_1_232), .A2(counter[4]), .ZN(n_0_1_358));
   AOI22_X1 i_0_1_549 (.A1(n_0_1_358), .A2(n_0_1_326), .B1(n_0_1_332), .B2(
      n_0_1_351), .ZN(n_0_1_359));
   AOI22_X1 i_0_1_550 (.A1(n_0_1_345), .A2(counter[1]), .B1(n_0_1_359), .B2(
      n_0_1_15), .ZN(n_0_1_360));
   OAI22_X1 i_0_1_551 (.A1(n_0_1_353), .A2(n_0_1_12), .B1(n_0_1_360), .B2(
      counter[0]), .ZN(n_0_110));
   NAND2_X1 i_0_1_552 (.A1(n_0_1_240), .A2(counter[4]), .ZN(n_0_1_361));
   AOI22_X1 i_0_1_553 (.A1(n_0_1_335), .A2(n_0_1_351), .B1(n_0_1_361), .B2(
      n_0_1_326), .ZN(n_0_1_362));
   AOI22_X1 i_0_1_554 (.A1(n_0_1_348), .A2(counter[1]), .B1(n_0_1_362), .B2(
      n_0_1_15), .ZN(n_0_1_363));
   OAI22_X1 i_0_1_555 (.A1(n_0_1_357), .A2(n_0_1_12), .B1(n_0_1_363), .B2(
      counter[0]), .ZN(n_0_111));
   NAND2_X1 i_0_1_556 (.A1(n_0_1_248), .A2(counter[4]), .ZN(n_0_1_364));
   AOI221_X1 i_0_1_557 (.A(counter[1]), .B1(n_0_1_364), .B2(n_0_1_326), .C1(
      n_0_1_338), .C2(n_0_1_351), .ZN(n_0_1_365));
   AOI21_X1 i_0_1_558 (.A(n_0_1_365), .B1(counter[1]), .B2(n_0_1_352), .ZN(
      n_0_1_366));
   OAI22_X1 i_0_1_559 (.A1(n_0_1_366), .A2(counter[0]), .B1(n_0_1_360), .B2(
      n_0_1_12), .ZN(n_0_112));
   NAND2_X1 i_0_1_560 (.A1(n_0_1_256), .A2(counter[4]), .ZN(n_0_1_367));
   AOI221_X1 i_0_1_561 (.A(counter[1]), .B1(n_0_1_367), .B2(n_0_1_326), .C1(
      n_0_1_341), .C2(n_0_1_351), .ZN(n_0_1_368));
   AOI21_X1 i_0_1_562 (.A(n_0_1_368), .B1(counter[1]), .B2(n_0_1_356), .ZN(
      n_0_1_369));
   OAI22_X1 i_0_1_563 (.A1(n_0_1_369), .A2(counter[0]), .B1(n_0_1_12), .B2(
      n_0_1_363), .ZN(n_0_113));
   NAND2_X1 i_0_1_564 (.A1(n_0_1_264), .A2(counter[4]), .ZN(n_0_1_370));
   AOI22_X1 i_0_1_565 (.A1(n_0_1_370), .A2(n_0_1_326), .B1(n_0_1_344), .B2(
      n_0_1_351), .ZN(n_0_1_371));
   OAI221_X1 i_0_1_566 (.A(n_0_1_12), .B1(n_0_1_359), .B2(n_0_1_15), .C1(
      counter[1]), .C2(n_0_1_371), .ZN(n_0_1_372));
   OAI21_X1 i_0_1_567 (.A(n_0_1_372), .B1(n_0_1_366), .B2(n_0_1_12), .ZN(n_0_114));
   OAI21_X1 i_0_1_568 (.A(n_0_1_270), .B1(n_0_1_8), .B2(n_0_1_9), .ZN(n_0_1_373));
   NAND3_X1 i_0_1_569 (.A1(n_0_1_149), .A2(counter[4]), .A3(counter[3]), 
      .ZN(n_0_1_374));
   NAND4_X1 i_0_1_570 (.A1(n_0_1_373), .A2(n_0_1_374), .A3(n_0_1_7), .A4(
      n_0_1_15), .ZN(n_0_1_375));
   NAND2_X1 i_0_1_571 (.A1(n_0_1_347), .A2(n_0_1_351), .ZN(n_0_1_376));
   OAI221_X1 i_0_1_572 (.A(n_0_1_375), .B1(n_0_1_376), .B2(counter[1]), .C1(
      n_0_1_362), .C2(n_0_1_15), .ZN(n_0_1_377));
   OAI22_X1 i_0_1_573 (.A1(n_0_1_369), .A2(n_0_1_12), .B1(n_0_1_377), .B2(
      counter[0]), .ZN(n_0_115));
   CLKGATETST_X1 clk_gate_counter_reg (.CK(clk), .E(enable), .SE(1'b0), .GCK(
      n_0_0));
   DFF_X1 \counter_reg[4]  (.D(n_0_263), .CK(n_0_0), .Q(counter[4]), .QN());
   DFF_X1 \counter_reg[3]  (.D(n_0_262), .CK(n_0_0), .Q(counter[3]), .QN());
   DFF_X1 \counter_reg[2]  (.D(n_0_261), .CK(n_0_0), .Q(counter[2]), .QN());
   DFF_X1 \counter_reg[1]  (.D(n_0_260), .CK(n_0_0), .Q(counter[1]), .QN());
   DFF_X1 \counter_reg[0]  (.D(n_0_259), .CK(n_0_0), .Q(counter[0]), .QN());
   DFF_X1 resetReg_reg (.D(n_0_264), .CK(clk), .Q(resetReg), .QN());
   MUX2_X1 resetReg_reg_enable_mux_0 (.A(resetReg), .B(n_0_129), .S(n_0_130), 
      .Z(n_0_264));
endmodule

module buffer__0_18(clk, rst, en, D, Q);
   input clk;
   input rst;
   input en;
   input [31:0]D;
   output [31:0]Q;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[31]  (.D(n_33), .CK(n_0), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_32), .CK(n_0), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_31), .CK(n_0), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_30), .CK(n_0), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_29), .CK(n_0), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_28), .CK(n_0), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_27), .CK(n_0), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_26), .CK(n_0), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_25), .CK(n_0), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_24), .CK(n_0), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_23), .CK(n_0), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_22), .CK(n_0), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_21), .CK(n_0), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_20), .CK(n_0), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_19), .CK(n_0), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_18), .CK(n_0), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_17), .CK(n_0), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_16), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_15), .CK(n_0), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_14), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_13), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_12), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_11), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_10), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_9), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_8), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_7), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_6), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_5), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_4), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_3), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_2), .CK(n_0), .Q(Q[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(rst), .ZN(n_1));
   INV_X1 i_0_1 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(D[31]), .ZN(n_33));
endmodule

module buffer(clk, rst, en, D, Q);
   input clk;
   input rst;
   input en;
   input [31:0]D;
   output [31:0]Q;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[31]  (.D(n_33), .CK(n_0), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_32), .CK(n_0), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_31), .CK(n_0), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_30), .CK(n_0), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_29), .CK(n_0), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_28), .CK(n_0), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_27), .CK(n_0), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_26), .CK(n_0), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_25), .CK(n_0), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_24), .CK(n_0), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_23), .CK(n_0), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_22), .CK(n_0), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_21), .CK(n_0), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_20), .CK(n_0), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_19), .CK(n_0), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_18), .CK(n_0), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_17), .CK(n_0), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_16), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_15), .CK(n_0), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_14), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_13), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_12), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_11), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_10), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_9), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_8), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_7), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_6), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_5), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_4), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_3), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_2), .CK(n_0), .Q(Q[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(rst), .ZN(n_1));
   INV_X1 i_0_1 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(D[31]), .ZN(n_33));
endmodule

module buffer__parameterized0(clk, rst, en, D, Q);
   input clk;
   input rst;
   input en;
   input [63:0]D;
   output [63:0]Q;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[63]  (.D(n_65), .CK(n_0), .Q(Q[63]), .QN());
   DFF_X1 \Q_reg[62]  (.D(n_64), .CK(n_0), .Q(Q[62]), .QN());
   DFF_X1 \Q_reg[61]  (.D(n_63), .CK(n_0), .Q(Q[61]), .QN());
   DFF_X1 \Q_reg[60]  (.D(n_62), .CK(n_0), .Q(Q[60]), .QN());
   DFF_X1 \Q_reg[59]  (.D(n_61), .CK(n_0), .Q(Q[59]), .QN());
   DFF_X1 \Q_reg[58]  (.D(n_60), .CK(n_0), .Q(Q[58]), .QN());
   DFF_X1 \Q_reg[57]  (.D(n_59), .CK(n_0), .Q(Q[57]), .QN());
   DFF_X1 \Q_reg[56]  (.D(n_58), .CK(n_0), .Q(Q[56]), .QN());
   DFF_X1 \Q_reg[55]  (.D(n_57), .CK(n_0), .Q(Q[55]), .QN());
   DFF_X1 \Q_reg[54]  (.D(n_56), .CK(n_0), .Q(Q[54]), .QN());
   DFF_X1 \Q_reg[53]  (.D(n_55), .CK(n_0), .Q(Q[53]), .QN());
   DFF_X1 \Q_reg[52]  (.D(n_54), .CK(n_0), .Q(Q[52]), .QN());
   DFF_X1 \Q_reg[51]  (.D(n_53), .CK(n_0), .Q(Q[51]), .QN());
   DFF_X1 \Q_reg[50]  (.D(n_52), .CK(n_0), .Q(Q[50]), .QN());
   DFF_X1 \Q_reg[49]  (.D(n_51), .CK(n_0), .Q(Q[49]), .QN());
   DFF_X1 \Q_reg[48]  (.D(n_50), .CK(n_0), .Q(Q[48]), .QN());
   DFF_X1 \Q_reg[47]  (.D(n_49), .CK(n_0), .Q(Q[47]), .QN());
   DFF_X1 \Q_reg[46]  (.D(n_48), .CK(n_0), .Q(Q[46]), .QN());
   DFF_X1 \Q_reg[45]  (.D(n_47), .CK(n_0), .Q(Q[45]), .QN());
   DFF_X1 \Q_reg[44]  (.D(n_46), .CK(n_0), .Q(Q[44]), .QN());
   DFF_X1 \Q_reg[43]  (.D(n_45), .CK(n_0), .Q(Q[43]), .QN());
   DFF_X1 \Q_reg[42]  (.D(n_44), .CK(n_0), .Q(Q[42]), .QN());
   DFF_X1 \Q_reg[41]  (.D(n_43), .CK(n_0), .Q(Q[41]), .QN());
   DFF_X1 \Q_reg[40]  (.D(n_42), .CK(n_0), .Q(Q[40]), .QN());
   DFF_X1 \Q_reg[39]  (.D(n_41), .CK(n_0), .Q(Q[39]), .QN());
   DFF_X1 \Q_reg[38]  (.D(n_40), .CK(n_0), .Q(Q[38]), .QN());
   DFF_X1 \Q_reg[37]  (.D(n_39), .CK(n_0), .Q(Q[37]), .QN());
   DFF_X1 \Q_reg[36]  (.D(n_38), .CK(n_0), .Q(Q[36]), .QN());
   DFF_X1 \Q_reg[35]  (.D(n_37), .CK(n_0), .Q(Q[35]), .QN());
   DFF_X1 \Q_reg[34]  (.D(n_36), .CK(n_0), .Q(Q[34]), .QN());
   DFF_X1 \Q_reg[33]  (.D(n_35), .CK(n_0), .Q(Q[33]), .QN());
   DFF_X1 \Q_reg[32]  (.D(n_34), .CK(n_0), .Q(Q[32]), .QN());
   DFF_X1 \Q_reg[31]  (.D(n_33), .CK(n_0), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_32), .CK(n_0), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_31), .CK(n_0), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_30), .CK(n_0), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_29), .CK(n_0), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_28), .CK(n_0), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_27), .CK(n_0), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_26), .CK(n_0), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_25), .CK(n_0), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_24), .CK(n_0), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_23), .CK(n_0), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_22), .CK(n_0), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_21), .CK(n_0), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_20), .CK(n_0), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_19), .CK(n_0), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_18), .CK(n_0), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_17), .CK(n_0), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_16), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_15), .CK(n_0), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_14), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_13), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_12), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_11), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_10), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_9), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_8), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_7), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_6), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_5), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_4), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_3), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_2), .CK(n_0), .Q(Q[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(rst), .ZN(n_1));
   INV_X1 i_0_1 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(D[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(D[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(D[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(D[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(D[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(D[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(D[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(D[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(D[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(D[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(D[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(D[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(D[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(D[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(D[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(D[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(D[31]), .ZN(n_33));
   AND2_X1 i_0_34 (.A1(n_0_0), .A2(D[32]), .ZN(n_34));
   AND2_X1 i_0_35 (.A1(n_0_0), .A2(D[33]), .ZN(n_35));
   AND2_X1 i_0_36 (.A1(n_0_0), .A2(D[34]), .ZN(n_36));
   AND2_X1 i_0_37 (.A1(n_0_0), .A2(D[35]), .ZN(n_37));
   AND2_X1 i_0_38 (.A1(n_0_0), .A2(D[36]), .ZN(n_38));
   AND2_X1 i_0_39 (.A1(n_0_0), .A2(D[37]), .ZN(n_39));
   AND2_X1 i_0_40 (.A1(n_0_0), .A2(D[38]), .ZN(n_40));
   AND2_X1 i_0_41 (.A1(n_0_0), .A2(D[39]), .ZN(n_41));
   AND2_X1 i_0_42 (.A1(n_0_0), .A2(D[40]), .ZN(n_42));
   AND2_X1 i_0_43 (.A1(n_0_0), .A2(D[41]), .ZN(n_43));
   AND2_X1 i_0_44 (.A1(n_0_0), .A2(D[42]), .ZN(n_44));
   AND2_X1 i_0_45 (.A1(n_0_0), .A2(D[43]), .ZN(n_45));
   AND2_X1 i_0_46 (.A1(n_0_0), .A2(D[44]), .ZN(n_46));
   AND2_X1 i_0_47 (.A1(n_0_0), .A2(D[45]), .ZN(n_47));
   AND2_X1 i_0_48 (.A1(n_0_0), .A2(D[46]), .ZN(n_48));
   AND2_X1 i_0_49 (.A1(n_0_0), .A2(D[47]), .ZN(n_49));
   AND2_X1 i_0_50 (.A1(n_0_0), .A2(D[48]), .ZN(n_50));
   AND2_X1 i_0_51 (.A1(n_0_0), .A2(D[49]), .ZN(n_51));
   AND2_X1 i_0_52 (.A1(n_0_0), .A2(D[50]), .ZN(n_52));
   AND2_X1 i_0_53 (.A1(n_0_0), .A2(D[51]), .ZN(n_53));
   AND2_X1 i_0_54 (.A1(n_0_0), .A2(D[52]), .ZN(n_54));
   AND2_X1 i_0_55 (.A1(n_0_0), .A2(D[53]), .ZN(n_55));
   AND2_X1 i_0_56 (.A1(n_0_0), .A2(D[54]), .ZN(n_56));
   AND2_X1 i_0_57 (.A1(n_0_0), .A2(D[55]), .ZN(n_57));
   AND2_X1 i_0_58 (.A1(n_0_0), .A2(D[56]), .ZN(n_58));
   AND2_X1 i_0_59 (.A1(n_0_0), .A2(D[57]), .ZN(n_59));
   AND2_X1 i_0_60 (.A1(n_0_0), .A2(D[58]), .ZN(n_60));
   AND2_X1 i_0_61 (.A1(n_0_0), .A2(D[59]), .ZN(n_61));
   AND2_X1 i_0_62 (.A1(n_0_0), .A2(D[60]), .ZN(n_62));
   AND2_X1 i_0_63 (.A1(n_0_0), .A2(D[61]), .ZN(n_63));
   AND2_X1 i_0_64 (.A1(n_0_0), .A2(D[62]), .ZN(n_64));
   AND2_X1 i_0_65 (.A1(n_0_0), .A2(D[63]), .ZN(n_65));
endmodule

module finalRadix4(inputA, inputB, clk, reset, en, result);
   input [31:0]inputA;
   input [31:0]inputB;
   input clk;
   input reset;
   input en;
   output [63:0]result;

   wire enableOutput;
   wire [63:0]result_out;
   wire [31:0]A_reg;
   wire [31:0]B_reg;

   RadixNoaman radixNoamanMult (.inputOne(A_reg), .inputTwo(B_reg), .finalResult(
      result_out), .clk(clk), .reset(reset), .enable(en), .enableRegisterOutput(
      enableOutput));
   buffer__0_18 regA (.clk(clk), .rst(reset), .en(en), .D(inputA), .Q(A_reg));
   buffer regB (.clk(clk), .rst(reset), .en(en), .D(inputB), .Q(B_reg));
   buffer__parameterized0 out (.clk(clk), .rst(reset), .en(enableOutput), 
      .D(result_out), .Q(result));
endmodule
