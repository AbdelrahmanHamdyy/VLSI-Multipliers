
// 	Fri Dec 23 03:07:13 2022
//	vlsi
//	localhost.localdomain

module buffer__parameterized0 (clk_CTS_0_PP_10, clk, rst, en, D, Q);

output [63:0] Q;
input [63:0] D;
input clk;
input en;
input rst;
input clk_CTS_0_PP_10;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_10;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire hfn_ipo_n5;
wire CTS_n_tid1_11;


AND2_X1 i_0_65 (.ZN (n_65), .A1 (hfn_ipo_n5), .A2 (D[63]));
AND2_X1 i_0_64 (.ZN (n_64), .A1 (hfn_ipo_n5), .A2 (D[62]));
AND2_X1 i_0_63 (.ZN (n_63), .A1 (hfn_ipo_n5), .A2 (D[61]));
AND2_X1 i_0_62 (.ZN (n_62), .A1 (hfn_ipo_n5), .A2 (D[60]));
AND2_X1 i_0_61 (.ZN (n_61), .A1 (hfn_ipo_n5), .A2 (D[59]));
AND2_X1 i_0_60 (.ZN (n_60), .A1 (hfn_ipo_n5), .A2 (D[58]));
AND2_X1 i_0_59 (.ZN (n_59), .A1 (hfn_ipo_n5), .A2 (D[57]));
AND2_X1 i_0_58 (.ZN (n_58), .A1 (hfn_ipo_n5), .A2 (D[56]));
AND2_X1 i_0_57 (.ZN (n_57), .A1 (hfn_ipo_n5), .A2 (D[55]));
AND2_X1 i_0_56 (.ZN (n_56), .A1 (n_0_0), .A2 (D[54]));
AND2_X1 i_0_55 (.ZN (n_55), .A1 (n_0_0), .A2 (D[53]));
AND2_X1 i_0_54 (.ZN (n_54), .A1 (n_0_0), .A2 (D[52]));
AND2_X1 i_0_53 (.ZN (n_53), .A1 (n_0_0), .A2 (D[51]));
AND2_X1 i_0_52 (.ZN (n_52), .A1 (n_0_0), .A2 (D[50]));
AND2_X1 i_0_51 (.ZN (n_51), .A1 (n_0_0), .A2 (D[49]));
AND2_X1 i_0_50 (.ZN (n_50), .A1 (n_0_0), .A2 (D[48]));
AND2_X1 i_0_49 (.ZN (n_49), .A1 (n_0_0), .A2 (D[47]));
AND2_X1 i_0_48 (.ZN (n_48), .A1 (n_0_0), .A2 (D[46]));
AND2_X1 i_0_47 (.ZN (n_47), .A1 (n_0_0), .A2 (D[45]));
AND2_X1 i_0_46 (.ZN (n_46), .A1 (n_0_0), .A2 (D[44]));
AND2_X1 i_0_45 (.ZN (n_45), .A1 (n_0_0), .A2 (D[43]));
AND2_X1 i_0_44 (.ZN (n_44), .A1 (n_0_0), .A2 (D[42]));
AND2_X1 i_0_43 (.ZN (n_43), .A1 (n_0_0), .A2 (D[41]));
AND2_X1 i_0_42 (.ZN (n_42), .A1 (n_0_0), .A2 (D[40]));
AND2_X1 i_0_41 (.ZN (n_41), .A1 (n_0_0), .A2 (D[39]));
AND2_X1 i_0_40 (.ZN (n_40), .A1 (n_0_0), .A2 (D[38]));
AND2_X1 i_0_39 (.ZN (n_39), .A1 (n_0_0), .A2 (D[37]));
AND2_X1 i_0_38 (.ZN (n_38), .A1 (n_0_0), .A2 (D[36]));
AND2_X1 i_0_37 (.ZN (n_37), .A1 (n_0_0), .A2 (D[35]));
AND2_X1 i_0_36 (.ZN (n_36), .A1 (n_0_0), .A2 (D[34]));
AND2_X1 i_0_35 (.ZN (n_35), .A1 (n_0_0), .A2 (D[33]));
AND2_X1 i_0_34 (.ZN (n_34), .A1 (n_0_0), .A2 (D[32]));
AND2_X1 i_0_33 (.ZN (n_33), .A1 (hfn_ipo_n5), .A2 (D[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (hfn_ipo_n5), .A2 (D[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (hfn_ipo_n5), .A2 (D[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (hfn_ipo_n5), .A2 (D[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (hfn_ipo_n5), .A2 (D[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (hfn_ipo_n5), .A2 (D[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (hfn_ipo_n5), .A2 (D[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (hfn_ipo_n5), .A2 (D[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (hfn_ipo_n5), .A2 (D[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (hfn_ipo_n5), .A2 (D[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (hfn_ipo_n5), .A2 (D[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (hfn_ipo_n5), .A2 (D[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (hfn_ipo_n5), .A2 (D[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (hfn_ipo_n5), .A2 (D[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (hfn_ipo_n5), .A2 (D[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (hfn_ipo_n5), .A2 (D[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (hfn_ipo_n5), .A2 (D[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (hfn_ipo_n5), .A2 (D[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (hfn_ipo_n5), .A2 (D[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (hfn_ipo_n5), .A2 (D[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (hfn_ipo_n5), .A2 (D[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (hfn_ipo_n5), .A2 (D[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (hfn_ipo_n5), .A2 (D[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (hfn_ipo_n5), .A2 (D[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (hfn_ipo_n5), .A2 (D[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (hfn_ipo_n5), .A2 (D[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (hfn_ipo_n5), .A2 (D[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (hfn_ipo_n5), .A2 (D[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (hfn_ipo_n5), .A2 (D[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (hfn_ipo_n5), .A2 (D[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (hfn_ipo_n5), .A2 (D[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (hfn_ipo_n5), .A2 (D[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (rst));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (rst));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (CTS_n_tid1_10), .D (n_2));
DFF_X1 \Q_reg[1]  (.Q (Q[1]), .CK (CTS_n_tid1_10), .D (n_3));
DFF_X1 \Q_reg[2]  (.Q (Q[2]), .CK (CTS_n_tid1_10), .D (n_4));
DFF_X1 \Q_reg[3]  (.Q (Q[3]), .CK (CTS_n_tid1_10), .D (n_5));
DFF_X1 \Q_reg[4]  (.Q (Q[4]), .CK (CTS_n_tid1_10), .D (n_6));
DFF_X1 \Q_reg[5]  (.Q (Q[5]), .CK (CTS_n_tid1_10), .D (n_7));
DFF_X1 \Q_reg[6]  (.Q (Q[6]), .CK (CTS_n_tid1_10), .D (n_8));
DFF_X1 \Q_reg[7]  (.Q (Q[7]), .CK (CTS_n_tid1_10), .D (n_9));
DFF_X1 \Q_reg[8]  (.Q (Q[8]), .CK (CTS_n_tid1_10), .D (n_10));
DFF_X1 \Q_reg[9]  (.Q (Q[9]), .CK (CTS_n_tid1_10), .D (n_11));
DFF_X1 \Q_reg[10]  (.Q (Q[10]), .CK (CTS_n_tid1_10), .D (n_12));
DFF_X1 \Q_reg[11]  (.Q (Q[11]), .CK (CTS_n_tid1_10), .D (n_13));
DFF_X1 \Q_reg[12]  (.Q (Q[12]), .CK (CTS_n_tid1_10), .D (n_14));
DFF_X1 \Q_reg[13]  (.Q (Q[13]), .CK (CTS_n_tid1_10), .D (n_15));
DFF_X1 \Q_reg[14]  (.Q (Q[14]), .CK (CTS_n_tid1_10), .D (n_16));
DFF_X1 \Q_reg[15]  (.Q (Q[15]), .CK (CTS_n_tid1_10), .D (n_17));
DFF_X1 \Q_reg[16]  (.Q (Q[16]), .CK (CTS_n_tid1_10), .D (n_18));
DFF_X1 \Q_reg[17]  (.Q (Q[17]), .CK (CTS_n_tid1_10), .D (n_19));
DFF_X1 \Q_reg[18]  (.Q (Q[18]), .CK (CTS_n_tid1_10), .D (n_20));
DFF_X1 \Q_reg[19]  (.Q (Q[19]), .CK (CTS_n_tid1_10), .D (n_21));
DFF_X1 \Q_reg[20]  (.Q (Q[20]), .CK (CTS_n_tid1_10), .D (n_22));
DFF_X1 \Q_reg[21]  (.Q (Q[21]), .CK (CTS_n_tid1_10), .D (n_23));
DFF_X1 \Q_reg[22]  (.Q (Q[22]), .CK (CTS_n_tid1_10), .D (n_24));
DFF_X1 \Q_reg[23]  (.Q (Q[23]), .CK (CTS_n_tid1_10), .D (n_25));
DFF_X1 \Q_reg[24]  (.Q (Q[24]), .CK (CTS_n_tid1_10), .D (n_26));
DFF_X1 \Q_reg[25]  (.Q (Q[25]), .CK (CTS_n_tid1_10), .D (n_27));
DFF_X1 \Q_reg[26]  (.Q (Q[26]), .CK (CTS_n_tid1_10), .D (n_28));
DFF_X1 \Q_reg[27]  (.Q (Q[27]), .CK (CTS_n_tid1_10), .D (n_29));
DFF_X1 \Q_reg[28]  (.Q (Q[28]), .CK (CTS_n_tid1_10), .D (n_30));
DFF_X1 \Q_reg[29]  (.Q (Q[29]), .CK (CTS_n_tid1_10), .D (n_31));
DFF_X1 \Q_reg[30]  (.Q (Q[30]), .CK (CTS_n_tid1_10), .D (n_32));
DFF_X1 \Q_reg[31]  (.Q (Q[31]), .CK (CTS_n_tid1_10), .D (n_33));
DFF_X1 \Q_reg[32]  (.Q (Q[32]), .CK (CTS_n_tid1_10), .D (n_34));
DFF_X1 \Q_reg[33]  (.Q (Q[33]), .CK (CTS_n_tid1_10), .D (n_35));
DFF_X1 \Q_reg[34]  (.Q (Q[34]), .CK (CTS_n_tid1_10), .D (n_36));
DFF_X1 \Q_reg[35]  (.Q (Q[35]), .CK (CTS_n_tid1_10), .D (n_37));
DFF_X1 \Q_reg[36]  (.Q (Q[36]), .CK (CTS_n_tid1_10), .D (n_38));
DFF_X1 \Q_reg[37]  (.Q (Q[37]), .CK (CTS_n_tid1_10), .D (n_39));
DFF_X1 \Q_reg[38]  (.Q (Q[38]), .CK (CTS_n_tid1_10), .D (n_40));
DFF_X1 \Q_reg[39]  (.Q (Q[39]), .CK (CTS_n_tid1_10), .D (n_41));
DFF_X1 \Q_reg[40]  (.Q (Q[40]), .CK (CTS_n_tid1_10), .D (n_42));
DFF_X1 \Q_reg[41]  (.Q (Q[41]), .CK (CTS_n_tid1_10), .D (n_43));
DFF_X1 \Q_reg[42]  (.Q (Q[42]), .CK (CTS_n_tid1_10), .D (n_44));
DFF_X1 \Q_reg[43]  (.Q (Q[43]), .CK (CTS_n_tid1_10), .D (n_45));
DFF_X1 \Q_reg[44]  (.Q (Q[44]), .CK (CTS_n_tid1_10), .D (n_46));
DFF_X1 \Q_reg[45]  (.Q (Q[45]), .CK (CTS_n_tid1_10), .D (n_47));
DFF_X1 \Q_reg[46]  (.Q (Q[46]), .CK (CTS_n_tid1_10), .D (n_48));
DFF_X1 \Q_reg[47]  (.Q (Q[47]), .CK (CTS_n_tid1_10), .D (n_49));
DFF_X1 \Q_reg[48]  (.Q (Q[48]), .CK (CTS_n_tid1_10), .D (n_50));
DFF_X1 \Q_reg[49]  (.Q (Q[49]), .CK (CTS_n_tid1_10), .D (n_51));
DFF_X1 \Q_reg[50]  (.Q (Q[50]), .CK (CTS_n_tid1_10), .D (n_52));
DFF_X1 \Q_reg[51]  (.Q (Q[51]), .CK (CTS_n_tid1_10), .D (n_53));
DFF_X1 \Q_reg[52]  (.Q (Q[52]), .CK (CTS_n_tid1_10), .D (n_54));
DFF_X1 \Q_reg[53]  (.Q (Q[53]), .CK (CTS_n_tid1_10), .D (n_55));
DFF_X1 \Q_reg[54]  (.Q (Q[54]), .CK (CTS_n_tid1_10), .D (n_56));
DFF_X1 \Q_reg[55]  (.Q (Q[55]), .CK (CTS_n_tid1_10), .D (n_57));
DFF_X1 \Q_reg[56]  (.Q (Q[56]), .CK (CTS_n_tid1_10), .D (n_58));
DFF_X1 \Q_reg[57]  (.Q (Q[57]), .CK (CTS_n_tid1_10), .D (n_59));
DFF_X1 \Q_reg[58]  (.Q (Q[58]), .CK (CTS_n_tid1_10), .D (n_60));
DFF_X1 \Q_reg[59]  (.Q (Q[59]), .CK (CTS_n_tid1_10), .D (n_61));
DFF_X1 \Q_reg[60]  (.Q (Q[60]), .CK (CTS_n_tid1_10), .D (n_62));
DFF_X1 \Q_reg[61]  (.Q (Q[61]), .CK (CTS_n_tid1_10), .D (n_63));
DFF_X1 \Q_reg[62]  (.Q (Q[62]), .CK (CTS_n_tid1_10), .D (n_64));
DFF_X1 \Q_reg[63]  (.Q (Q[63]), .CK (CTS_n_tid1_10), .D (n_65));
CLKGATETST_X8 clk_gate_Q_reg (.GCK (CTS_n_tid1_11), .CK (clk_CTS_0_PP_10), .E (n_1), .SE (1'b0 ));
BUF_X2 hfn_ipo_c5 (.Z (hfn_ipo_n5), .A (n_0_0));
CLKBUF_X3 CTS_L3_c_tid1_11 (.Z (CTS_n_tid1_10), .A (CTS_n_tid1_11));

endmodule //buffer__parameterized0

module buffer (clk_CTS_0_PP_11, clk, rst, en, D, Q);

output [31:0] Q;
input [31:0] D;
input clk;
input en;
input rst;
input clk_CTS_0_PP_11;
wire CLOCK_slh__n69;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CLOCK_slh__n70;
wire CLOCK_slh__n68;
wire CLOCK_slh__n74;
wire CLOCK_slh__n75;
wire CLOCK_slh__n76;
wire CLOCK_slh__n80;
wire CLOCK_slh__n81;
wire CLOCK_slh__n82;
wire CLOCK_slh__n86;
wire CLOCK_slh__n87;
wire CLOCK_slh__n88;
wire CLOCK_slh__n92;
wire CLOCK_slh__n93;
wire CLOCK_slh__n94;
wire CLOCK_slh__n98;
wire CLOCK_slh__n99;
wire CLOCK_slh__n100;
wire CLOCK_slh__n104;
wire CLOCK_slh__n105;
wire CLOCK_slh__n106;
wire CLOCK_slh__n110;
wire CLOCK_slh__n111;
wire CLOCK_slh__n112;
wire CLOCK_slh__n116;
wire CLOCK_slh__n117;
wire CLOCK_slh__n118;
wire CLOCK_slh__n122;
wire CLOCK_slh__n123;
wire CLOCK_slh__n124;
wire CLOCK_slh__n128;
wire CLOCK_slh__n129;
wire CLOCK_slh__n130;
wire CLOCK_slh__n134;
wire CLOCK_slh__n135;
wire CLOCK_slh__n136;
wire CLOCK_slh__n140;
wire CLOCK_slh__n141;
wire CLOCK_slh__n142;
wire CLOCK_slh__n146;
wire CLOCK_slh__n147;
wire CLOCK_slh__n148;
wire CLOCK_slh__n152;
wire CLOCK_slh__n153;
wire CLOCK_slh__n154;
wire CLOCK_slh__n158;
wire CLOCK_slh__n159;
wire CLOCK_slh__n160;
wire CLOCK_slh__n164;
wire CLOCK_slh__n165;
wire CLOCK_slh__n166;
wire CLOCK_slh__n170;
wire CLOCK_slh__n171;
wire CLOCK_slh__n172;
wire CLOCK_slh__n176;
wire CLOCK_slh__n177;
wire CLOCK_slh__n178;
wire CLOCK_slh__n182;
wire CLOCK_slh__n183;
wire CLOCK_slh__n184;
wire CLOCK_slh__n188;
wire CLOCK_slh__n189;
wire CLOCK_slh__n190;
wire CLOCK_slh__n194;
wire CLOCK_slh__n195;
wire CLOCK_slh__n196;
wire CLOCK_slh__n200;
wire CLOCK_slh__n201;
wire CLOCK_slh__n202;
wire CLOCK_slh__n206;
wire CLOCK_slh__n207;
wire CLOCK_slh__n208;
wire CLOCK_slh__n209;
wire CLOCK_slh__n210;
wire CLOCK_slh__n211;
wire CLOCK_slh__n212;
wire CLOCK_slh__n213;
wire CLOCK_slh__n214;
wire CLOCK_slh__n215;
wire CLOCK_slh__n216;
wire CLOCK_slh__n217;
wire CLOCK_slh__n218;
wire CLOCK_slh__n219;
wire CLOCK_slh__n220;
wire CLOCK_slh__n221;
wire CLOCK_slh__n222;
wire CLOCK_slh__n223;
wire CLOCK_slh__n224;
wire CLOCK_slh__n225;
wire CLOCK_slh__n226;
wire CLOCK_slh__n227;
wire CLOCK_slh__n228;
wire CLOCK_slh__n229;
wire CLOCK_slh__n230;
wire CLOCK_slh__n231;
wire CLOCK_slh__n232;
wire CLOCK_sph__n254;
wire CLOCK_sph__n256;
wire CLOCK_sph__n258;
wire CLOCK_sph__n260;
wire CLOCK_sph__n262;
wire CLOCK_sph__n264;
wire CLOCK_sph__n266;
wire CLOCK_sph__n268;
wire CLOCK_sph__n270;
wire CLOCK_sph__n272;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n86), .A1 (n_0_0), .A2 (D[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n212), .A1 (n_0_0), .A2 (D[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n221), .A1 (n_0_0), .A2 (D[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n182), .A1 (n_0_0), .A2 (D[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n110), .A1 (n_0_0), .A2 (D[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n74), .A1 (n_0_0), .A2 (D[26]));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n134), .A1 (n_0_0), .A2 (D[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n152), .A1 (n_0_0), .A2 (D[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n116), .A1 (n_0_0), .A2 (D[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n170), .A1 (n_0_0), .A2 (D[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n209), .A1 (n_0_0), .A2 (D[21]));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n92), .A1 (n_0_0), .A2 (D[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n146), .A1 (n_0_0), .A2 (D[19]));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n98), .A1 (n_0_0), .A2 (D[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n230), .A1 (n_0_0), .A2 (D[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n140), .A1 (n_0_0), .A2 (D[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n68), .A1 (n_0_0), .A2 (D[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n218), .A1 (n_0_0), .A2 (D[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n206), .A1 (n_0_0), .A2 (D[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n128), .A1 (n_0_0), .A2 (D[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n164), .A1 (n_0_0), .A2 (D[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n200), .A1 (n_0_0), .A2 (D[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n227), .A1 (n_0_0), .A2 (D[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n176), .A1 (n_0_0), .A2 (D[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n80), .A1 (n_0_0), .A2 (D[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n194), .A1 (n_0_0), .A2 (D[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n158), .A1 (n_0_0), .A2 (D[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n104), .A1 (n_0_0), .A2 (D[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n122), .A1 (n_0_0), .A2 (D[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n224), .A1 (n_0_0), .A2 (D[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n188), .A1 (n_0_0), .A2 (D[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n215), .A1 (n_0_0), .A2 (D[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (rst));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (rst));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (n_0), .D (n_2));
DFF_X1 \Q_reg[1]  (.Q (Q[1]), .CK (n_0), .D (n_3));
DFF_X1 \Q_reg[2]  (.Q (Q[2]), .CK (n_0), .D (n_4));
DFF_X1 \Q_reg[3]  (.Q (Q[3]), .CK (n_0), .D (n_5));
DFF_X1 \Q_reg[4]  (.Q (Q[4]), .CK (n_0), .D (n_6));
DFF_X1 \Q_reg[5]  (.Q (Q[5]), .CK (n_0), .D (n_7));
DFF_X1 \Q_reg[6]  (.Q (Q[6]), .CK (n_0), .D (n_8));
DFF_X1 \Q_reg[7]  (.Q (Q[7]), .CK (n_0), .D (n_9));
DFF_X1 \Q_reg[8]  (.Q (Q[8]), .CK (n_0), .D (n_10));
DFF_X1 \Q_reg[9]  (.Q (Q[9]), .CK (n_0), .D (n_11));
DFF_X1 \Q_reg[10]  (.Q (Q[10]), .CK (n_0), .D (n_12));
DFF_X1 \Q_reg[11]  (.Q (Q[11]), .CK (n_0), .D (n_13));
DFF_X1 \Q_reg[12]  (.Q (Q[12]), .CK (n_0), .D (n_14));
DFF_X1 \Q_reg[13]  (.Q (Q[13]), .CK (n_0), .D (n_15));
DFF_X1 \Q_reg[14]  (.Q (Q[14]), .CK (n_0), .D (n_16));
DFF_X1 \Q_reg[15]  (.Q (Q[15]), .CK (n_0), .D (n_17));
DFF_X1 \Q_reg[16]  (.Q (Q[16]), .CK (n_0), .D (n_18));
DFF_X1 \Q_reg[17]  (.Q (Q[17]), .CK (n_0), .D (n_19));
DFF_X1 \Q_reg[18]  (.Q (Q[18]), .CK (n_0), .D (n_20));
DFF_X1 \Q_reg[19]  (.Q (Q[19]), .CK (n_0), .D (n_21));
DFF_X1 \Q_reg[20]  (.Q (Q[20]), .CK (n_0), .D (n_22));
DFF_X1 \Q_reg[21]  (.Q (Q[21]), .CK (n_0), .D (n_23));
DFF_X1 \Q_reg[22]  (.Q (Q[22]), .CK (n_0), .D (n_24));
DFF_X1 \Q_reg[23]  (.Q (Q[23]), .CK (n_0), .D (n_25));
DFF_X1 \Q_reg[24]  (.Q (Q[24]), .CK (n_0), .D (n_26));
DFF_X1 \Q_reg[25]  (.Q (Q[25]), .CK (n_0), .D (n_27));
DFF_X1 \Q_reg[26]  (.Q (Q[26]), .CK (n_0), .D (n_28));
DFF_X1 \Q_reg[27]  (.Q (Q[27]), .CK (n_0), .D (n_29));
DFF_X1 \Q_reg[28]  (.Q (Q[28]), .CK (n_0), .D (n_30));
DFF_X1 \Q_reg[29]  (.Q (Q[29]), .CK (n_0), .D (n_31));
DFF_X1 \Q_reg[30]  (.Q (Q[30]), .CK (n_0), .D (n_32));
DFF_X1 \Q_reg[31]  (.Q (Q[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_Q_reg (.GCK (n_0), .CK (clk_CTS_0_PP_11), .E (n_1), .SE (1'b0 ));
CLKBUF_X1 CLOCK_slh__c17 (.Z (CLOCK_slh__n69), .A (CLOCK_slh__n68));
CLKBUF_X1 CLOCK_slh__c18 (.Z (CLOCK_slh__n70), .A (CLOCK_slh__n69));
CLKBUF_X1 CLOCK_slh__c19 (.Z (n_17), .A (CLOCK_slh__n70));
CLKBUF_X1 CLOCK_slh__c23 (.Z (CLOCK_slh__n75), .A (CLOCK_slh__n74));
CLKBUF_X1 CLOCK_slh__c24 (.Z (CLOCK_slh__n76), .A (CLOCK_slh__n75));
CLKBUF_X1 CLOCK_slh__c25 (.Z (n_28), .A (CLOCK_slh__n76));
CLKBUF_X1 CLOCK_slh__c29 (.Z (CLOCK_slh__n81), .A (CLOCK_slh__n80));
CLKBUF_X1 CLOCK_slh__c30 (.Z (CLOCK_slh__n82), .A (CLOCK_slh__n81));
CLKBUF_X1 CLOCK_slh__c31 (.Z (n_9), .A (CLOCK_slh__n82));
CLKBUF_X1 CLOCK_slh__c35 (.Z (CLOCK_slh__n87), .A (CLOCK_slh__n86));
CLKBUF_X1 CLOCK_slh__c36 (.Z (CLOCK_slh__n88), .A (CLOCK_slh__n87));
CLKBUF_X1 CLOCK_slh__c37 (.Z (n_33), .A (CLOCK_slh__n88));
CLKBUF_X1 CLOCK_slh__c41 (.Z (CLOCK_slh__n93), .A (CLOCK_slh__n92));
CLKBUF_X1 CLOCK_slh__c42 (.Z (CLOCK_slh__n94), .A (CLOCK_slh__n93));
CLKBUF_X1 CLOCK_slh__c43 (.Z (n_22), .A (CLOCK_slh__n94));
CLKBUF_X1 CLOCK_slh__c47 (.Z (CLOCK_slh__n99), .A (CLOCK_slh__n98));
CLKBUF_X1 CLOCK_slh__c48 (.Z (CLOCK_slh__n100), .A (CLOCK_slh__n99));
CLKBUF_X1 CLOCK_slh__c49 (.Z (n_20), .A (CLOCK_slh__n100));
CLKBUF_X1 CLOCK_slh__c53 (.Z (CLOCK_slh__n105), .A (CLOCK_slh__n104));
CLKBUF_X1 CLOCK_slh__c54 (.Z (CLOCK_slh__n106), .A (CLOCK_slh__n105));
CLKBUF_X1 CLOCK_slh__c55 (.Z (n_6), .A (CLOCK_slh__n106));
CLKBUF_X1 CLOCK_slh__c59 (.Z (CLOCK_slh__n111), .A (CLOCK_slh__n110));
CLKBUF_X1 CLOCK_slh__c60 (.Z (CLOCK_slh__n112), .A (CLOCK_slh__n111));
CLKBUF_X1 CLOCK_slh__c61 (.Z (n_29), .A (CLOCK_slh__n112));
CLKBUF_X1 CLOCK_slh__c65 (.Z (CLOCK_slh__n117), .A (CLOCK_slh__n116));
CLKBUF_X1 CLOCK_slh__c66 (.Z (CLOCK_slh__n118), .A (CLOCK_slh__n117));
CLKBUF_X1 CLOCK_slh__c67 (.Z (CLOCK_sph__n262), .A (CLOCK_slh__n118));
CLKBUF_X1 CLOCK_slh__c71 (.Z (CLOCK_slh__n123), .A (CLOCK_slh__n122));
CLKBUF_X1 CLOCK_slh__c72 (.Z (CLOCK_slh__n124), .A (CLOCK_slh__n123));
CLKBUF_X1 CLOCK_slh__c73 (.Z (n_5), .A (CLOCK_slh__n124));
CLKBUF_X1 CLOCK_slh__c77 (.Z (CLOCK_slh__n129), .A (CLOCK_slh__n128));
CLKBUF_X1 CLOCK_slh__c78 (.Z (CLOCK_slh__n130), .A (CLOCK_slh__n129));
CLKBUF_X1 CLOCK_slh__c79 (.Z (n_14), .A (CLOCK_slh__n130));
CLKBUF_X1 CLOCK_slh__c83 (.Z (CLOCK_slh__n135), .A (CLOCK_slh__n134));
CLKBUF_X1 CLOCK_slh__c84 (.Z (CLOCK_slh__n136), .A (CLOCK_slh__n135));
CLKBUF_X1 CLOCK_slh__c85 (.Z (CLOCK_sph__n258), .A (CLOCK_slh__n136));
CLKBUF_X1 CLOCK_slh__c89 (.Z (CLOCK_slh__n141), .A (CLOCK_slh__n140));
CLKBUF_X1 CLOCK_slh__c90 (.Z (CLOCK_slh__n142), .A (CLOCK_slh__n141));
CLKBUF_X1 CLOCK_slh__c91 (.Z (n_18), .A (CLOCK_slh__n142));
CLKBUF_X1 CLOCK_slh__c95 (.Z (CLOCK_slh__n147), .A (CLOCK_slh__n146));
CLKBUF_X1 CLOCK_slh__c96 (.Z (CLOCK_slh__n148), .A (CLOCK_slh__n147));
CLKBUF_X1 CLOCK_slh__c97 (.Z (n_21), .A (CLOCK_slh__n148));
CLKBUF_X1 CLOCK_slh__c101 (.Z (CLOCK_slh__n153), .A (CLOCK_slh__n152));
CLKBUF_X1 CLOCK_slh__c102 (.Z (CLOCK_slh__n154), .A (CLOCK_slh__n153));
CLKBUF_X1 CLOCK_slh__c103 (.Z (CLOCK_sph__n266), .A (CLOCK_slh__n154));
CLKBUF_X1 CLOCK_slh__c107 (.Z (CLOCK_slh__n159), .A (CLOCK_slh__n158));
CLKBUF_X1 CLOCK_slh__c108 (.Z (CLOCK_slh__n160), .A (CLOCK_slh__n159));
CLKBUF_X1 CLOCK_slh__c109 (.Z (n_7), .A (CLOCK_slh__n160));
CLKBUF_X1 CLOCK_slh__c113 (.Z (CLOCK_slh__n165), .A (CLOCK_slh__n164));
CLKBUF_X1 CLOCK_slh__c114 (.Z (CLOCK_slh__n166), .A (CLOCK_slh__n165));
CLKBUF_X1 CLOCK_slh__c115 (.Z (n_13), .A (CLOCK_slh__n166));
CLKBUF_X1 CLOCK_slh__c119 (.Z (CLOCK_slh__n171), .A (CLOCK_slh__n170));
CLKBUF_X1 CLOCK_slh__c120 (.Z (CLOCK_slh__n172), .A (CLOCK_slh__n171));
CLKBUF_X1 CLOCK_slh__c121 (.Z (CLOCK_sph__n268), .A (CLOCK_slh__n172));
CLKBUF_X1 CLOCK_slh__c125 (.Z (CLOCK_slh__n177), .A (CLOCK_slh__n176));
CLKBUF_X1 CLOCK_slh__c126 (.Z (CLOCK_slh__n178), .A (CLOCK_slh__n177));
CLKBUF_X1 CLOCK_slh__c127 (.Z (CLOCK_sph__n264), .A (CLOCK_slh__n178));
CLKBUF_X1 CLOCK_slh__c131 (.Z (CLOCK_slh__n183), .A (CLOCK_slh__n182));
CLKBUF_X1 CLOCK_slh__c132 (.Z (CLOCK_slh__n184), .A (CLOCK_slh__n183));
CLKBUF_X1 CLOCK_slh__c133 (.Z (CLOCK_sph__n272), .A (CLOCK_slh__n184));
CLKBUF_X1 CLOCK_slh__c137 (.Z (CLOCK_slh__n189), .A (CLOCK_slh__n188));
CLKBUF_X1 CLOCK_slh__c138 (.Z (CLOCK_slh__n190), .A (CLOCK_slh__n189));
CLKBUF_X1 CLOCK_slh__c139 (.Z (n_3), .A (CLOCK_slh__n190));
CLKBUF_X1 CLOCK_slh__c143 (.Z (CLOCK_slh__n195), .A (CLOCK_slh__n194));
CLKBUF_X1 CLOCK_slh__c144 (.Z (CLOCK_slh__n196), .A (CLOCK_slh__n195));
CLKBUF_X1 CLOCK_slh__c145 (.Z (CLOCK_sph__n256), .A (CLOCK_slh__n196));
CLKBUF_X1 CLOCK_slh__c149 (.Z (CLOCK_slh__n201), .A (CLOCK_slh__n200));
CLKBUF_X1 CLOCK_slh__c150 (.Z (CLOCK_slh__n202), .A (CLOCK_slh__n201));
CLKBUF_X1 CLOCK_slh__c151 (.Z (n_12), .A (CLOCK_slh__n202));
CLKBUF_X1 CLOCK_slh__c155 (.Z (CLOCK_slh__n207), .A (CLOCK_slh__n206));
CLKBUF_X1 CLOCK_slh__c156 (.Z (CLOCK_slh__n208), .A (CLOCK_slh__n207));
CLKBUF_X1 CLOCK_slh__c157 (.Z (n_15), .A (CLOCK_slh__n208));
CLKBUF_X1 CLOCK_slh__c158 (.Z (CLOCK_slh__n210), .A (CLOCK_slh__n209));
CLKBUF_X1 CLOCK_slh__c159 (.Z (CLOCK_slh__n211), .A (CLOCK_slh__n210));
CLKBUF_X1 CLOCK_slh__c160 (.Z (n_23), .A (CLOCK_slh__n211));
CLKBUF_X1 CLOCK_slh__c161 (.Z (CLOCK_slh__n213), .A (CLOCK_slh__n212));
CLKBUF_X1 CLOCK_slh__c162 (.Z (CLOCK_slh__n214), .A (CLOCK_slh__n213));
CLKBUF_X1 CLOCK_slh__c163 (.Z (n_32), .A (CLOCK_slh__n214));
CLKBUF_X1 CLOCK_slh__c164 (.Z (CLOCK_slh__n216), .A (CLOCK_slh__n215));
CLKBUF_X1 CLOCK_slh__c165 (.Z (CLOCK_slh__n217), .A (CLOCK_slh__n216));
CLKBUF_X1 CLOCK_slh__c166 (.Z (CLOCK_sph__n254), .A (CLOCK_slh__n217));
CLKBUF_X1 CLOCK_slh__c167 (.Z (CLOCK_slh__n219), .A (CLOCK_slh__n218));
CLKBUF_X1 CLOCK_slh__c168 (.Z (CLOCK_slh__n220), .A (CLOCK_slh__n219));
CLKBUF_X1 CLOCK_slh__c169 (.Z (CLOCK_sph__n260), .A (CLOCK_slh__n220));
CLKBUF_X1 CLOCK_slh__c170 (.Z (CLOCK_slh__n222), .A (CLOCK_slh__n221));
CLKBUF_X1 CLOCK_slh__c171 (.Z (CLOCK_slh__n223), .A (CLOCK_slh__n222));
CLKBUF_X1 CLOCK_slh__c172 (.Z (CLOCK_sph__n270), .A (CLOCK_slh__n223));
CLKBUF_X1 CLOCK_slh__c173 (.Z (CLOCK_slh__n225), .A (CLOCK_slh__n224));
CLKBUF_X1 CLOCK_slh__c174 (.Z (CLOCK_slh__n226), .A (CLOCK_slh__n225));
CLKBUF_X1 CLOCK_slh__c175 (.Z (n_4), .A (CLOCK_slh__n226));
CLKBUF_X1 CLOCK_slh__c176 (.Z (CLOCK_slh__n228), .A (CLOCK_slh__n227));
CLKBUF_X1 CLOCK_slh__c177 (.Z (CLOCK_slh__n229), .A (CLOCK_slh__n228));
CLKBUF_X1 CLOCK_slh__c178 (.Z (n_11), .A (CLOCK_slh__n229));
CLKBUF_X1 CLOCK_slh__c179 (.Z (CLOCK_slh__n231), .A (CLOCK_slh__n230));
CLKBUF_X1 CLOCK_slh__c180 (.Z (CLOCK_slh__n232), .A (CLOCK_slh__n231));
CLKBUF_X1 CLOCK_slh__c181 (.Z (n_19), .A (CLOCK_slh__n232));
CLKBUF_X1 CLOCK_sph__c203 (.Z (n_2), .A (CLOCK_sph__n254));
CLKBUF_X1 CLOCK_sph__c205 (.Z (n_8), .A (CLOCK_sph__n256));
CLKBUF_X1 CLOCK_sph__c207 (.Z (n_27), .A (CLOCK_sph__n258));
CLKBUF_X1 CLOCK_sph__c209 (.Z (n_16), .A (CLOCK_sph__n260));
CLKBUF_X1 CLOCK_sph__c211 (.Z (n_25), .A (CLOCK_sph__n262));
CLKBUF_X1 CLOCK_sph__c213 (.Z (n_10), .A (CLOCK_sph__n264));
CLKBUF_X1 CLOCK_sph__c215 (.Z (n_26), .A (CLOCK_sph__n266));
CLKBUF_X1 CLOCK_sph__c217 (.Z (n_24), .A (CLOCK_sph__n268));
CLKBUF_X1 CLOCK_sph__c219 (.Z (n_31), .A (CLOCK_sph__n270));
CLKBUF_X1 CLOCK_sph__c221 (.Z (n_30), .A (CLOCK_sph__n272));

endmodule //buffer

module buffer__0_18 (clk_CTS_0_PP_10, clk, rst, en, D, Q);

output [31:0] Q;
input [31:0] D;
input clk;
input en;
input rst;
input clk_CTS_0_PP_10;
wire CLOCK_slh__n62;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CLOCK_slh__n61;
wire CLOCK_slh__n63;
wire CLOCK_slh__n67;
wire CLOCK_slh__n68;
wire CLOCK_slh__n69;
wire CLOCK_slh__n73;
wire CLOCK_slh__n74;
wire CLOCK_slh__n75;
wire CLOCK_slh__n79;
wire CLOCK_slh__n80;
wire CLOCK_slh__n81;
wire CLOCK_slh__n85;
wire CLOCK_slh__n86;
wire CLOCK_slh__n87;
wire CLOCK_slh__n91;
wire CLOCK_slh__n92;
wire CLOCK_slh__n93;
wire CLOCK_slh__n97;
wire CLOCK_slh__n98;
wire CLOCK_slh__n99;
wire CLOCK_slh__n103;
wire CLOCK_slh__n104;
wire CLOCK_slh__n105;
wire CLOCK_slh__n109;
wire CLOCK_slh__n110;
wire CLOCK_slh__n111;
wire CLOCK_slh__n115;
wire CLOCK_slh__n116;
wire CLOCK_slh__n117;
wire CLOCK_slh__n121;
wire CLOCK_slh__n122;
wire CLOCK_slh__n123;
wire CLOCK_slh__n127;
wire CLOCK_slh__n128;
wire CLOCK_slh__n129;
wire CLOCK_slh__n133;
wire CLOCK_slh__n134;
wire CLOCK_slh__n135;
wire CLOCK_slh__n139;
wire CLOCK_slh__n140;
wire CLOCK_slh__n141;
wire CLOCK_slh__n145;
wire CLOCK_slh__n146;
wire CLOCK_slh__n147;
wire CLOCK_slh__n151;
wire CLOCK_slh__n152;
wire CLOCK_slh__n153;
wire CLOCK_slh__n157;
wire CLOCK_slh__n158;
wire CLOCK_slh__n159;
wire CLOCK_slh__n163;
wire CLOCK_slh__n164;
wire CLOCK_slh__n165;
wire CLOCK_slh__n169;
wire CLOCK_slh__n170;
wire CLOCK_slh__n171;
wire CLOCK_slh__n175;
wire CLOCK_slh__n176;
wire CLOCK_slh__n177;
wire CLOCK_slh__n181;
wire CLOCK_slh__n182;
wire CLOCK_slh__n183;
wire CLOCK_slh__n187;
wire CLOCK_slh__n188;
wire CLOCK_slh__n189;
wire CLOCK_slh__n193;
wire CLOCK_slh__n194;
wire CLOCK_slh__n195;
wire CLOCK_slh__n199;
wire CLOCK_slh__n200;
wire CLOCK_slh__n201;
wire CLOCK_slh__n205;
wire CLOCK_slh__n206;
wire CLOCK_slh__n207;
wire CLOCK_slh__n211;
wire CLOCK_slh__n212;
wire CLOCK_slh__n213;
wire CLOCK_slh__n217;
wire CLOCK_slh__n218;
wire CLOCK_slh__n219;
wire CLOCK_slh__n223;
wire CLOCK_slh__n224;
wire CLOCK_slh__n225;
wire CLOCK_slh__n229;
wire CLOCK_slh__n230;
wire CLOCK_slh__n231;
wire CLOCK_slh__n235;
wire CLOCK_slh__n236;
wire CLOCK_slh__n237;
wire CLOCK_slh__n238;
wire CLOCK_slh__n239;
wire CLOCK_slh__n240;
wire CLOCK_slh__n241;
wire CLOCK_slh__n242;
wire CLOCK_slh__n243;
wire CLOCK_sph__n244;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n223), .A1 (n_0_0), .A2 (D[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n175), .A1 (n_0_0), .A2 (D[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n235), .A1 (n_0_0), .A2 (D[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n238), .A1 (n_0_0), .A2 (D[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n229), .A1 (n_0_0), .A2 (D[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n217), .A1 (n_0_0), .A2 (D[26]));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n157), .A1 (n_0_0), .A2 (D[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n109), .A1 (n_0_0), .A2 (D[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n199), .A1 (n_0_0), .A2 (D[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n211), .A1 (n_0_0), .A2 (D[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n205), .A1 (n_0_0), .A2 (D[21]));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n193), .A1 (n_0_0), .A2 (D[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n139), .A1 (n_0_0), .A2 (D[19]));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n61), .A1 (n_0_0), .A2 (D[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n91), .A1 (n_0_0), .A2 (D[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n85), .A1 (n_0_0), .A2 (D[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n169), .A1 (n_0_0), .A2 (D[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n187), .A1 (n_0_0), .A2 (D[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n241), .A1 (n_0_0), .A2 (D[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n151), .A1 (n_0_0), .A2 (D[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n97), .A1 (n_0_0), .A2 (D[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n115), .A1 (n_0_0), .A2 (D[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n79), .A1 (n_0_0), .A2 (D[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n73), .A1 (n_0_0), .A2 (D[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n145), .A1 (n_0_0), .A2 (D[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n163), .A1 (n_0_0), .A2 (D[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n127), .A1 (n_0_0), .A2 (D[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n121), .A1 (n_0_0), .A2 (D[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n67), .A1 (n_0_0), .A2 (D[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n181), .A1 (n_0_0), .A2 (D[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n133), .A1 (n_0_0), .A2 (D[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n103), .A1 (n_0_0), .A2 (D[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (rst));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (rst));
DFF_X1 \Q_reg[0]  (.Q (Q[0]), .CK (n_0), .D (n_2));
DFF_X1 \Q_reg[1]  (.Q (Q[1]), .CK (n_0), .D (n_3));
DFF_X1 \Q_reg[2]  (.Q (Q[2]), .CK (n_0), .D (n_4));
DFF_X1 \Q_reg[3]  (.Q (Q[3]), .CK (n_0), .D (n_5));
DFF_X1 \Q_reg[4]  (.Q (Q[4]), .CK (n_0), .D (n_6));
DFF_X1 \Q_reg[5]  (.Q (Q[5]), .CK (n_0), .D (n_7));
DFF_X1 \Q_reg[6]  (.Q (Q[6]), .CK (n_0), .D (n_8));
DFF_X1 \Q_reg[7]  (.Q (Q[7]), .CK (n_0), .D (n_9));
DFF_X1 \Q_reg[8]  (.Q (Q[8]), .CK (n_0), .D (n_10));
DFF_X1 \Q_reg[9]  (.Q (Q[9]), .CK (n_0), .D (n_11));
DFF_X1 \Q_reg[10]  (.Q (Q[10]), .CK (n_0), .D (n_12));
DFF_X1 \Q_reg[11]  (.Q (Q[11]), .CK (n_0), .D (n_13));
DFF_X1 \Q_reg[12]  (.Q (Q[12]), .CK (n_0), .D (n_14));
DFF_X1 \Q_reg[13]  (.Q (Q[13]), .CK (n_0), .D (n_15));
DFF_X1 \Q_reg[14]  (.Q (Q[14]), .CK (n_0), .D (n_16));
DFF_X1 \Q_reg[15]  (.Q (Q[15]), .CK (n_0), .D (n_17));
DFF_X1 \Q_reg[16]  (.Q (Q[16]), .CK (n_0), .D (n_18));
DFF_X1 \Q_reg[17]  (.Q (Q[17]), .CK (n_0), .D (n_19));
DFF_X1 \Q_reg[18]  (.Q (Q[18]), .CK (n_0), .D (n_20));
DFF_X1 \Q_reg[19]  (.Q (Q[19]), .CK (n_0), .D (n_21));
DFF_X1 \Q_reg[20]  (.Q (Q[20]), .CK (n_0), .D (n_22));
DFF_X1 \Q_reg[21]  (.Q (Q[21]), .CK (n_0), .D (n_23));
DFF_X1 \Q_reg[22]  (.Q (Q[22]), .CK (n_0), .D (n_24));
DFF_X1 \Q_reg[23]  (.Q (Q[23]), .CK (n_0), .D (n_25));
DFF_X1 \Q_reg[24]  (.Q (Q[24]), .CK (n_0), .D (n_26));
DFF_X1 \Q_reg[25]  (.Q (Q[25]), .CK (n_0), .D (n_27));
DFF_X1 \Q_reg[26]  (.Q (Q[26]), .CK (n_0), .D (n_28));
DFF_X1 \Q_reg[27]  (.Q (Q[27]), .CK (n_0), .D (n_29));
DFF_X1 \Q_reg[28]  (.Q (Q[28]), .CK (n_0), .D (n_30));
DFF_X1 \Q_reg[29]  (.Q (Q[29]), .CK (n_0), .D (n_31));
DFF_X1 \Q_reg[30]  (.Q (Q[30]), .CK (n_0), .D (n_32));
DFF_X1 \Q_reg[31]  (.Q (Q[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_Q_reg (.GCK (n_0), .CK (clk_CTS_0_PP_10), .E (n_1), .SE (1'b0 ));
CLKBUF_X1 CLOCK_slh__c7 (.Z (CLOCK_slh__n62), .A (CLOCK_slh__n61));
CLKBUF_X1 CLOCK_slh__c8 (.Z (CLOCK_slh__n63), .A (CLOCK_slh__n62));
CLKBUF_X1 CLOCK_slh__c9 (.Z (n_20), .A (CLOCK_slh__n63));
CLKBUF_X1 CLOCK_slh__c13 (.Z (CLOCK_slh__n68), .A (CLOCK_slh__n67));
CLKBUF_X1 CLOCK_slh__c14 (.Z (CLOCK_slh__n69), .A (CLOCK_slh__n68));
CLKBUF_X1 CLOCK_slh__c15 (.Z (n_5), .A (CLOCK_slh__n69));
CLKBUF_X1 CLOCK_slh__c19 (.Z (CLOCK_slh__n74), .A (CLOCK_slh__n73));
CLKBUF_X1 CLOCK_slh__c20 (.Z (CLOCK_slh__n75), .A (CLOCK_slh__n74));
CLKBUF_X1 CLOCK_slh__c21 (.Z (n_10), .A (CLOCK_slh__n75));
CLKBUF_X1 CLOCK_slh__c25 (.Z (CLOCK_slh__n80), .A (CLOCK_slh__n79));
CLKBUF_X1 CLOCK_slh__c26 (.Z (CLOCK_slh__n81), .A (CLOCK_slh__n80));
CLKBUF_X1 CLOCK_slh__c27 (.Z (n_11), .A (CLOCK_slh__n81));
CLKBUF_X1 CLOCK_slh__c31 (.Z (CLOCK_slh__n86), .A (CLOCK_slh__n85));
CLKBUF_X1 CLOCK_slh__c32 (.Z (CLOCK_slh__n87), .A (CLOCK_slh__n86));
CLKBUF_X1 CLOCK_slh__c33 (.Z (n_18), .A (CLOCK_slh__n87));
CLKBUF_X1 CLOCK_slh__c37 (.Z (CLOCK_slh__n92), .A (CLOCK_slh__n91));
CLKBUF_X1 CLOCK_slh__c38 (.Z (CLOCK_slh__n93), .A (CLOCK_slh__n92));
CLKBUF_X1 CLOCK_slh__c39 (.Z (n_19), .A (CLOCK_slh__n93));
CLKBUF_X1 CLOCK_slh__c43 (.Z (CLOCK_slh__n98), .A (CLOCK_slh__n97));
CLKBUF_X1 CLOCK_slh__c44 (.Z (CLOCK_slh__n99), .A (CLOCK_slh__n98));
CLKBUF_X1 CLOCK_slh__c45 (.Z (n_13), .A (CLOCK_slh__n99));
CLKBUF_X1 CLOCK_slh__c49 (.Z (CLOCK_slh__n104), .A (CLOCK_slh__n103));
CLKBUF_X1 CLOCK_slh__c50 (.Z (CLOCK_slh__n105), .A (CLOCK_slh__n104));
CLKBUF_X1 CLOCK_slh__c51 (.Z (n_2), .A (CLOCK_slh__n105));
CLKBUF_X1 CLOCK_slh__c55 (.Z (CLOCK_slh__n110), .A (CLOCK_slh__n109));
CLKBUF_X1 CLOCK_slh__c56 (.Z (CLOCK_slh__n111), .A (CLOCK_slh__n110));
CLKBUF_X1 CLOCK_slh__c57 (.Z (n_26), .A (CLOCK_slh__n111));
CLKBUF_X1 CLOCK_slh__c61 (.Z (CLOCK_slh__n116), .A (CLOCK_slh__n115));
CLKBUF_X1 CLOCK_slh__c62 (.Z (CLOCK_slh__n117), .A (CLOCK_slh__n116));
CLKBUF_X1 CLOCK_slh__c63 (.Z (n_12), .A (CLOCK_slh__n117));
CLKBUF_X1 CLOCK_slh__c67 (.Z (CLOCK_slh__n122), .A (CLOCK_slh__n121));
CLKBUF_X1 CLOCK_slh__c68 (.Z (CLOCK_slh__n123), .A (CLOCK_slh__n122));
CLKBUF_X1 CLOCK_slh__c69 (.Z (n_6), .A (CLOCK_slh__n123));
CLKBUF_X1 CLOCK_slh__c73 (.Z (CLOCK_slh__n128), .A (CLOCK_slh__n127));
CLKBUF_X1 CLOCK_slh__c74 (.Z (CLOCK_slh__n129), .A (CLOCK_slh__n128));
CLKBUF_X1 CLOCK_slh__c75 (.Z (n_7), .A (CLOCK_slh__n129));
CLKBUF_X1 CLOCK_slh__c79 (.Z (CLOCK_slh__n134), .A (CLOCK_slh__n133));
CLKBUF_X1 CLOCK_slh__c80 (.Z (CLOCK_slh__n135), .A (CLOCK_slh__n134));
CLKBUF_X1 CLOCK_slh__c81 (.Z (n_3), .A (CLOCK_slh__n135));
CLKBUF_X1 CLOCK_slh__c85 (.Z (CLOCK_slh__n140), .A (CLOCK_slh__n139));
CLKBUF_X1 CLOCK_slh__c86 (.Z (CLOCK_slh__n141), .A (CLOCK_slh__n140));
CLKBUF_X1 CLOCK_slh__c87 (.Z (n_21), .A (CLOCK_slh__n141));
CLKBUF_X1 CLOCK_slh__c91 (.Z (CLOCK_slh__n146), .A (CLOCK_slh__n145));
CLKBUF_X1 CLOCK_slh__c92 (.Z (CLOCK_slh__n147), .A (CLOCK_slh__n146));
CLKBUF_X1 CLOCK_slh__c93 (.Z (n_9), .A (CLOCK_slh__n147));
CLKBUF_X1 CLOCK_slh__c97 (.Z (CLOCK_slh__n152), .A (CLOCK_slh__n151));
CLKBUF_X1 CLOCK_slh__c98 (.Z (CLOCK_slh__n153), .A (CLOCK_slh__n152));
CLKBUF_X1 CLOCK_slh__c99 (.Z (n_14), .A (CLOCK_slh__n153));
CLKBUF_X1 CLOCK_slh__c103 (.Z (CLOCK_slh__n158), .A (CLOCK_slh__n157));
CLKBUF_X1 CLOCK_slh__c104 (.Z (CLOCK_slh__n159), .A (CLOCK_slh__n158));
CLKBUF_X1 CLOCK_slh__c105 (.Z (n_27), .A (CLOCK_slh__n159));
CLKBUF_X1 CLOCK_slh__c109 (.Z (CLOCK_slh__n164), .A (CLOCK_slh__n163));
CLKBUF_X1 CLOCK_slh__c110 (.Z (CLOCK_slh__n165), .A (CLOCK_slh__n164));
CLKBUF_X1 CLOCK_slh__c111 (.Z (n_8), .A (CLOCK_slh__n165));
CLKBUF_X1 CLOCK_slh__c115 (.Z (CLOCK_slh__n170), .A (CLOCK_slh__n169));
CLKBUF_X1 CLOCK_slh__c116 (.Z (CLOCK_slh__n171), .A (CLOCK_slh__n170));
CLKBUF_X1 CLOCK_slh__c117 (.Z (n_17), .A (CLOCK_slh__n171));
CLKBUF_X1 CLOCK_slh__c121 (.Z (CLOCK_slh__n176), .A (CLOCK_slh__n175));
CLKBUF_X1 CLOCK_slh__c122 (.Z (CLOCK_slh__n177), .A (CLOCK_slh__n176));
CLKBUF_X1 CLOCK_slh__c123 (.Z (n_32), .A (CLOCK_slh__n177));
CLKBUF_X1 CLOCK_slh__c127 (.Z (CLOCK_slh__n182), .A (CLOCK_slh__n181));
CLKBUF_X1 CLOCK_slh__c128 (.Z (CLOCK_slh__n183), .A (CLOCK_slh__n182));
CLKBUF_X1 CLOCK_slh__c129 (.Z (n_4), .A (CLOCK_slh__n183));
CLKBUF_X1 CLOCK_slh__c133 (.Z (CLOCK_slh__n188), .A (CLOCK_slh__n187));
CLKBUF_X1 CLOCK_slh__c134 (.Z (CLOCK_slh__n189), .A (CLOCK_slh__n188));
CLKBUF_X1 CLOCK_slh__c135 (.Z (n_16), .A (CLOCK_slh__n189));
CLKBUF_X1 CLOCK_slh__c139 (.Z (CLOCK_slh__n194), .A (CLOCK_slh__n193));
CLKBUF_X1 CLOCK_slh__c140 (.Z (CLOCK_slh__n195), .A (CLOCK_slh__n194));
CLKBUF_X1 CLOCK_slh__c141 (.Z (n_22), .A (CLOCK_slh__n195));
CLKBUF_X1 CLOCK_slh__c145 (.Z (CLOCK_slh__n200), .A (CLOCK_slh__n199));
CLKBUF_X1 CLOCK_slh__c146 (.Z (CLOCK_slh__n201), .A (CLOCK_slh__n200));
CLKBUF_X1 CLOCK_slh__c147 (.Z (n_25), .A (CLOCK_slh__n201));
CLKBUF_X1 CLOCK_slh__c151 (.Z (CLOCK_slh__n206), .A (CLOCK_slh__n205));
CLKBUF_X1 CLOCK_slh__c152 (.Z (CLOCK_slh__n207), .A (CLOCK_slh__n206));
CLKBUF_X1 CLOCK_slh__c153 (.Z (n_23), .A (CLOCK_slh__n207));
CLKBUF_X1 CLOCK_slh__c157 (.Z (CLOCK_slh__n212), .A (CLOCK_slh__n211));
CLKBUF_X1 CLOCK_slh__c158 (.Z (CLOCK_slh__n213), .A (CLOCK_slh__n212));
CLKBUF_X1 CLOCK_slh__c159 (.Z (n_24), .A (CLOCK_slh__n213));
CLKBUF_X1 CLOCK_slh__c163 (.Z (CLOCK_slh__n218), .A (CLOCK_slh__n217));
CLKBUF_X1 CLOCK_slh__c164 (.Z (CLOCK_slh__n219), .A (CLOCK_slh__n218));
CLKBUF_X1 CLOCK_slh__c165 (.Z (n_28), .A (CLOCK_slh__n219));
CLKBUF_X1 CLOCK_slh__c169 (.Z (CLOCK_slh__n224), .A (CLOCK_slh__n223));
CLKBUF_X1 CLOCK_slh__c170 (.Z (CLOCK_slh__n225), .A (CLOCK_slh__n224));
CLKBUF_X1 CLOCK_slh__c171 (.Z (CLOCK_sph__n244), .A (CLOCK_slh__n225));
CLKBUF_X1 CLOCK_slh__c175 (.Z (CLOCK_slh__n230), .A (CLOCK_slh__n229));
CLKBUF_X1 CLOCK_slh__c176 (.Z (CLOCK_slh__n231), .A (CLOCK_slh__n230));
CLKBUF_X1 CLOCK_slh__c177 (.Z (n_29), .A (CLOCK_slh__n231));
CLKBUF_X1 CLOCK_slh__c181 (.Z (CLOCK_slh__n236), .A (CLOCK_slh__n235));
CLKBUF_X1 CLOCK_slh__c182 (.Z (CLOCK_slh__n237), .A (CLOCK_slh__n236));
CLKBUF_X1 CLOCK_slh__c183 (.Z (n_31), .A (CLOCK_slh__n237));
CLKBUF_X1 CLOCK_slh__c184 (.Z (CLOCK_slh__n239), .A (CLOCK_slh__n238));
CLKBUF_X1 CLOCK_slh__c185 (.Z (CLOCK_slh__n240), .A (CLOCK_slh__n239));
CLKBUF_X1 CLOCK_slh__c186 (.Z (n_30), .A (CLOCK_slh__n240));
CLKBUF_X1 CLOCK_slh__c187 (.Z (CLOCK_slh__n242), .A (CLOCK_slh__n241));
CLKBUF_X1 CLOCK_slh__c188 (.Z (CLOCK_slh__n243), .A (CLOCK_slh__n242));
CLKBUF_X1 CLOCK_slh__c189 (.Z (n_15), .A (CLOCK_slh__n243));
CLKBUF_X1 CLOCK_sph__c190 (.Z (n_33), .A (CLOCK_sph__n244));

endmodule //buffer__0_18

module datapath__0_10 (p_0, finalResult, p_1);

output [63:0] p_1;
input [63:0] finalResult;
input [63:0] p_0;
wire n_0;
wire n_366;
wire n_1;
wire n_365;
wire n_364;
wire n_2;
wire n_369;
wire n_363;
wire n_3;
wire n_370;
wire n_376;
wire n_372;
wire n_361;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_358;
wire n_349;
wire n_11;
wire n_5;
wire n_359;
wire n_353;
wire n_8;
wire n_356;
wire n_354;
wire n_360;
wire n_351;
wire n_347;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_344;
wire n_335;
wire n_19;
wire n_13;
wire n_345;
wire n_339;
wire n_16;
wire n_342;
wire n_340;
wire n_346;
wire n_337;
wire n_333;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_330;
wire n_321;
wire n_27;
wire n_21;
wire n_331;
wire n_325;
wire n_24;
wire n_328;
wire n_326;
wire n_332;
wire n_323;
wire n_319;
wire n_34;
wire n_33;
wire n_30;
wire n_31;
wire n_28;
wire n_285;
wire n_275;
wire n_35;
wire n_29;
wire n_284;
wire n_287;
wire n_277;
wire n_32;
wire n_286;
wire n_282;
wire n_279;
wire n_289;
wire n_63;
wire n_42;
wire n_41;
wire n_38;
wire n_39;
wire n_36;
wire n_313;
wire n_257;
wire n_43;
wire n_37;
wire n_312;
wire n_315;
wire n_259;
wire n_40;
wire n_314;
wire n_318;
wire n_261;
wire n_317;
wire n_61;
wire n_50;
wire n_49;
wire n_46;
wire n_47;
wire n_44;
wire n_296;
wire n_269;
wire n_51;
wire n_45;
wire n_295;
wire n_298;
wire n_271;
wire n_48;
wire n_297;
wire n_293;
wire n_273;
wire n_300;
wire n_59;
wire n_58;
wire n_57;
wire n_54;
wire n_55;
wire n_52;
wire n_305;
wire n_263;
wire n_65;
wire n_53;
wire n_304;
wire n_307;
wire n_266;
wire n_56;
wire n_306;
wire n_302;
wire n_267;
wire n_60;
wire n_268;
wire n_292;
wire n_62;
wire n_256;
wire n_310;
wire n_64;
wire n_274;
wire n_281;
wire n_308;
wire n_377;
wire n_373;
wire n_254;
wire n_72;
wire n_71;
wire n_68;
wire n_69;
wire n_66;
wire n_223;
wire n_213;
wire n_73;
wire n_67;
wire n_222;
wire n_225;
wire n_215;
wire n_70;
wire n_224;
wire n_220;
wire n_217;
wire n_227;
wire n_101;
wire n_80;
wire n_79;
wire n_76;
wire n_77;
wire n_74;
wire n_248;
wire n_206;
wire n_81;
wire n_75;
wire n_247;
wire n_250;
wire n_208;
wire n_78;
wire n_249;
wire n_253;
wire n_210;
wire n_252;
wire n_99;
wire n_88;
wire n_87;
wire n_84;
wire n_85;
wire n_82;
wire n_234;
wire n_192;
wire n_89;
wire n_83;
wire n_233;
wire n_236;
wire n_194;
wire n_86;
wire n_235;
wire n_231;
wire n_196;
wire n_238;
wire n_98;
wire n_97;
wire n_95;
wire n_94;
wire n_91;
wire n_90;
wire n_202;
wire n_242;
wire n_199;
wire n_103;
wire n_92;
wire n_93;
wire n_241;
wire n_200;
wire n_96;
wire n_243;
wire n_203;
wire n_204;
wire n_191;
wire n_230;
wire n_100;
wire n_205;
wire n_245;
wire n_102;
wire n_212;
wire n_219;
wire n_244;
wire n_189;
wire n_110;
wire n_109;
wire n_106;
wire n_107;
wire n_104;
wire n_186;
wire n_177;
wire n_111;
wire n_105;
wire n_187;
wire n_181;
wire n_108;
wire n_184;
wire n_182;
wire n_188;
wire n_179;
wire n_175;
wire n_118;
wire n_117;
wire n_114;
wire n_115;
wire n_112;
wire n_164;
wire n_154;
wire n_119;
wire n_113;
wire n_163;
wire n_166;
wire n_156;
wire n_116;
wire n_165;
wire n_161;
wire n_158;
wire n_168;
wire n_128;
wire n_127;
wire n_125;
wire n_124;
wire n_121;
wire n_120;
wire n_149;
wire n_172;
wire n_145;
wire n_129;
wire n_122;
wire n_123;
wire n_171;
wire n_146;
wire n_126;
wire n_173;
wire n_150;
wire n_151;
wire n_153;
wire n_160;
wire n_174;
wire n_143;
wire n_142;
wire n_140;
wire n_136;
wire n_141;
wire n_135;
wire n_137;
wire n_379;
wire n_375;
wire n_170;
wire n_148;
wire n_155;
wire n_167;
wire n_162;
wire n_157;
wire n_178;
wire n_195;
wire n_209;
wire n_216;
wire n_232;
wire n_246;
wire n_311;
wire n_260;
wire n_258;
wire n_264;
wire n_265;
wire n_294;
wire n_272;
wire n_270;
wire n_283;
wire n_278;
wire n_276;
wire n_288;
wire n_299;
wire n_316;
wire n_322;
wire n_320;
wire n_329;
wire n_324;
wire n_327;
wire n_334;
wire n_338;
wire n_341;
wire n_336;
wire n_343;
wire n_348;
wire n_352;
wire n_355;
wire n_350;
wire n_357;
wire n_362;
wire n_368;
wire n_367;
wire n_374;
wire n_378;
wire n_412;
wire n_228;
wire n_479;
wire n_130;
wire n_478;
wire n_229;
wire n_240;
wire n_131;
wire n_371;
wire n_290;
wire n_301;
wire n_132;
wire n_415;
wire n_405;
wire n_385;
wire n_133;
wire n_421;
wire n_417;
wire n_406;
wire n_396;
wire n_472;
wire n_394;
wire n_400;
wire n_410;
wire n_420;
wire n_431;
wire n_432;
wire n_434;
wire n_440;
wire n_447;
wire n_134;
wire n_144;
wire n_138;
wire n_139;
wire n_180;
wire n_169;
wire n_147;
wire n_176;
wire n_159;
wire n_152;
wire n_211;
wire n_226;
wire n_183;
wire n_190;
wire n_197;
wire n_185;
wire n_207;
wire n_214;
wire n_201;
wire n_193;
wire n_198;
wire n_221;
wire n_218;
wire n_237;
wire n_280;
wire n_239;
wire n_251;
wire n_255;
wire n_262;
wire n_291;
wire n_303;
wire n_382;
wire n_309;
wire n_380;
wire n_384;
wire n_414;
wire n_381;
wire n_383;
wire n_386;
wire n_395;
wire n_387;
wire n_388;
wire n_389;
wire n_468;
wire n_392;
wire n_390;
wire n_391;
wire n_469;
wire n_393;
wire n_465;
wire n_397;
wire n_403;
wire n_398;
wire n_399;
wire n_402;
wire n_401;
wire n_404;
wire n_477;
wire n_411;
wire n_407;
wire n_408;
wire n_409;
wire n_413;
wire n_476;
wire n_416;
wire n_418;
wire n_419;
wire n_459;
wire n_457;
wire n_422;
wire n_423;
wire n_441;
wire n_433;
wire n_424;
wire n_446;
wire n_453;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_430;
wire n_429;
wire n_436;
wire n_439;
wire n_438;
wire n_437;
wire n_442;
wire n_443;
wire n_456;
wire n_455;
wire n_445;
wire n_449;
wire n_452;
wire n_451;
wire n_450;
wire n_454;
wire n_464;
wire n_458;
wire n_461;
wire n_460;
wire n_463;
wire n_462;
wire n_466;
wire n_467;
wire n_475;
wire n_471;
wire n_470;
wire n_474;
wire n_473;


NAND2_X1 i_543 (.ZN (n_479), .A1 (p_0[60]), .A2 (finalResult[60]));
OR2_X1 i_542 (.ZN (n_478), .A1 (p_0[60]), .A2 (finalResult[60]));
INV_X1 i_541 (.ZN (n_477), .A (n_230));
INV_X1 i_540 (.ZN (n_476), .A (n_245));
OR2_X1 i_539 (.ZN (n_475), .A1 (p_0[44]), .A2 (finalResult[44]));
INV_X1 i_538 (.ZN (n_474), .A (p_0[45]));
INV_X1 i_537 (.ZN (n_473), .A (finalResult[45]));
NAND2_X1 i_536 (.ZN (n_472), .A1 (n_474), .A2 (n_473));
INV_X1 i_535 (.ZN (n_471), .A (p_0[47]));
INV_X1 i_534 (.ZN (n_470), .A (finalResult[47]));
NAND2_X1 i_533 (.ZN (n_469), .A1 (n_471), .A2 (n_470));
OAI211_X1 i_532 (.ZN (n_468), .A (n_469), .B (n_472), .C1 (p_0[46]), .C2 (finalResult[46]));
INV_X1 i_531 (.ZN (n_467), .A (n_468));
NAND2_X1 i_530 (.ZN (n_466), .A1 (n_467), .A2 (n_475));
INV_X1 i_529 (.ZN (n_465), .A (n_466));
INV_X1 i_528 (.ZN (n_464), .A (n_220));
INV_X1 i_527 (.ZN (n_463), .A (p_0[33]));
INV_X1 i_526 (.ZN (n_462), .A (finalResult[33]));
NAND2_X1 i_525 (.ZN (n_224), .A1 (n_463), .A2 (n_462));
INV_X1 i_524 (.ZN (n_461), .A (p_0[35]));
INV_X1 i_523 (.ZN (n_460), .A (finalResult[35]));
NAND2_X1 i_522 (.ZN (n_459), .A1 (n_461), .A2 (n_460));
NOR2_X1 i_521 (.ZN (n_223), .A1 (p_0[34]), .A2 (finalResult[34]));
INV_X1 i_520 (.ZN (n_222), .A (n_223));
NAND3_X1 i_519 (.ZN (n_458), .A1 (n_222), .A2 (n_224), .A3 (n_459));
INV_X1 i_518 (.ZN (n_457), .A (n_458));
NAND2_X1 i_517 (.ZN (n_219), .A1 (n_457), .A2 (n_464));
NOR2_X1 i_516 (.ZN (n_456), .A1 (p_0[31]), .A2 (finalResult[31]));
INV_X1 i_515 (.ZN (n_308), .A (n_456));
NOR2_X1 i_514 (.ZN (n_455), .A1 (n_305), .A2 (n_307));
OAI21_X1 i_513 (.ZN (n_454), .A (n_455), .B1 (p_0[28]), .B2 (finalResult[28]));
INV_X1 i_512 (.ZN (n_453), .A (n_454));
INV_X1 i_511 (.ZN (n_452), .A (p_0[27]));
INV_X1 i_510 (.ZN (n_451), .A (finalResult[27]));
INV_X1 i_509 (.ZN (n_450), .A (n_269));
INV_X1 i_508 (.ZN (n_449), .A (n_270));
OAI221_X1 i_506 (.ZN (n_447), .A (n_449), .B1 (n_452), .B2 (n_451), .C1 (n_450), .C2 (n_300));
NAND3_X1 i_505 (.ZN (n_446), .A1 (n_453), .A2 (n_308), .A3 (n_447));
INV_X1 i_504 (.ZN (n_445), .A (n_265));
AOI21_X1 i_502 (.ZN (n_443), .A (n_263), .B1 (n_455), .B2 (n_445));
OAI22_X1 i_501 (.ZN (n_442), .A1 (n_443), .A2 (n_456), .B1 (n_377), .B2 (n_373));
INV_X1 i_500 (.ZN (n_441), .A (n_442));
NOR2_X1 i_499 (.ZN (n_440), .A1 (n_294), .A2 (n_293));
INV_X1 i_498 (.ZN (n_439), .A (p_0[23]));
INV_X1 i_497 (.ZN (n_438), .A (finalResult[23]));
INV_X1 i_496 (.ZN (n_437), .A (n_257));
INV_X1 i_495 (.ZN (n_436), .A (n_258));
OAI221_X1 i_493 (.ZN (n_434), .A (n_436), .B1 (n_439), .B2 (n_438), .C1 (n_437), .C2 (n_317));
NAND4_X1 i_492 (.ZN (n_433), .A1 (n_453), .A2 (n_308), .A3 (n_440), .A4 (n_434));
INV_X1 i_491 (.ZN (n_432), .A (n_318));
INV_X1 i_490 (.ZN (n_431), .A (n_311));
OR2_X1 i_489 (.ZN (n_281), .A1 (n_283), .A2 (n_282));
NOR4_X4 i_488 (.ZN (n_319), .A1 (n_327), .A2 (n_323), .A3 (n_320), .A4 (n_324));
INV_X1 i_487 (.ZN (n_430), .A (n_276));
AOI22_X1 i_486 (.ZN (n_429), .A1 (n_288), .A2 (n_275), .B1 (p_0[19]), .B2 (finalResult[19]));
NAND2_X1 i_485 (.ZN (n_428), .A1 (n_430), .A2 (n_429));
INV_X1 i_484 (.ZN (n_274), .A (n_428));
OAI21_X2 i_483 (.ZN (n_427), .A (n_274), .B1 (n_319), .B2 (n_281));
NAND3_X1 i_482 (.ZN (n_426), .A1 (n_431), .A2 (n_432), .A3 (n_427));
INV_X2 i_481 (.ZN (n_425), .A (n_426));
NAND4_X1 i_480 (.ZN (n_424), .A1 (n_453), .A2 (n_308), .A3 (n_440), .A4 (n_425));
NAND4_X1 i_479 (.ZN (n_423), .A1 (n_441), .A2 (n_433), .A3 (n_424), .A4 (n_446));
INV_X1 i_478 (.ZN (n_254), .A (n_423));
NAND2_X1 i_477 (.ZN (n_217), .A1 (p_0[32]), .A2 (finalResult[32]));
NAND2_X1 i_476 (.ZN (n_216), .A1 (p_0[33]), .A2 (finalResult[33]));
NAND2_X1 i_475 (.ZN (n_422), .A1 (n_217), .A2 (n_216));
NAND2_X1 i_474 (.ZN (n_421), .A1 (n_457), .A2 (n_422));
INV_X1 i_473 (.ZN (n_227), .A (n_459));
NAND2_X1 i_472 (.ZN (n_420), .A1 (p_0[34]), .A2 (finalResult[34]));
NAND2_X1 i_471 (.ZN (n_419), .A1 (p_0[35]), .A2 (finalResult[35]));
OAI21_X1 i_470 (.ZN (n_418), .A (n_419), .B1 (n_227), .B2 (n_420));
INV_X1 i_469 (.ZN (n_417), .A (n_418));
OAI211_X1 i_468 (.ZN (n_416), .A (n_421), .B (n_417), .C1 (n_219), .C2 (n_254));
NAND4_X1 i_467 (.ZN (n_415), .A1 (n_476), .A2 (n_477), .A3 (n_465), .A4 (n_416));
INV_X1 i_466 (.ZN (n_414), .A (n_415));
NAND2_X1 i_465 (.ZN (n_210), .A1 (p_0[36]), .A2 (finalResult[36]));
NAND2_X1 i_464 (.ZN (n_209), .A1 (p_0[37]), .A2 (finalResult[37]));
NAND2_X1 i_463 (.ZN (n_413), .A1 (n_210), .A2 (n_209));
NOR2_X1 i_462 (.ZN (n_252), .A1 (p_0[39]), .A2 (finalResult[39]));
INV_X1 i_461 (.ZN (n_412), .A (n_252));
NOR2_X1 i_460 (.ZN (n_250), .A1 (p_0[37]), .A2 (finalResult[37]));
INV_X1 i_459 (.ZN (n_249), .A (n_250));
NOR2_X1 i_458 (.ZN (n_248), .A1 (p_0[38]), .A2 (finalResult[38]));
INV_X1 i_457 (.ZN (n_247), .A (n_248));
NAND4_X1 i_456 (.ZN (n_411), .A1 (n_413), .A2 (n_412), .A3 (n_247), .A4 (n_249));
NAND2_X1 i_455 (.ZN (n_410), .A1 (p_0[38]), .A2 (finalResult[38]));
NAND2_X1 i_454 (.ZN (n_409), .A1 (p_0[39]), .A2 (finalResult[39]));
OAI21_X1 i_453 (.ZN (n_408), .A (n_409), .B1 (n_252), .B2 (n_410));
INV_X1 i_452 (.ZN (n_407), .A (n_408));
NAND2_X1 i_451 (.ZN (n_406), .A1 (n_411), .A2 (n_407));
NAND3_X1 i_450 (.ZN (n_405), .A1 (n_477), .A2 (n_465), .A3 (n_406));
NAND2_X1 i_449 (.ZN (n_196), .A1 (p_0[40]), .A2 (finalResult[40]));
NAND2_X1 i_448 (.ZN (n_195), .A1 (p_0[41]), .A2 (finalResult[41]));
NAND2_X1 i_447 (.ZN (n_404), .A1 (n_196), .A2 (n_195));
INV_X1 i_446 (.ZN (n_403), .A (n_404));
INV_X1 i_445 (.ZN (n_402), .A (p_0[41]));
INV_X1 i_444 (.ZN (n_401), .A (finalResult[41]));
NAND2_X1 i_435 (.ZN (n_235), .A1 (n_402), .A2 (n_401));
NOR2_X1 i_383 (.ZN (n_234), .A1 (p_0[42]), .A2 (finalResult[42]));
INV_X1 i_374 (.ZN (n_233), .A (n_234));
OAI211_X1 i_373 (.ZN (n_232), .A (n_233), .B (n_235), .C1 (p_0[43]), .C2 (finalResult[43]));
NOR2_X1 i_372 (.ZN (n_238), .A1 (p_0[43]), .A2 (finalResult[43]));
NAND2_X1 i_370 (.ZN (n_400), .A1 (p_0[42]), .A2 (finalResult[42]));
NAND2_X1 i_368 (.ZN (n_399), .A1 (p_0[43]), .A2 (finalResult[43]));
OAI21_X1 i_367 (.ZN (n_398), .A (n_399), .B1 (n_238), .B2 (n_400));
INV_X1 i_366 (.ZN (n_397), .A (n_398));
OAI21_X1 i_365 (.ZN (n_396), .A (n_397), .B1 (n_232), .B2 (n_403));
NAND2_X1 i_356 (.ZN (n_395), .A1 (n_465), .A2 (n_396));
NAND2_X1 i_355 (.ZN (n_394), .A1 (p_0[45]), .A2 (finalResult[45]));
NAND2_X1 i_354 (.ZN (n_393), .A1 (n_204), .A2 (n_394));
INV_X1 i_345 (.ZN (n_392), .A (n_393));
INV_X1 i_344 (.ZN (n_244), .A (n_469));
NAND2_X1 i_338 (.ZN (n_200), .A1 (p_0[46]), .A2 (finalResult[46]));
NAND2_X1 i_332 (.ZN (n_391), .A1 (p_0[47]), .A2 (finalResult[47]));
OAI21_X1 i_326 (.ZN (n_390), .A (n_391), .B1 (n_244), .B2 (n_200));
INV_X1 i_320 (.ZN (n_389), .A (n_390));
OAI21_X1 i_319 (.ZN (n_388), .A (n_389), .B1 (n_468), .B2 (n_392));
INV_X1 i_318 (.ZN (n_387), .A (n_388));
NAND2_X1 i_316 (.ZN (n_386), .A1 (n_395), .A2 (n_387));
INV_X1 i_315 (.ZN (n_385), .A (n_386));
NAND2_X1 i_314 (.ZN (n_384), .A1 (n_405), .A2 (n_385));
OR3_X1 i_313 (.ZN (n_383), .A1 (n_187), .A2 (n_188), .A3 (n_186));
INV_X1 i_312 (.ZN (n_382), .A (n_383));
OAI21_X1 i_311 (.ZN (n_381), .A (n_382), .B1 (p_0[48]), .B2 (finalResult[48]));
INV_X1 i_310 (.ZN (n_380), .A (n_381));
OAI21_X1 i_308 (.ZN (n_371), .A (n_380), .B1 (n_384), .B2 (n_414));
NAND2_X1 i_307 (.ZN (n_309), .A1 (n_182), .A2 (n_181));
NAND2_X1 i_306 (.ZN (n_303), .A1 (n_382), .A2 (n_309));
NAND2_X1 i_304 (.ZN (n_301), .A1 (p_0[51]), .A2 (finalResult[51]));
OAI211_X1 i_303 (.ZN (n_291), .A (n_303), .B (n_301), .C1 (n_188), .C2 (n_178));
INV_X1 i_302 (.ZN (n_290), .A (n_291));
OAI21_X1 i_301 (.ZN (n_280), .A (n_170), .B1 (p_0[56]), .B2 (finalResult[56]));
INV_X1 i_300 (.ZN (n_262), .A (n_161));
INV_X1 i_299 (.ZN (n_255), .A (n_162));
NAND2_X1 i_298 (.ZN (n_160), .A1 (n_255), .A2 (n_262));
OR2_X1 i_297 (.ZN (n_251), .A1 (n_160), .A2 (n_280));
AOI21_X1 i_296 (.ZN (n_240), .A (n_251), .B1 (n_371), .B2 (n_290));
OAI221_X1 i_293 (.ZN (n_239), .A (n_148), .B1 (n_146), .B2 (n_174), .C1 (n_378), .C2 (n_374));
INV_X1 i_292 (.ZN (n_237), .A (n_239));
OAI21_X1 i_291 (.ZN (n_229), .A (n_237), .B1 (n_153), .B2 (n_280));
OAI21_X1 i_290 (.ZN (n_228), .A (n_478), .B1 (n_229), .B2 (n_240));
NAND2_X1 i_289 (.ZN (n_226), .A1 (p_0[62]), .A2 (finalResult[62]));
INV_X1 i_288 (.ZN (n_221), .A (n_226));
NOR2_X1 i_287 (.ZN (n_218), .A1 (n_136), .A2 (n_221));
NAND3_X1 i_286 (.ZN (n_214), .A1 (n_228), .A2 (n_479), .A3 (n_218));
OR2_X1 i_285 (.ZN (n_211), .A1 (p_0[62]), .A2 (finalResult[62]));
NAND2_X1 i_283 (.ZN (n_137), .A1 (n_379), .A2 (n_375));
OAI21_X1 i_282 (.ZN (n_207), .A (n_211), .B1 (n_137), .B2 (n_221));
INV_X1 i_281 (.ZN (n_201), .A (n_207));
INV_X1 i_280 (.ZN (n_198), .A (finalResult[63]));
XNOR2_X1 i_278 (.ZN (n_197), .A (p_0[63]), .B (n_198));
INV_X1 i_277 (.ZN (n_193), .A (n_197));
NAND3_X1 i_276 (.ZN (n_190), .A1 (n_214), .A2 (n_201), .A3 (n_193));
INV_X1 i_275 (.ZN (n_185), .A (n_214));
OAI21_X1 i_274 (.ZN (n_183), .A (n_197), .B1 (n_185), .B2 (n_207));
NAND2_X1 i_273 (.ZN (p_1[63]), .A1 (n_183), .A2 (n_190));
NAND2_X1 i_271 (.ZN (n_180), .A1 (n_211), .A2 (n_226));
INV_X1 i_270 (.ZN (n_176), .A (n_180));
NAND2_X1 i_269 (.ZN (n_169), .A1 (p_0[61]), .A2 (finalResult[61]));
INV_X1 i_267 (.ZN (n_159), .A (n_169));
INV_X1 i_266 (.ZN (n_152), .A (n_137));
AOI21_X1 i_265 (.ZN (n_147), .A (n_152), .B1 (n_228), .B2 (n_479));
OAI21_X1 i_264 (.ZN (n_144), .A (n_176), .B1 (n_147), .B2 (n_159));
INV_X1 i_262 (.ZN (n_139), .A (n_147));
NAND3_X1 i_261 (.ZN (n_138), .A1 (n_139), .A2 (n_180), .A3 (n_169));
NAND2_X1 i_260 (.ZN (n_134), .A1 (n_144), .A2 (n_138));
INV_X1 i_259 (.ZN (p_1[62]), .A (n_134));
INV_X1 i_257 (.ZN (n_304), .A (n_305));
INV_X1 i_256 (.ZN (n_306), .A (n_307));
NOR2_X1 i_255 (.ZN (n_302), .A1 (p_0[28]), .A2 (finalResult[28]));
INV_X1 i_254 (.ZN (n_268), .A (n_447));
INV_X1 i_253 (.ZN (n_292), .A (n_440));
INV_X1 i_249 (.ZN (n_256), .A (n_434));
NAND2_X1 i_248 (.ZN (n_310), .A1 (n_431), .A2 (n_432));
INV_X1 i_247 (.ZN (n_213), .A (n_420));
INV_X1 i_244 (.ZN (n_225), .A (n_224));
INV_X1 i_243 (.ZN (n_206), .A (n_410));
INV_X1 i_240 (.ZN (n_192), .A (n_400));
INV_X1 i_239 (.ZN (n_236), .A (n_235));
INV_X1 i_233 (.ZN (n_202), .A (n_394));
NOR2_X1 i_224 (.ZN (n_242), .A1 (p_0[46]), .A2 (finalResult[46]));
INV_X1 i_223 (.ZN (n_243), .A (n_472));
INV_X1 i_216 (.ZN (n_203), .A (n_204));
INV_X1 i_211 (.ZN (n_191), .A (n_396));
INV_X1 i_208 (.ZN (n_205), .A (n_406));
NAND2_X1 i_207 (.ZN (n_133), .A1 (n_421), .A2 (n_417));
INV_X1 i_206 (.ZN (n_212), .A (n_133));
NAND3_X1 i_205 (.ZN (n_132), .A1 (n_415), .A2 (n_405), .A3 (n_385));
INV_X1 i_204 (.ZN (n_189), .A (n_132));
NOR2_X1 i_203 (.ZN (n_184), .A1 (p_0[48]), .A2 (finalResult[48]));
INV_X1 i_202 (.ZN (n_179), .A (n_301));
NAND2_X1 i_201 (.ZN (n_131), .A1 (n_371), .A2 (n_290));
INV_X1 i_199 (.ZN (n_175), .A (n_131));
NOR2_X1 i_198 (.ZN (n_143), .A1 (n_229), .A2 (n_240));
NAND2_X1 i_197 (.ZN (n_130), .A1 (n_478), .A2 (n_479));
INV_X1 i_196 (.ZN (n_142), .A (n_130));
NAND2_X1 i_195 (.ZN (n_141), .A1 (n_228), .A2 (n_479));
INV_X1 i_194 (.ZN (n_140), .A (n_141));
INV_X1 i_193 (.ZN (n_135), .A (n_136));
NAND3_X1 i_192 (.ZN (n_246), .A1 (n_412), .A2 (n_247), .A3 (n_249));
INV_X1 i_443 (.ZN (n_379), .A (p_0[61]));
INV_X1 i_442 (.ZN (n_378), .A (p_0[59]));
INV_X1 i_441 (.ZN (n_377), .A (p_0[31]));
INV_X1 i_440 (.ZN (n_376), .A (p_0[3]));
INV_X1 i_439 (.ZN (n_375), .A (finalResult[61]));
INV_X1 i_438 (.ZN (n_374), .A (finalResult[59]));
INV_X1 i_437 (.ZN (n_373), .A (finalResult[31]));
INV_X1 i_436 (.ZN (n_372), .A (finalResult[3]));
NAND2_X1 i_434 (.ZN (n_370), .A1 (n_376), .A2 (n_372));
NAND2_X1 i_433 (.ZN (n_369), .A1 (p_0[2]), .A2 (finalResult[2]));
INV_X1 i_432 (.ZN (n_368), .A (n_369));
NOR2_X1 i_431 (.ZN (n_367), .A1 (p_0[1]), .A2 (finalResult[1]));
NAND2_X1 i_430 (.ZN (n_366), .A1 (p_0[0]), .A2 (finalResult[0]));
NAND2_X1 i_429 (.ZN (n_365), .A1 (p_0[1]), .A2 (finalResult[1]));
AOI21_X1 i_428 (.ZN (n_364), .A (n_367), .B1 (n_366), .B2 (n_365));
OAI22_X2 i_427 (.ZN (n_363), .A1 (p_0[2]), .A2 (finalResult[2]), .B1 (n_368), .B2 (n_364));
OAI21_X1 i_426 (.ZN (n_362), .A (n_363), .B1 (n_376), .B2 (n_372));
NAND2_X2 i_425 (.ZN (n_361), .A1 (n_370), .A2 (n_362));
NOR2_X2 i_424 (.ZN (n_360), .A1 (p_0[7]), .A2 (finalResult[7]));
NOR2_X2 i_423 (.ZN (n_359), .A1 (p_0[5]), .A2 (finalResult[5]));
NOR2_X1 i_422 (.ZN (n_358), .A1 (p_0[6]), .A2 (finalResult[6]));
OR3_X2 i_421 (.ZN (n_357), .A1 (n_360), .A2 (n_358), .A3 (n_359));
NOR2_X1 i_420 (.ZN (n_356), .A1 (p_0[4]), .A2 (finalResult[4]));
NOR3_X2 i_419 (.ZN (n_355), .A1 (n_357), .A2 (n_356), .A3 (n_361));
NAND2_X1 i_418 (.ZN (n_354), .A1 (p_0[4]), .A2 (finalResult[4]));
NAND2_X1 i_417 (.ZN (n_353), .A1 (p_0[5]), .A2 (finalResult[5]));
AOI21_X2 i_416 (.ZN (n_352), .A (n_357), .B1 (n_354), .B2 (n_353));
AND2_X1 i_415 (.ZN (n_351), .A1 (p_0[7]), .A2 (finalResult[7]));
NAND2_X1 i_414 (.ZN (n_350), .A1 (p_0[6]), .A2 (finalResult[6]));
INV_X1 i_413 (.ZN (n_349), .A (n_350));
NOR2_X1 i_412 (.ZN (n_348), .A1 (n_360), .A2 (n_350));
NOR4_X4 i_411 (.ZN (n_347), .A1 (n_351), .A2 (n_348), .A3 (n_352), .A4 (n_355));
NOR2_X1 i_410 (.ZN (n_346), .A1 (p_0[11]), .A2 (finalResult[11]));
NOR2_X1 i_409 (.ZN (n_345), .A1 (p_0[9]), .A2 (finalResult[9]));
NOR2_X1 i_408 (.ZN (n_344), .A1 (p_0[10]), .A2 (finalResult[10]));
OR3_X1 i_407 (.ZN (n_343), .A1 (n_346), .A2 (n_344), .A3 (n_345));
NOR2_X1 i_406 (.ZN (n_342), .A1 (p_0[8]), .A2 (finalResult[8]));
NOR3_X2 i_405 (.ZN (n_341), .A1 (n_343), .A2 (n_342), .A3 (n_347));
NAND2_X1 i_404 (.ZN (n_340), .A1 (p_0[8]), .A2 (finalResult[8]));
NAND2_X1 i_403 (.ZN (n_339), .A1 (p_0[9]), .A2 (finalResult[9]));
AOI21_X1 i_402 (.ZN (n_338), .A (n_343), .B1 (n_340), .B2 (n_339));
AND2_X1 i_401 (.ZN (n_337), .A1 (p_0[11]), .A2 (finalResult[11]));
NAND2_X1 i_400 (.ZN (n_336), .A1 (p_0[10]), .A2 (finalResult[10]));
INV_X1 i_399 (.ZN (n_335), .A (n_336));
NOR2_X1 i_398 (.ZN (n_334), .A1 (n_346), .A2 (n_336));
NOR4_X4 i_397 (.ZN (n_333), .A1 (n_337), .A2 (n_334), .A3 (n_338), .A4 (n_341));
NOR2_X1 i_396 (.ZN (n_332), .A1 (p_0[15]), .A2 (finalResult[15]));
NOR2_X1 i_395 (.ZN (n_331), .A1 (p_0[13]), .A2 (finalResult[13]));
NOR2_X1 i_394 (.ZN (n_330), .A1 (p_0[14]), .A2 (finalResult[14]));
OR3_X1 i_393 (.ZN (n_329), .A1 (n_332), .A2 (n_330), .A3 (n_331));
NOR2_X1 i_392 (.ZN (n_328), .A1 (p_0[12]), .A2 (finalResult[12]));
NOR3_X1 i_391 (.ZN (n_327), .A1 (n_329), .A2 (n_328), .A3 (n_333));
NAND2_X1 i_390 (.ZN (n_326), .A1 (p_0[12]), .A2 (finalResult[12]));
NAND2_X1 i_389 (.ZN (n_325), .A1 (p_0[13]), .A2 (finalResult[13]));
AOI21_X1 i_388 (.ZN (n_324), .A (n_329), .B1 (n_326), .B2 (n_325));
AND2_X1 i_387 (.ZN (n_323), .A1 (p_0[15]), .A2 (finalResult[15]));
NAND2_X1 i_386 (.ZN (n_322), .A1 (p_0[14]), .A2 (finalResult[14]));
INV_X1 i_385 (.ZN (n_321), .A (n_322));
NOR2_X1 i_384 (.ZN (n_320), .A1 (n_332), .A2 (n_322));
NOR2_X1 i_382 (.ZN (n_318), .A1 (p_0[20]), .A2 (finalResult[20]));
NOR2_X1 i_381 (.ZN (n_317), .A1 (p_0[23]), .A2 (finalResult[23]));
INV_X1 i_380 (.ZN (n_316), .A (n_317));
NOR2_X1 i_379 (.ZN (n_315), .A1 (p_0[21]), .A2 (finalResult[21]));
INV_X1 i_378 (.ZN (n_314), .A (n_315));
NOR2_X1 i_377 (.ZN (n_313), .A1 (p_0[22]), .A2 (finalResult[22]));
INV_X1 i_376 (.ZN (n_312), .A (n_313));
NAND3_X1 i_375 (.ZN (n_311), .A1 (n_316), .A2 (n_312), .A3 (n_314));
NOR2_X1 i_371 (.ZN (n_307), .A1 (p_0[29]), .A2 (finalResult[29]));
NOR2_X1 i_369 (.ZN (n_305), .A1 (p_0[30]), .A2 (finalResult[30]));
NOR2_X1 i_364 (.ZN (n_300), .A1 (p_0[27]), .A2 (finalResult[27]));
INV_X1 i_363 (.ZN (n_299), .A (n_300));
NOR2_X1 i_362 (.ZN (n_298), .A1 (p_0[25]), .A2 (finalResult[25]));
INV_X1 i_361 (.ZN (n_297), .A (n_298));
NOR2_X1 i_360 (.ZN (n_296), .A1 (p_0[26]), .A2 (finalResult[26]));
INV_X1 i_359 (.ZN (n_295), .A (n_296));
NAND3_X1 i_358 (.ZN (n_294), .A1 (n_299), .A2 (n_295), .A3 (n_297));
NOR2_X1 i_357 (.ZN (n_293), .A1 (p_0[24]), .A2 (finalResult[24]));
NOR2_X1 i_353 (.ZN (n_289), .A1 (p_0[19]), .A2 (finalResult[19]));
INV_X1 i_352 (.ZN (n_288), .A (n_289));
NOR2_X1 i_351 (.ZN (n_287), .A1 (p_0[17]), .A2 (finalResult[17]));
INV_X1 i_350 (.ZN (n_286), .A (n_287));
NOR2_X1 i_349 (.ZN (n_285), .A1 (p_0[18]), .A2 (finalResult[18]));
INV_X1 i_348 (.ZN (n_284), .A (n_285));
NAND3_X1 i_347 (.ZN (n_283), .A1 (n_288), .A2 (n_284), .A3 (n_286));
NOR2_X1 i_346 (.ZN (n_282), .A1 (p_0[16]), .A2 (finalResult[16]));
NAND2_X1 i_343 (.ZN (n_279), .A1 (p_0[16]), .A2 (finalResult[16]));
NAND2_X1 i_342 (.ZN (n_278), .A1 (p_0[17]), .A2 (finalResult[17]));
INV_X1 i_341 (.ZN (n_277), .A (n_278));
AOI21_X1 i_340 (.ZN (n_276), .A (n_283), .B1 (n_279), .B2 (n_278));
AND2_X1 i_339 (.ZN (n_275), .A1 (p_0[18]), .A2 (finalResult[18]));
NAND2_X1 i_337 (.ZN (n_273), .A1 (p_0[24]), .A2 (finalResult[24]));
NAND2_X1 i_336 (.ZN (n_272), .A1 (p_0[25]), .A2 (finalResult[25]));
INV_X1 i_335 (.ZN (n_271), .A (n_272));
AOI21_X1 i_334 (.ZN (n_270), .A (n_294), .B1 (n_273), .B2 (n_272));
AND2_X1 i_333 (.ZN (n_269), .A1 (p_0[26]), .A2 (finalResult[26]));
NAND2_X1 i_331 (.ZN (n_267), .A1 (p_0[28]), .A2 (finalResult[28]));
AND2_X1 i_330 (.ZN (n_266), .A1 (p_0[29]), .A2 (finalResult[29]));
AOI21_X1 i_329 (.ZN (n_265), .A (n_266), .B1 (p_0[28]), .B2 (finalResult[28]));
NAND2_X1 i_328 (.ZN (n_264), .A1 (p_0[30]), .A2 (finalResult[30]));
INV_X1 i_327 (.ZN (n_263), .A (n_264));
NAND2_X1 i_325 (.ZN (n_261), .A1 (p_0[20]), .A2 (finalResult[20]));
NAND2_X1 i_324 (.ZN (n_260), .A1 (p_0[21]), .A2 (finalResult[21]));
INV_X1 i_323 (.ZN (n_259), .A (n_260));
AOI21_X1 i_322 (.ZN (n_258), .A (n_311), .B1 (n_261), .B2 (n_260));
AND2_X1 i_321 (.ZN (n_257), .A1 (p_0[22]), .A2 (finalResult[22]));
NOR2_X1 i_317 (.ZN (n_253), .A1 (p_0[36]), .A2 (finalResult[36]));
OR2_X1 i_309 (.ZN (n_245), .A1 (n_253), .A2 (n_246));
NOR2_X1 i_305 (.ZN (n_241), .A1 (n_243), .A2 (n_242));
NOR2_X1 i_295 (.ZN (n_231), .A1 (p_0[40]), .A2 (finalResult[40]));
OR2_X1 i_294 (.ZN (n_230), .A1 (n_232), .A2 (n_231));
NOR2_X1 i_284 (.ZN (n_220), .A1 (p_0[32]), .A2 (finalResult[32]));
INV_X1 i_279 (.ZN (n_215), .A (n_216));
INV_X1 i_272 (.ZN (n_208), .A (n_209));
NAND2_X1 i_268 (.ZN (n_204), .A1 (p_0[44]), .A2 (finalResult[44]));
INV_X1 i_263 (.ZN (n_199), .A (n_200));
INV_X1 i_258 (.ZN (n_194), .A (n_195));
NOR2_X1 i_252 (.ZN (n_188), .A1 (p_0[51]), .A2 (finalResult[51]));
NOR2_X1 i_251 (.ZN (n_187), .A1 (p_0[49]), .A2 (finalResult[49]));
NOR2_X1 i_250 (.ZN (n_186), .A1 (p_0[50]), .A2 (finalResult[50]));
NAND2_X1 i_246 (.ZN (n_182), .A1 (p_0[48]), .A2 (finalResult[48]));
NAND2_X1 i_245 (.ZN (n_181), .A1 (p_0[49]), .A2 (finalResult[49]));
NAND2_X1 i_242 (.ZN (n_178), .A1 (p_0[50]), .A2 (finalResult[50]));
INV_X1 i_241 (.ZN (n_177), .A (n_178));
NOR2_X1 i_238 (.ZN (n_174), .A1 (p_0[59]), .A2 (finalResult[59]));
NOR2_X1 i_237 (.ZN (n_173), .A1 (p_0[57]), .A2 (finalResult[57]));
NOR2_X1 i_236 (.ZN (n_172), .A1 (p_0[58]), .A2 (finalResult[58]));
NOR2_X1 i_235 (.ZN (n_171), .A1 (n_173), .A2 (n_172));
NOR3_X1 i_234 (.ZN (n_170), .A1 (n_174), .A2 (n_172), .A3 (n_173));
NOR2_X1 i_232 (.ZN (n_168), .A1 (p_0[55]), .A2 (finalResult[55]));
INV_X1 i_231 (.ZN (n_167), .A (n_168));
NOR2_X1 i_230 (.ZN (n_166), .A1 (p_0[53]), .A2 (finalResult[53]));
INV_X1 i_229 (.ZN (n_165), .A (n_166));
NOR2_X1 i_228 (.ZN (n_164), .A1 (p_0[54]), .A2 (finalResult[54]));
INV_X1 i_227 (.ZN (n_163), .A (n_164));
NAND3_X1 i_226 (.ZN (n_162), .A1 (n_167), .A2 (n_163), .A3 (n_165));
NOR2_X1 i_225 (.ZN (n_161), .A1 (p_0[52]), .A2 (finalResult[52]));
NAND2_X1 i_222 (.ZN (n_158), .A1 (p_0[52]), .A2 (finalResult[52]));
NAND2_X1 i_221 (.ZN (n_157), .A1 (p_0[53]), .A2 (finalResult[53]));
INV_X1 i_220 (.ZN (n_156), .A (n_157));
AOI21_X1 i_219 (.ZN (n_155), .A (n_162), .B1 (n_158), .B2 (n_157));
AND2_X1 i_218 (.ZN (n_154), .A1 (p_0[54]), .A2 (finalResult[54]));
AOI221_X1 i_217 (.ZN (n_153), .A (n_155), .B1 (p_0[55]), .B2 (finalResult[55]), .C1 (n_167), .C2 (n_154));
NAND2_X1 i_215 (.ZN (n_151), .A1 (p_0[56]), .A2 (finalResult[56]));
INV_X1 i_214 (.ZN (n_150), .A (n_151));
AND2_X1 i_213 (.ZN (n_149), .A1 (p_0[57]), .A2 (finalResult[57]));
OAI21_X1 i_212 (.ZN (n_148), .A (n_170), .B1 (n_150), .B2 (n_149));
NAND2_X1 i_210 (.ZN (n_146), .A1 (p_0[58]), .A2 (finalResult[58]));
INV_X1 i_209 (.ZN (n_145), .A (n_146));
OAI21_X1 i_200 (.ZN (n_136), .A (n_137), .B1 (n_379), .B2 (n_375));
AOI22_X1 i_191 (.ZN (p_1[61]), .A1 (n_140), .A2 (n_136), .B1 (n_141), .B2 (n_135));
XNOR2_X1 i_190 (.ZN (p_1[60]), .A (n_143), .B (n_142));
AOI21_X1 i_189 (.ZN (n_129), .A (n_174), .B1 (p_0[59]), .B2 (finalResult[59]));
OAI21_X1 i_188 (.ZN (n_128), .A (n_153), .B1 (n_175), .B2 (n_160));
OAI21_X1 i_187 (.ZN (n_127), .A (n_151), .B1 (p_0[56]), .B2 (finalResult[56]));
OAI22_X1 i_186 (.ZN (n_126), .A1 (p_0[56]), .A2 (finalResult[56]), .B1 (n_150), .B2 (n_128));
INV_X1 i_185 (.ZN (n_125), .A (n_126));
NOR2_X1 i_184 (.ZN (n_124), .A1 (n_173), .A2 (n_149));
NAND3_X1 i_183 (.ZN (n_123), .A1 (n_146), .A2 (n_124), .A3 (n_126));
OAI21_X1 i_182 (.ZN (n_122), .A (n_123), .B1 (n_171), .B2 (n_145));
XNOR2_X1 i_181 (.ZN (p_1[59]), .A (n_129), .B (n_122));
NOR2_X1 i_180 (.ZN (n_121), .A1 (n_172), .A2 (n_145));
OAI22_X1 i_179 (.ZN (n_120), .A1 (p_0[57]), .A2 (finalResult[57]), .B1 (n_149), .B2 (n_125));
XNOR2_X1 i_178 (.ZN (p_1[58]), .A (n_121), .B (n_120));
XOR2_X1 i_177 (.Z (p_1[57]), .A (n_125), .B (n_124));
XNOR2_X1 i_176 (.ZN (p_1[56]), .A (n_128), .B (n_127));
AOI21_X1 i_175 (.ZN (n_119), .A (n_168), .B1 (p_0[55]), .B2 (finalResult[55]));
OAI21_X1 i_174 (.ZN (n_118), .A (n_158), .B1 (p_0[52]), .B2 (finalResult[52]));
AOI21_X1 i_173 (.ZN (n_117), .A (n_161), .B1 (n_175), .B2 (n_158));
OAI21_X1 i_172 (.ZN (n_116), .A (n_165), .B1 (n_156), .B2 (n_117));
INV_X1 i_171 (.ZN (n_115), .A (n_116));
NOR2_X1 i_170 (.ZN (n_114), .A1 (n_166), .A2 (n_156));
OAI21_X1 i_169 (.ZN (n_113), .A (n_163), .B1 (n_154), .B2 (n_115));
XNOR2_X1 i_168 (.ZN (p_1[55]), .A (n_119), .B (n_113));
NOR2_X1 i_167 (.ZN (n_112), .A1 (n_164), .A2 (n_154));
XOR2_X1 i_166 (.Z (p_1[54]), .A (n_115), .B (n_112));
XOR2_X1 i_165 (.Z (p_1[53]), .A (n_117), .B (n_114));
XOR2_X1 i_164 (.Z (p_1[52]), .A (n_175), .B (n_118));
NOR2_X1 i_163 (.ZN (n_111), .A1 (n_188), .A2 (n_179));
OAI21_X1 i_162 (.ZN (n_110), .A (n_182), .B1 (p_0[48]), .B2 (finalResult[48]));
AOI21_X1 i_161 (.ZN (n_109), .A (n_184), .B1 (n_189), .B2 (n_182));
INV_X1 i_160 (.ZN (n_108), .A (n_109));
AOI21_X1 i_159 (.ZN (n_107), .A (n_187), .B1 (n_181), .B2 (n_108));
AOI21_X1 i_158 (.ZN (n_106), .A (n_187), .B1 (p_0[49]), .B2 (finalResult[49]));
OAI22_X1 i_157 (.ZN (n_105), .A1 (p_0[50]), .A2 (finalResult[50]), .B1 (n_177), .B2 (n_107));
XNOR2_X1 i_156 (.ZN (p_1[51]), .A (n_111), .B (n_105));
NOR2_X1 i_155 (.ZN (n_104), .A1 (n_186), .A2 (n_177));
XOR2_X1 i_154 (.Z (p_1[50]), .A (n_107), .B (n_104));
XOR2_X1 i_153 (.Z (p_1[49]), .A (n_109), .B (n_106));
XOR2_X1 i_152 (.Z (p_1[48]), .A (n_189), .B (n_110));
AOI21_X1 i_151 (.ZN (n_103), .A (n_244), .B1 (p_0[47]), .B2 (finalResult[47]));
OAI21_X1 i_150 (.ZN (n_102), .A (n_212), .B1 (n_254), .B2 (n_219));
INV_X1 i_149 (.ZN (n_101), .A (n_102));
OAI21_X1 i_148 (.ZN (n_100), .A (n_205), .B1 (n_245), .B2 (n_101));
INV_X1 i_147 (.ZN (n_99), .A (n_100));
OAI21_X1 i_146 (.ZN (n_98), .A (n_191), .B1 (n_230), .B2 (n_99));
OAI21_X1 i_145 (.ZN (n_97), .A (n_204), .B1 (p_0[44]), .B2 (finalResult[44]));
OAI22_X1 i_144 (.ZN (n_96), .A1 (p_0[44]), .A2 (finalResult[44]), .B1 (n_203), .B2 (n_98));
INV_X1 i_143 (.ZN (n_95), .A (n_96));
NOR2_X1 i_142 (.ZN (n_94), .A1 (n_243), .A2 (n_202));
NAND3_X1 i_141 (.ZN (n_93), .A1 (n_200), .A2 (n_94), .A3 (n_96));
OAI21_X1 i_140 (.ZN (n_92), .A (n_93), .B1 (n_241), .B2 (n_199));
XNOR2_X1 i_139 (.ZN (p_1[47]), .A (n_103), .B (n_92));
NOR2_X1 i_138 (.ZN (n_91), .A1 (n_242), .A2 (n_199));
OAI22_X1 i_137 (.ZN (n_90), .A1 (p_0[45]), .A2 (finalResult[45]), .B1 (n_202), .B2 (n_95));
XNOR2_X1 i_136 (.ZN (p_1[46]), .A (n_91), .B (n_90));
XOR2_X1 i_135 (.Z (p_1[45]), .A (n_95), .B (n_94));
XNOR2_X1 i_134 (.ZN (p_1[44]), .A (n_98), .B (n_97));
AOI21_X1 i_133 (.ZN (n_89), .A (n_238), .B1 (p_0[43]), .B2 (finalResult[43]));
OAI21_X1 i_132 (.ZN (n_88), .A (n_196), .B1 (p_0[40]), .B2 (finalResult[40]));
AOI21_X1 i_131 (.ZN (n_87), .A (n_231), .B1 (n_196), .B2 (n_99));
OAI21_X1 i_130 (.ZN (n_86), .A (n_235), .B1 (n_194), .B2 (n_87));
INV_X1 i_129 (.ZN (n_85), .A (n_86));
NOR2_X1 i_128 (.ZN (n_84), .A1 (n_236), .A2 (n_194));
OAI21_X1 i_127 (.ZN (n_83), .A (n_233), .B1 (n_192), .B2 (n_85));
XNOR2_X1 i_126 (.ZN (p_1[43]), .A (n_89), .B (n_83));
NOR2_X1 i_125 (.ZN (n_82), .A1 (n_234), .A2 (n_192));
XOR2_X1 i_124 (.Z (p_1[42]), .A (n_85), .B (n_82));
XOR2_X1 i_123 (.Z (p_1[41]), .A (n_87), .B (n_84));
XOR2_X1 i_122 (.Z (p_1[40]), .A (n_99), .B (n_88));
AOI21_X1 i_121 (.ZN (n_81), .A (n_252), .B1 (p_0[39]), .B2 (finalResult[39]));
OAI21_X1 i_120 (.ZN (n_80), .A (n_210), .B1 (p_0[36]), .B2 (finalResult[36]));
AOI21_X1 i_119 (.ZN (n_79), .A (n_253), .B1 (n_210), .B2 (n_101));
OAI21_X1 i_118 (.ZN (n_78), .A (n_249), .B1 (n_208), .B2 (n_79));
INV_X1 i_117 (.ZN (n_77), .A (n_78));
NOR2_X1 i_116 (.ZN (n_76), .A1 (n_250), .A2 (n_208));
OAI21_X1 i_115 (.ZN (n_75), .A (n_247), .B1 (n_206), .B2 (n_77));
XNOR2_X1 i_114 (.ZN (p_1[39]), .A (n_81), .B (n_75));
NOR2_X1 i_113 (.ZN (n_74), .A1 (n_248), .A2 (n_206));
XOR2_X1 i_112 (.Z (p_1[38]), .A (n_77), .B (n_74));
XOR2_X1 i_111 (.Z (p_1[37]), .A (n_79), .B (n_76));
XOR2_X1 i_110 (.Z (p_1[36]), .A (n_101), .B (n_80));
AOI21_X1 i_109 (.ZN (n_73), .A (n_227), .B1 (p_0[35]), .B2 (finalResult[35]));
OAI21_X1 i_108 (.ZN (n_72), .A (n_217), .B1 (p_0[32]), .B2 (finalResult[32]));
AOI21_X1 i_107 (.ZN (n_71), .A (n_220), .B1 (n_254), .B2 (n_217));
OAI21_X1 i_106 (.ZN (n_70), .A (n_224), .B1 (n_215), .B2 (n_71));
INV_X1 i_105 (.ZN (n_69), .A (n_70));
NOR2_X1 i_104 (.ZN (n_68), .A1 (n_225), .A2 (n_215));
OAI21_X1 i_103 (.ZN (n_67), .A (n_222), .B1 (n_213), .B2 (n_69));
XNOR2_X1 i_102 (.ZN (p_1[35]), .A (n_73), .B (n_67));
NOR2_X1 i_101 (.ZN (n_66), .A1 (n_223), .A2 (n_213));
XOR2_X1 i_100 (.Z (p_1[34]), .A (n_69), .B (n_66));
XOR2_X1 i_99 (.Z (p_1[33]), .A (n_71), .B (n_68));
XOR2_X1 i_98 (.Z (p_1[32]), .A (n_254), .B (n_72));
OAI21_X1 i_97 (.ZN (n_65), .A (n_308), .B1 (n_377), .B2 (n_373));
OAI21_X1 i_96 (.ZN (n_64), .A (n_274), .B1 (n_319), .B2 (n_281));
INV_X1 i_95 (.ZN (n_63), .A (n_64));
OAI21_X1 i_94 (.ZN (n_62), .A (n_256), .B1 (n_310), .B2 (n_63));
INV_X1 i_93 (.ZN (n_61), .A (n_62));
OAI21_X1 i_92 (.ZN (n_60), .A (n_268), .B1 (n_292), .B2 (n_61));
INV_X1 i_91 (.ZN (n_59), .A (n_60));
OAI21_X1 i_90 (.ZN (n_58), .A (n_267), .B1 (p_0[28]), .B2 (finalResult[28]));
AOI21_X1 i_89 (.ZN (n_57), .A (n_302), .B1 (n_267), .B2 (n_59));
OAI21_X1 i_88 (.ZN (n_56), .A (n_306), .B1 (n_266), .B2 (n_57));
INV_X1 i_87 (.ZN (n_55), .A (n_56));
NOR2_X1 i_86 (.ZN (n_54), .A1 (n_307), .A2 (n_266));
OAI21_X1 i_85 (.ZN (n_53), .A (n_304), .B1 (n_263), .B2 (n_55));
XOR2_X1 i_84 (.Z (p_1[31]), .A (n_65), .B (n_53));
NOR2_X1 i_83 (.ZN (n_52), .A1 (n_305), .A2 (n_263));
XOR2_X1 i_82 (.Z (p_1[30]), .A (n_55), .B (n_52));
XOR2_X1 i_81 (.Z (p_1[29]), .A (n_57), .B (n_54));
XOR2_X1 i_80 (.Z (p_1[28]), .A (n_59), .B (n_58));
AOI21_X1 i_79 (.ZN (n_51), .A (n_300), .B1 (p_0[27]), .B2 (finalResult[27]));
OAI21_X1 i_78 (.ZN (n_50), .A (n_273), .B1 (p_0[24]), .B2 (finalResult[24]));
AOI21_X1 i_77 (.ZN (n_49), .A (n_293), .B1 (n_273), .B2 (n_61));
OAI21_X1 i_76 (.ZN (n_48), .A (n_297), .B1 (n_271), .B2 (n_49));
INV_X1 i_75 (.ZN (n_47), .A (n_48));
NOR2_X1 i_74 (.ZN (n_46), .A1 (n_298), .A2 (n_271));
OAI21_X1 i_73 (.ZN (n_45), .A (n_295), .B1 (n_269), .B2 (n_47));
XNOR2_X1 i_72 (.ZN (p_1[27]), .A (n_51), .B (n_45));
NOR2_X1 i_71 (.ZN (n_44), .A1 (n_296), .A2 (n_269));
XOR2_X1 i_70 (.Z (p_1[26]), .A (n_47), .B (n_44));
XOR2_X1 i_69 (.Z (p_1[25]), .A (n_49), .B (n_46));
XOR2_X1 i_68 (.Z (p_1[24]), .A (n_61), .B (n_50));
AOI21_X1 i_67 (.ZN (n_43), .A (n_317), .B1 (p_0[23]), .B2 (finalResult[23]));
OAI21_X1 i_66 (.ZN (n_42), .A (n_261), .B1 (p_0[20]), .B2 (finalResult[20]));
AOI21_X1 i_65 (.ZN (n_41), .A (n_318), .B1 (n_261), .B2 (n_63));
OAI21_X1 i_64 (.ZN (n_40), .A (n_314), .B1 (n_259), .B2 (n_41));
INV_X1 i_63 (.ZN (n_39), .A (n_40));
NOR2_X1 i_62 (.ZN (n_38), .A1 (n_315), .A2 (n_259));
OAI21_X1 i_61 (.ZN (n_37), .A (n_312), .B1 (n_257), .B2 (n_39));
XNOR2_X1 i_60 (.ZN (p_1[23]), .A (n_43), .B (n_37));
NOR2_X1 i_59 (.ZN (n_36), .A1 (n_313), .A2 (n_257));
XOR2_X1 i_58 (.Z (p_1[22]), .A (n_39), .B (n_36));
XOR2_X1 i_57 (.Z (p_1[21]), .A (n_41), .B (n_38));
XOR2_X1 i_56 (.Z (p_1[20]), .A (n_63), .B (n_42));
AOI21_X1 i_55 (.ZN (n_35), .A (n_289), .B1 (p_0[19]), .B2 (finalResult[19]));
OAI21_X1 i_54 (.ZN (n_34), .A (n_279), .B1 (p_0[16]), .B2 (finalResult[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_282), .B1 (n_319), .B2 (n_279));
OAI21_X1 i_52 (.ZN (n_32), .A (n_286), .B1 (n_277), .B2 (n_33));
INV_X1 i_51 (.ZN (n_31), .A (n_32));
NOR2_X1 i_50 (.ZN (n_30), .A1 (n_287), .A2 (n_277));
OAI21_X1 i_49 (.ZN (n_29), .A (n_284), .B1 (n_275), .B2 (n_31));
XNOR2_X1 i_48 (.ZN (p_1[19]), .A (n_35), .B (n_29));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_285), .A2 (n_275));
XOR2_X1 i_46 (.Z (p_1[18]), .A (n_31), .B (n_28));
XOR2_X1 i_45 (.Z (p_1[17]), .A (n_33), .B (n_30));
XOR2_X1 i_44 (.Z (p_1[16]), .A (n_319), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_332), .A2 (n_323));
OAI21_X1 i_42 (.ZN (n_26), .A (n_326), .B1 (p_0[12]), .B2 (finalResult[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_328), .B1 (n_333), .B2 (n_326));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_331), .B1 (n_325), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_331), .B1 (p_0[13]), .B2 (finalResult[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (p_0[14]), .A2 (finalResult[14]), .B1 (n_321), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (p_1[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_330), .A2 (n_321));
XOR2_X1 i_34 (.Z (p_1[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (p_1[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (p_1[12]), .A (n_333), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_346), .A2 (n_337));
AOI21_X1 i_30 (.ZN (n_18), .A (n_342), .B1 (p_0[8]), .B2 (finalResult[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_342), .B1 (n_347), .B2 (n_340));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_345), .B1 (n_339), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_345), .B1 (p_0[9]), .B2 (finalResult[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (p_0[10]), .A2 (finalResult[10]), .B1 (n_335), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (p_1[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_344), .A2 (n_335));
XOR2_X1 i_22 (.Z (p_1[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (p_1[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (p_1[8]), .A (n_347), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_360), .A2 (n_351));
OAI21_X1 i_18 (.ZN (n_10), .A (n_354), .B1 (p_0[4]), .B2 (finalResult[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_356), .B1 (n_361), .B2 (n_354));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_359), .B1 (n_353), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_359), .B1 (p_0[5]), .B2 (finalResult[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (p_0[6]), .A2 (finalResult[6]), .B1 (n_349), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (p_1[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_358), .A2 (n_349));
XOR2_X1 i_10 (.Z (p_1[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (p_1[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (p_1[4]), .A (n_361), .B (n_10));
OAI21_X1 i_7 (.ZN (n_3), .A (n_370), .B1 (n_376), .B2 (n_372));
XOR2_X1 i_6 (.Z (p_1[3]), .A (n_363), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_369), .B1 (p_0[2]), .B2 (finalResult[2]));
XNOR2_X1 i_4 (.ZN (p_1[2]), .A (n_364), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_365), .B1 (p_0[1]), .B2 (finalResult[1]));
XOR2_X1 i_2 (.Z (p_1[1]), .A (n_366), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_366), .B1 (p_0[0]), .B2 (finalResult[0]));
INV_X1 i_0 (.ZN (p_1[0]), .A (n_0));

endmodule //datapath__0_10

module datapath (firstInputComplement, inputOne);

output [31:0] firstInputComplement;
input [31:0] inputOne;
wire n_3;
wire n_12;
wire n_5;
wire n_10;
wire n_11;
wire n_22;
wire n_0;
wire n_8;
wire n_20;
wire n_21;
wire n_18;
wire n_19;
wire n_38;
wire n_30;
wire n_36;
wire n_37;
wire n_51;
wire n_44;
wire n_49;
wire n_50;
wire n_61;
wire n_56;
wire n_77;
wire n_63;
wire n_68;
wire n_69;
wire n_80;
wire n_74;
wire n_83;
wire n_1;
wire n_2;
wire n_4;
wire n_6;
wire n_9;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_32;
wire n_29;
wire n_33;
wire n_31;
wire n_34;
wire n_35;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_46;
wire n_43;
wire n_45;
wire n_47;
wire n_48;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_58;
wire n_57;
wire n_59;
wire n_60;
wire n_62;
wire n_65;
wire n_64;
wire n_66;
wire n_67;
wire n_71;
wire n_70;
wire n_72;
wire n_73;
wire n_76;
wire n_75;
wire n_78;
wire n_79;
wire n_82;
wire n_81;
wire n_84;
wire n_85;
wire n_86;


INV_X1 i_117 (.ZN (n_86), .A (inputOne[31]));
NAND4_X1 i_116 (.ZN (n_85), .A1 (n_62), .A2 (n_70), .A3 (n_75), .A4 (n_82));
AND4_X1 i_115 (.ZN (n_84), .A1 (n_86), .A2 (n_77), .A3 (n_75), .A4 (n_82));
AOI21_X1 i_114 (.ZN (firstInputComplement[31]), .A (n_84), .B1 (inputOne[31]), .B2 (n_85));
NOR2_X1 i_113 (.ZN (n_83), .A1 (inputOne[29]), .A2 (inputOne[28]));
NOR3_X1 i_112 (.ZN (n_82), .A1 (inputOne[29]), .A2 (inputOne[28]), .A3 (inputOne[30]));
NAND3_X1 i_111 (.ZN (n_81), .A1 (n_77), .A2 (n_75), .A3 (n_83));
AOI22_X1 i_110 (.ZN (firstInputComplement[30]), .A1 (n_74), .A2 (n_82), .B1 (inputOne[30]), .B2 (n_81));
INV_X1 i_109 (.ZN (n_80), .A (n_79));
AOI21_X1 i_108 (.ZN (firstInputComplement[28]), .A (n_79), .B1 (inputOne[28]), .B2 (n_78));
NOR2_X1 i_107 (.ZN (n_79), .A1 (n_78), .A2 (inputOne[28]));
NAND2_X1 i_106 (.ZN (n_78), .A1 (n_77), .A2 (n_75));
INV_X1 i_105 (.ZN (n_77), .A (n_69));
INV_X1 i_104 (.ZN (n_76), .A (n_72));
NOR2_X1 i_103 (.ZN (n_75), .A1 (n_73), .A2 (inputOne[27]));
NOR3_X1 i_102 (.ZN (n_74), .A1 (n_73), .A2 (inputOne[27]), .A3 (n_69));
AOI21_X1 i_101 (.ZN (firstInputComplement[27]), .A (n_74), .B1 (inputOne[27]), .B2 (n_76));
OR3_X1 i_100 (.ZN (n_73), .A1 (inputOne[26]), .A2 (inputOne[24]), .A3 (inputOne[25]));
NOR2_X1 i_99 (.ZN (n_72), .A1 (n_69), .A2 (n_73));
AOI21_X1 i_98 (.ZN (firstInputComplement[26]), .A (n_72), .B1 (inputOne[26]), .B2 (n_67));
INV_X1 i_97 (.ZN (n_71), .A (inputOne[25]));
INV_X1 i_96 (.ZN (n_70), .A (inputOne[23]));
NAND4_X1 i_95 (.ZN (n_69), .A1 (n_70), .A2 (n_43), .A3 (n_57), .A4 (n_64));
NOR2_X1 i_94 (.ZN (n_68), .A1 (inputOne[24]), .A2 (n_69));
NAND2_X1 i_93 (.ZN (n_67), .A1 (n_71), .A2 (n_68));
OAI21_X1 i_92 (.ZN (n_66), .A (n_67), .B1 (n_71), .B2 (n_68));
INV_X1 i_91 (.ZN (firstInputComplement[25]), .A (n_66));
INV_X1 i_90 (.ZN (n_65), .A (n_59));
NOR3_X1 i_89 (.ZN (n_64), .A1 (inputOne[22]), .A2 (inputOne[20]), .A3 (inputOne[21]));
NAND4_X1 i_88 (.ZN (n_63), .A1 (n_29), .A2 (n_45), .A3 (n_57), .A4 (n_64));
INV_X1 i_87 (.ZN (n_62), .A (n_63));
AOI21_X1 i_86 (.ZN (firstInputComplement[22]), .A (n_62), .B1 (inputOne[22]), .B2 (n_65));
NOR2_X1 i_85 (.ZN (n_61), .A1 (inputOne[20]), .A2 (n_56));
INV_X1 i_84 (.ZN (n_60), .A (n_61));
NOR2_X1 i_83 (.ZN (n_59), .A1 (inputOne[21]), .A2 (n_60));
AOI21_X1 i_82 (.ZN (firstInputComplement[21]), .A (n_59), .B1 (inputOne[21]), .B2 (n_60));
INV_X1 i_81 (.ZN (n_58), .A (inputOne[19]));
AND4_X1 i_80 (.ZN (n_57), .A1 (n_53), .A2 (n_52), .A3 (n_58), .A4 (n_54));
NAND2_X1 i_79 (.ZN (n_56), .A1 (n_43), .A2 (n_57));
OAI21_X1 i_78 (.ZN (n_55), .A (n_56), .B1 (n_58), .B2 (n_47));
INV_X1 i_77 (.ZN (firstInputComplement[19]), .A (n_55));
INV_X1 i_76 (.ZN (n_54), .A (inputOne[18]));
INV_X1 i_75 (.ZN (n_53), .A (inputOne[17]));
INV_X1 i_74 (.ZN (n_52), .A (inputOne[16]));
NOR2_X1 i_73 (.ZN (n_51), .A1 (inputOne[16]), .A2 (n_44));
INV_X1 i_72 (.ZN (n_50), .A (n_51));
NOR2_X1 i_71 (.ZN (n_49), .A1 (inputOne[17]), .A2 (n_50));
INV_X1 i_70 (.ZN (n_48), .A (n_49));
NOR2_X1 i_69 (.ZN (n_47), .A1 (inputOne[18]), .A2 (n_48));
AOI21_X1 i_68 (.ZN (firstInputComplement[18]), .A (n_47), .B1 (inputOne[18]), .B2 (n_48));
INV_X1 i_67 (.ZN (n_46), .A (inputOne[15]));
AND4_X1 i_66 (.ZN (n_45), .A1 (n_40), .A2 (n_39), .A3 (n_46), .A4 (n_41));
NAND4_X1 i_65 (.ZN (n_44), .A1 (n_6), .A2 (n_31), .A3 (n_45), .A4 (n_33));
INV_X1 i_64 (.ZN (n_43), .A (n_44));
OAI21_X1 i_63 (.ZN (n_42), .A (n_44), .B1 (n_46), .B2 (n_34));
INV_X1 i_62 (.ZN (firstInputComplement[15]), .A (n_42));
INV_X1 i_61 (.ZN (n_41), .A (inputOne[14]));
INV_X1 i_60 (.ZN (n_40), .A (inputOne[13]));
INV_X1 i_59 (.ZN (n_39), .A (inputOne[12]));
NOR2_X1 i_58 (.ZN (n_38), .A1 (inputOne[12]), .A2 (n_30));
INV_X1 i_57 (.ZN (n_37), .A (n_38));
NOR2_X1 i_56 (.ZN (n_36), .A1 (inputOne[13]), .A2 (n_37));
INV_X1 i_55 (.ZN (n_35), .A (n_36));
NOR2_X1 i_54 (.ZN (n_34), .A1 (inputOne[14]), .A2 (n_35));
AOI21_X1 i_53 (.ZN (firstInputComplement[14]), .A (n_34), .B1 (inputOne[14]), .B2 (n_35));
INV_X1 i_52 (.ZN (n_33), .A (n_23));
INV_X1 i_51 (.ZN (n_32), .A (inputOne[11]));
AND4_X1 i_50 (.ZN (n_31), .A1 (n_26), .A2 (n_25), .A3 (n_32), .A4 (n_27));
NAND3_X1 i_49 (.ZN (n_30), .A1 (n_33), .A2 (n_6), .A3 (n_31));
INV_X1 i_48 (.ZN (n_29), .A (n_30));
OAI21_X1 i_47 (.ZN (n_28), .A (n_30), .B1 (n_32), .B2 (n_16));
INV_X1 i_46 (.ZN (firstInputComplement[11]), .A (n_28));
INV_X1 i_45 (.ZN (n_27), .A (inputOne[10]));
INV_X1 i_44 (.ZN (n_26), .A (inputOne[9]));
INV_X1 i_42 (.ZN (n_25), .A (inputOne[8]));
INV_X1 i_41 (.ZN (n_24), .A (inputOne[7]));
NAND4_X1 i_40 (.ZN (n_23), .A1 (n_14), .A2 (n_13), .A3 (n_24), .A4 (n_15));
NOR2_X1 i_39 (.ZN (n_22), .A1 (n_5), .A2 (n_23));
INV_X1 i_38 (.ZN (n_21), .A (n_22));
NOR2_X1 i_37 (.ZN (n_20), .A1 (inputOne[8]), .A2 (n_21));
INV_X1 i_36 (.ZN (n_19), .A (n_20));
NOR2_X1 i_35 (.ZN (n_18), .A1 (inputOne[9]), .A2 (n_19));
INV_X1 i_32 (.ZN (n_17), .A (n_18));
NOR2_X1 i_31 (.ZN (n_16), .A1 (inputOne[10]), .A2 (n_17));
AOI21_X1 i_30 (.ZN (firstInputComplement[10]), .A (n_16), .B1 (inputOne[10]), .B2 (n_17));
INV_X1 i_29 (.ZN (n_15), .A (inputOne[6]));
INV_X1 i_28 (.ZN (n_14), .A (inputOne[5]));
INV_X1 i_27 (.ZN (n_13), .A (inputOne[4]));
NOR2_X1 i_26 (.ZN (n_12), .A1 (inputOne[4]), .A2 (n_5));
INV_X1 i_25 (.ZN (n_11), .A (n_12));
NOR2_X1 i_22 (.ZN (n_10), .A1 (inputOne[5]), .A2 (n_11));
INV_X1 i_21 (.ZN (n_9), .A (n_10));
NOR2_X1 i_20 (.ZN (n_8), .A1 (inputOne[6]), .A2 (n_9));
AOI21_X1 i_19 (.ZN (firstInputComplement[6]), .A (n_8), .B1 (inputOne[6]), .B2 (n_9));
NOR4_X1 i_17 (.ZN (n_6), .A1 (inputOne[3]), .A2 (inputOne[0]), .A3 (inputOne[2]), .A4 (inputOne[1]));
INV_X1 i_16 (.ZN (n_5), .A (n_6));
AOI21_X1 i_15 (.ZN (firstInputComplement[3]), .A (n_6), .B1 (inputOne[3]), .B2 (n_2));
INV_X1 i_14 (.ZN (n_4), .A (inputOne[2]));
NOR2_X1 i_13 (.ZN (n_3), .A1 (inputOne[1]), .A2 (inputOne[0]));
NAND2_X1 i_12 (.ZN (n_2), .A1 (n_4), .A2 (n_3));
OAI21_X1 i_11 (.ZN (n_1), .A (n_2), .B1 (n_4), .B2 (n_3));
INV_X1 i_10 (.ZN (firstInputComplement[2]), .A (n_1));
AOI22_X1 i_9 (.ZN (firstInputComplement[29]), .A1 (n_80), .A2 (inputOne[29]), .B1 (n_74), .B2 (n_83));
AOI21_X1 i_8 (.ZN (firstInputComplement[24]), .A (n_68), .B1 (inputOne[24]), .B2 (n_69));
AOI21_X1 i_7 (.ZN (firstInputComplement[23]), .A (n_77), .B1 (inputOne[23]), .B2 (n_63));
AOI21_X1 i_43 (.ZN (firstInputComplement[20]), .A (n_61), .B1 (inputOne[20]), .B2 (n_56));
AOI21_X1 i_34 (.ZN (firstInputComplement[17]), .A (n_49), .B1 (inputOne[17]), .B2 (n_50));
AOI21_X1 i_33 (.ZN (firstInputComplement[16]), .A (n_51), .B1 (inputOne[16]), .B2 (n_44));
AOI21_X1 i_24 (.ZN (firstInputComplement[13]), .A (n_36), .B1 (inputOne[13]), .B2 (n_37));
AOI21_X1 i_23 (.ZN (firstInputComplement[12]), .A (n_38), .B1 (inputOne[12]), .B2 (n_30));
AOI21_X1 i_6 (.ZN (firstInputComplement[9]), .A (n_18), .B1 (inputOne[9]), .B2 (n_19));
AOI21_X1 i_5 (.ZN (firstInputComplement[8]), .A (n_20), .B1 (inputOne[8]), .B2 (n_21));
INV_X1 i_4 (.ZN (n_0), .A (n_8));
AOI21_X1 i_3 (.ZN (firstInputComplement[7]), .A (n_22), .B1 (inputOne[7]), .B2 (n_0));
AOI21_X1 i_2 (.ZN (firstInputComplement[5]), .A (n_10), .B1 (inputOne[5]), .B2 (n_11));
AOI21_X1 i_1 (.ZN (firstInputComplement[4]), .A (n_12), .B1 (inputOne[4]), .B2 (n_5));
AOI21_X1 i_0 (.ZN (firstInputComplement[1]), .A (n_3), .B1 (inputOne[1]), .B2 (inputOne[0]));

endmodule //datapath

module RadixNoaman (clk_CTS_0_PP_10, clk_CTS_0_PP_11, inputOne, inputTwo, finalResult, 
    clk, reset, enable, enableRegisterOutput);

output enableRegisterOutput;
output [63:0] finalResult;
input clk;
input enable;
input [31:0] inputOne;
input [31:0] inputTwo;
input reset;
input clk_CTS_0_PP_10;
input clk_CTS_0_PP_11;
wire CTS_n_tid0_63;
wire \firstInputComplement[31] ;
wire \firstInputComplement[30] ;
wire \firstInputComplement[29] ;
wire \firstInputComplement[28] ;
wire \firstInputComplement[27] ;
wire \firstInputComplement[26] ;
wire \firstInputComplement[25] ;
wire \firstInputComplement[24] ;
wire \firstInputComplement[23] ;
wire \firstInputComplement[22] ;
wire \firstInputComplement[21] ;
wire \firstInputComplement[20] ;
wire \firstInputComplement[19] ;
wire \firstInputComplement[18] ;
wire \firstInputComplement[17] ;
wire \firstInputComplement[16] ;
wire \firstInputComplement[15] ;
wire \firstInputComplement[14] ;
wire \firstInputComplement[13] ;
wire \firstInputComplement[12] ;
wire \firstInputComplement[11] ;
wire \firstInputComplement[10] ;
wire \firstInputComplement[9] ;
wire \firstInputComplement[8] ;
wire \firstInputComplement[7] ;
wire \firstInputComplement[6] ;
wire \firstInputComplement[5] ;
wire \firstInputComplement[4] ;
wire \firstInputComplement[3] ;
wire \firstInputComplement[2] ;
wire \firstInputComplement[1] ;
wire hfn_ipo_n35;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_1_3;
wire n_0_1_0;
wire n_0_1_4;
wire n_0_1_1;
wire n_0_1_5;
wire n_0_1_2;
wire n_0_1_6;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_185;
wire n_0_186;
wire n_0_187;
wire n_0_188;
wire n_0_189;
wire n_0_190;
wire n_0_191;
wire n_0_192;
wire n_0_193;
wire n_0_194;
wire n_0_1_7;
wire n_0_1_8;
wire n_0_1_9;
wire n_0_1_10;
wire n_0_1_11;
wire n_0_1_12;
wire n_0_1_13;
wire n_0_195;
wire n_0_196;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_201;
wire n_0_202;
wire n_0_203;
wire n_0_204;
wire n_0_205;
wire n_0_206;
wire n_0_207;
wire n_0_208;
wire n_0_209;
wire n_0_210;
wire n_0_211;
wire n_0_212;
wire n_0_213;
wire n_0_214;
wire n_0_215;
wire n_0_216;
wire n_0_217;
wire n_0_218;
wire n_0_219;
wire n_0_220;
wire n_0_221;
wire n_0_222;
wire n_0_223;
wire n_0_224;
wire n_0_225;
wire n_0_226;
wire n_0_227;
wire n_0_228;
wire n_0_229;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_233;
wire n_0_234;
wire n_0_235;
wire n_0_236;
wire n_0_237;
wire n_0_238;
wire n_0_239;
wire n_0_240;
wire n_0_241;
wire n_0_242;
wire n_0_243;
wire n_0_244;
wire n_0_245;
wire n_0_246;
wire n_0_247;
wire n_0_248;
wire n_0_249;
wire n_0_250;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_257;
wire n_0_258;
wire n_0_1_14;
wire n_0_1_15;
wire n_0_1_16;
wire n_0_1_17;
wire n_0_1_18;
wire n_0_259;
wire n_0_1_19;
wire n_0_260;
wire n_0_261;
wire n_0_262;
wire n_0_1_20;
wire n_0_263;
wire n_0_130;
wire n_0_129;
wire n_0_1_21;
wire n_0_1_22;
wire n_0_1_23;
wire n_0_1_24;
wire n_0_1_25;
wire n_0_1_26;
wire n_0_1_27;
wire n_0_1_28;
wire n_0_1_29;
wire n_0_1_30;
wire n_0_1_31;
wire n_0_1_32;
wire n_0_1_33;
wire n_0_1_34;
wire n_0_1_35;
wire n_0_1_36;
wire n_0_1_37;
wire n_0_1_38;
wire n_0_1_39;
wire n_0_1_40;
wire n_0_1_41;
wire n_0_1_42;
wire n_0_1_43;
wire n_0_1_44;
wire n_0_1_45;
wire n_0_1_46;
wire n_0_1_47;
wire n_0_1_48;
wire n_0_1_49;
wire n_0_1_50;
wire n_0_1_51;
wire n_0_1_52;
wire n_0_1_53;
wire n_0_1_54;
wire n_0_52;
wire n_0_1_55;
wire n_0_1_56;
wire n_0_1_57;
wire n_0_1_58;
wire n_0_1_59;
wire n_0_1_60;
wire n_0_1_61;
wire n_0_1_62;
wire n_0_1_63;
wire n_0_1_64;
wire n_0_1_65;
wire n_0_1_66;
wire n_0_1_67;
wire n_0_1_68;
wire n_0_1_69;
wire n_0_53;
wire n_0_1_70;
wire n_0_1_71;
wire n_0_1_72;
wire n_0_1_73;
wire n_0_1_74;
wire n_0_1_75;
wire n_0_54;
wire n_0_1_76;
wire n_0_1_77;
wire n_0_1_78;
wire n_0_1_79;
wire n_0_55;
wire n_0_1_80;
wire n_0_1_81;
wire n_0_1_82;
wire n_0_1_83;
wire n_0_1_84;
wire n_0_1_85;
wire n_0_56;
wire n_0_1_86;
wire n_0_1_87;
wire n_0_1_88;
wire n_0_1_89;
wire n_0_1_90;
wire n_0_57;
wire n_0_1_91;
wire n_0_1_92;
wire n_0_1_93;
wire n_0_1_94;
wire n_0_58;
wire n_0_1_95;
wire n_0_1_96;
wire n_0_1_97;
wire n_0_1_98;
wire n_0_59;
wire n_0_1_99;
wire n_0_1_100;
wire n_0_1_101;
wire n_0_1_102;
wire n_0_1_103;
wire n_0_1_104;
wire n_0_1_105;
wire n_0_1_106;
wire n_0_60;
wire n_0_1_107;
wire n_0_1_108;
wire n_0_1_109;
wire n_0_1_110;
wire n_0_1_111;
wire n_0_1_112;
wire n_0_61;
wire n_0_1_113;
wire n_0_1_114;
wire n_0_1_115;
wire n_0_1_116;
wire n_0_1_117;
wire n_0_1_118;
wire n_0_62;
wire n_0_1_119;
wire n_0_1_120;
wire n_0_1_121;
wire n_0_1_122;
wire n_0_1_123;
wire n_0_1_124;
wire n_0_63;
wire n_0_1_125;
wire n_0_1_126;
wire n_0_1_127;
wire n_0_1_128;
wire n_0_1_129;
wire n_0_1_130;
wire n_0_1_131;
wire n_0_64;
wire n_0_1_132;
wire n_0_1_133;
wire n_0_1_134;
wire n_0_1_135;
wire n_0_1_136;
wire n_0_1_137;
wire n_0_1_138;
wire n_0_65;
wire n_0_1_139;
wire n_0_1_140;
wire n_0_1_141;
wire n_0_1_142;
wire n_0_1_143;
wire n_0_1_144;
wire n_0_1_145;
wire n_0_66;
wire n_0_1_146;
wire n_0_1_147;
wire n_0_1_148;
wire n_0_1_149;
wire n_0_1_150;
wire n_0_1_151;
wire n_0_1_152;
wire n_0_67;
wire n_0_1_153;
wire n_0_1_154;
wire n_0_1_155;
wire n_0_1_156;
wire n_0_1_157;
wire n_0_1_158;
wire n_0_1_159;
wire n_0_1_160;
wire n_0_68;
wire n_0_1_161;
wire n_0_1_162;
wire n_0_1_163;
wire n_0_1_164;
wire n_0_1_165;
wire n_0_1_166;
wire n_0_1_167;
wire n_0_1_168;
wire n_0_69;
wire n_0_1_169;
wire n_0_1_170;
wire n_0_1_171;
wire n_0_1_172;
wire n_0_1_173;
wire n_0_1_174;
wire n_0_1_175;
wire n_0_1_176;
wire n_0_70;
wire n_0_1_177;
wire n_0_1_178;
wire n_0_1_179;
wire n_0_1_180;
wire n_0_1_181;
wire n_0_1_182;
wire n_0_1_183;
wire n_0_1_184;
wire n_0_71;
wire n_0_1_185;
wire n_0_1_186;
wire n_0_1_187;
wire n_0_1_188;
wire n_0_1_189;
wire n_0_1_190;
wire n_0_1_191;
wire n_0_1_192;
wire n_0_72;
wire n_0_1_193;
wire n_0_1_194;
wire n_0_1_195;
wire n_0_1_196;
wire n_0_1_197;
wire n_0_1_198;
wire n_0_1_199;
wire n_0_73;
wire n_0_1_200;
wire n_0_1_201;
wire n_0_1_202;
wire n_0_1_203;
wire n_0_1_204;
wire n_0_1_205;
wire n_0_74;
wire n_0_1_206;
wire n_0_1_207;
wire n_0_1_208;
wire n_0_1_209;
wire n_0_1_210;
wire n_0_1_211;
wire n_0_75;
wire n_0_1_212;
wire n_0_1_213;
wire n_0_1_214;
wire n_0_1_215;
wire n_0_1_216;
wire n_0_1_217;
wire n_0_1_218;
wire n_0_1_219;
wire n_0_76;
wire n_0_1_220;
wire n_0_1_221;
wire n_0_1_222;
wire n_0_1_223;
wire n_0_1_224;
wire n_0_1_225;
wire n_0_1_226;
wire n_0_1_227;
wire n_0_77;
wire n_0_1_228;
wire n_0_1_229;
wire n_0_1_230;
wire n_0_1_231;
wire n_0_1_232;
wire n_0_1_233;
wire n_0_1_234;
wire n_0_1_235;
wire n_0_78;
wire n_0_1_236;
wire n_0_1_237;
wire n_0_1_238;
wire n_0_1_239;
wire n_0_1_240;
wire n_0_1_241;
wire n_0_1_242;
wire n_0_1_243;
wire n_0_79;
wire n_0_1_244;
wire n_0_1_245;
wire n_0_1_246;
wire n_0_1_247;
wire n_0_1_248;
wire n_0_1_249;
wire n_0_1_250;
wire n_0_1_251;
wire n_0_80;
wire n_0_1_252;
wire n_0_1_253;
wire n_0_1_254;
wire n_0_1_255;
wire n_0_1_256;
wire n_0_1_257;
wire n_0_1_258;
wire n_0_1_259;
wire n_0_81;
wire n_0_1_260;
wire n_0_1_261;
wire n_0_1_262;
wire n_0_1_263;
wire n_0_1_264;
wire n_0_1_265;
wire n_0_1_266;
wire n_0_1_267;
wire n_0_82;
wire n_0_1_268;
wire n_0_1_269;
wire n_0_1_270;
wire n_0_1_271;
wire n_0_1_272;
wire n_0_1_273;
wire n_0_1_274;
wire n_0_1_275;
wire n_0_1_276;
wire n_0_83;
wire n_0_1_277;
wire n_0_1_278;
wire n_0_1_279;
wire n_0_84;
wire n_0_1_280;
wire n_0_1_281;
wire n_0_1_282;
wire n_0_85;
wire n_0_1_283;
wire n_0_1_284;
wire n_0_1_285;
wire n_0_86;
wire n_0_1_286;
wire n_0_1_287;
wire n_0_1_288;
wire n_0_87;
wire n_0_1_289;
wire n_0_1_290;
wire n_0_1_291;
wire n_0_88;
wire n_0_1_292;
wire n_0_1_293;
wire n_0_1_294;
wire n_0_89;
wire n_0_1_295;
wire n_0_1_296;
wire n_0_1_297;
wire n_0_90;
wire n_0_1_298;
wire n_0_1_299;
wire n_0_1_300;
wire n_0_91;
wire n_0_1_301;
wire n_0_1_302;
wire n_0_1_303;
wire n_0_92;
wire n_0_1_304;
wire n_0_1_305;
wire n_0_1_306;
wire n_0_93;
wire n_0_1_307;
wire n_0_1_308;
wire n_0_1_309;
wire n_0_94;
wire n_0_1_310;
wire n_0_1_311;
wire n_0_1_312;
wire n_0_95;
wire n_0_1_313;
wire n_0_1_314;
wire n_0_1_315;
wire n_0_96;
wire n_0_1_316;
wire n_0_1_317;
wire n_0_1_318;
wire n_0_97;
wire n_0_1_319;
wire n_0_1_320;
wire n_0_1_321;
wire n_0_98;
wire n_0_1_322;
wire n_0_1_323;
wire n_0_1_324;
wire n_0_99;
wire n_0_1_325;
wire n_0_1_326;
wire n_0_1_327;
wire n_0_1_328;
wire n_0_100;
wire n_0_1_329;
wire n_0_1_330;
wire n_0_1_331;
wire n_0_101;
wire n_0_1_332;
wire n_0_1_333;
wire n_0_1_334;
wire n_0_102;
wire n_0_1_335;
wire n_0_1_336;
wire n_0_1_337;
wire n_0_103;
wire n_0_1_338;
wire n_0_1_339;
wire n_0_1_340;
wire n_0_104;
wire n_0_1_341;
wire n_0_1_342;
wire n_0_1_343;
wire n_0_105;
wire n_0_1_344;
wire n_0_1_345;
wire n_0_1_346;
wire n_0_106;
wire n_0_1_347;
wire n_0_1_348;
wire n_0_1_349;
wire n_0_107;
wire n_0_1_350;
wire n_0_1_351;
wire n_0_1_352;
wire n_0_1_353;
wire n_0_108;
wire n_0_1_354;
wire n_0_1_355;
wire n_0_1_356;
wire n_0_1_357;
wire n_0_109;
wire n_0_1_358;
wire n_0_1_359;
wire n_0_1_360;
wire n_0_110;
wire n_0_1_361;
wire n_0_1_362;
wire n_0_1_363;
wire n_0_111;
wire n_0_1_364;
wire n_0_1_365;
wire n_0_1_366;
wire n_0_112;
wire n_0_1_367;
wire n_0_1_368;
wire n_0_1_369;
wire n_0_113;
wire n_0_1_370;
wire n_0_1_371;
wire n_0_1_372;
wire n_0_114;
wire n_0_1_373;
wire n_0_1_374;
wire n_0_1_375;
wire n_0_1_376;
wire n_0_1_377;
wire n_0_115;
wire n_0_0;
wire \counter[4] ;
wire \counter[3] ;
wire \counter[2] ;
wire \counter[1] ;
wire \counter[0] ;
wire resetReg;
wire n_0_264;
wire n_64;
wire n_0;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire uc_0;
wire hfn_ipo_n36;
wire drc_ipo_n47;
wire drc_ipo_n48;
wire hfn_ipo_n37;
wire CTS_n_tid0_64;
wire hfn_ipo_n42;
wire hfn_ipo_n43;
wire hfn_ipo_n41;
wire hfn_ipo_n44;
wire hfn_ipo_n45;
wire hfn_ipo_n46;
wire hfn_ipo_n33;
wire hfn_ipo_n34;
wire hfn_ipo_n40;


MUX2_X1 resetReg_reg_enable_mux_0 (.Z (n_0_264), .A (resetReg), .B (n_0_129), .S (n_0_130));
DFF_X1 resetReg_reg (.Q (resetReg), .CK (CTS_n_tid0_63), .D (n_0_264));
DFF_X1 \counter_reg[0]  (.Q (\counter[0] ), .CK (n_0_0), .D (n_0_259));
DFF_X1 \counter_reg[1]  (.Q (\counter[1] ), .CK (n_0_0), .D (n_0_260));
DFF_X1 \counter_reg[2]  (.Q (\counter[2] ), .CK (n_0_0), .D (n_0_261));
DFF_X1 \counter_reg[3]  (.Q (\counter[3] ), .CK (n_0_0), .D (n_0_262));
DFF_X1 \counter_reg[4]  (.Q (\counter[4] ), .CK (n_0_0), .D (n_0_263));
CLKGATETST_X1 clk_gate_counter_reg (.GCK (n_0_0), .CK (clk_CTS_0_PP_10), .E (enable), .SE (1'b0 ));
OAI22_X1 i_0_1_573 (.ZN (n_0_115), .A1 (n_0_1_369), .A2 (hfn_ipo_n36), .B1 (n_0_1_377), .B2 (hfn_ipo_n44));
OAI221_X1 i_0_1_572 (.ZN (n_0_1_377), .A (n_0_1_375), .B1 (n_0_1_376), .B2 (hfn_ipo_n41)
    , .C1 (n_0_1_362), .C2 (n_0_1_15));
NAND2_X1 i_0_1_571 (.ZN (n_0_1_376), .A1 (n_0_1_347), .A2 (n_0_1_351));
NAND4_X1 i_0_1_570 (.ZN (n_0_1_375), .A1 (n_0_1_373), .A2 (n_0_1_374), .A3 (n_0_1_7), .A4 (n_0_1_15));
NAND3_X1 i_0_1_569 (.ZN (n_0_1_374), .A1 (n_0_1_149), .A2 (\counter[4] ), .A3 (\counter[3] ));
OAI21_X1 i_0_1_568 (.ZN (n_0_1_373), .A (n_0_1_270), .B1 (n_0_1_8), .B2 (n_0_1_9));
OAI21_X1 i_0_1_567 (.ZN (n_0_114), .A (n_0_1_372), .B1 (n_0_1_366), .B2 (hfn_ipo_n36));
OAI221_X1 i_0_1_566 (.ZN (n_0_1_372), .A (hfn_ipo_n36), .B1 (n_0_1_359), .B2 (n_0_1_15)
    , .C1 (hfn_ipo_n41), .C2 (n_0_1_371));
AOI22_X1 i_0_1_565 (.ZN (n_0_1_371), .A1 (n_0_1_370), .A2 (n_0_1_326), .B1 (n_0_1_344), .B2 (n_0_1_351));
NAND2_X1 i_0_1_564 (.ZN (n_0_1_370), .A1 (n_0_1_264), .A2 (\counter[4] ));
OAI22_X1 i_0_1_563 (.ZN (n_0_113), .A1 (n_0_1_369), .A2 (hfn_ipo_n44), .B1 (hfn_ipo_n36), .B2 (n_0_1_363));
AOI21_X1 i_0_1_562 (.ZN (n_0_1_369), .A (n_0_1_368), .B1 (hfn_ipo_n41), .B2 (n_0_1_356));
AOI221_X1 i_0_1_561 (.ZN (n_0_1_368), .A (hfn_ipo_n41), .B1 (n_0_1_367), .B2 (n_0_1_326)
    , .C1 (n_0_1_341), .C2 (n_0_1_351));
NAND2_X1 i_0_1_560 (.ZN (n_0_1_367), .A1 (n_0_1_256), .A2 (\counter[4] ));
OAI22_X1 i_0_1_559 (.ZN (n_0_112), .A1 (n_0_1_366), .A2 (hfn_ipo_n44), .B1 (n_0_1_360), .B2 (hfn_ipo_n36));
AOI21_X1 i_0_1_558 (.ZN (n_0_1_366), .A (n_0_1_365), .B1 (hfn_ipo_n41), .B2 (n_0_1_352));
AOI221_X1 i_0_1_557 (.ZN (n_0_1_365), .A (hfn_ipo_n41), .B1 (n_0_1_364), .B2 (n_0_1_326)
    , .C1 (n_0_1_338), .C2 (n_0_1_351));
NAND2_X1 i_0_1_556 (.ZN (n_0_1_364), .A1 (n_0_1_248), .A2 (\counter[4] ));
OAI22_X1 i_0_1_555 (.ZN (n_0_111), .A1 (n_0_1_357), .A2 (hfn_ipo_n36), .B1 (n_0_1_363), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_554 (.ZN (n_0_1_363), .A1 (n_0_1_348), .A2 (hfn_ipo_n41), .B1 (n_0_1_362), .B2 (n_0_1_15));
AOI22_X1 i_0_1_553 (.ZN (n_0_1_362), .A1 (n_0_1_335), .A2 (n_0_1_351), .B1 (n_0_1_361), .B2 (n_0_1_326));
NAND2_X1 i_0_1_552 (.ZN (n_0_1_361), .A1 (n_0_1_240), .A2 (\counter[4] ));
OAI22_X1 i_0_1_551 (.ZN (n_0_110), .A1 (n_0_1_353), .A2 (hfn_ipo_n36), .B1 (n_0_1_360), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_550 (.ZN (n_0_1_360), .A1 (n_0_1_345), .A2 (hfn_ipo_n41), .B1 (n_0_1_359), .B2 (n_0_1_15));
AOI22_X1 i_0_1_549 (.ZN (n_0_1_359), .A1 (n_0_1_358), .A2 (n_0_1_326), .B1 (n_0_1_332), .B2 (n_0_1_351));
NAND2_X1 i_0_1_548 (.ZN (n_0_1_358), .A1 (n_0_1_232), .A2 (\counter[4] ));
OAI22_X1 i_0_1_547 (.ZN (n_0_109), .A1 (n_0_1_349), .A2 (hfn_ipo_n36), .B1 (n_0_1_357), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_546 (.ZN (n_0_1_357), .A1 (n_0_1_342), .A2 (hfn_ipo_n41), .B1 (n_0_1_356), .B2 (n_0_1_15));
AOI21_X1 i_0_1_545 (.ZN (n_0_1_356), .A (n_0_1_355), .B1 (n_0_1_329), .B2 (n_0_1_351));
AOI21_X1 i_0_1_544 (.ZN (n_0_1_355), .A (n_0_1_354), .B1 (n_0_1_224), .B2 (\counter[4] ));
INV_X1 i_0_1_543 (.ZN (n_0_1_354), .A (n_0_1_326));
OAI22_X1 i_0_1_542 (.ZN (n_0_108), .A1 (n_0_1_346), .A2 (hfn_ipo_n36), .B1 (n_0_1_353), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_541 (.ZN (n_0_1_353), .A1 (n_0_1_339), .A2 (hfn_ipo_n41), .B1 (n_0_1_15), .B2 (n_0_1_352));
AOI22_X1 i_0_1_540 (.ZN (n_0_1_352), .A1 (n_0_1_350), .A2 (n_0_1_326), .B1 (n_0_1_325), .B2 (n_0_1_351));
NOR2_X1 i_0_1_539 (.ZN (n_0_1_351), .A1 (n_0_1_271), .A2 (n_0_1_7));
NAND2_X1 i_0_1_538 (.ZN (n_0_1_350), .A1 (n_0_1_216), .A2 (\counter[4] ));
OAI22_X1 i_0_1_537 (.ZN (n_0_107), .A1 (n_0_1_343), .A2 (hfn_ipo_n36), .B1 (n_0_1_349), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_536 (.ZN (n_0_1_349), .A1 (n_0_1_336), .A2 (hfn_ipo_n41), .B1 (n_0_1_15), .B2 (n_0_1_348));
AOI22_X1 i_0_1_535 (.ZN (n_0_1_348), .A1 (n_0_1_347), .A2 (n_0_1_326), .B1 (n_0_1_322), .B2 (drc_ipo_n47));
OR2_X1 i_0_1_534 (.ZN (n_0_1_347), .A1 (n_0_1_209), .A2 (n_0_1_8));
OAI22_X1 i_0_1_533 (.ZN (n_0_106), .A1 (n_0_1_340), .A2 (hfn_ipo_n36), .B1 (n_0_1_346), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_532 (.ZN (n_0_1_346), .A1 (n_0_1_345), .A2 (n_0_1_15), .B1 (n_0_1_333), .B2 (hfn_ipo_n41));
AOI22_X1 i_0_1_531 (.ZN (n_0_1_345), .A1 (n_0_1_319), .A2 (drc_ipo_n47), .B1 (n_0_1_344), .B2 (n_0_1_326));
OR2_X1 i_0_1_530 (.ZN (n_0_1_344), .A1 (n_0_1_203), .A2 (n_0_1_8));
OAI22_X1 i_0_1_529 (.ZN (n_0_105), .A1 (n_0_1_337), .A2 (hfn_ipo_n36), .B1 (n_0_1_343), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_528 (.ZN (n_0_1_343), .A1 (n_0_1_330), .A2 (hfn_ipo_n42), .B1 (n_0_1_342), .B2 (n_0_1_15));
AOI22_X1 i_0_1_527 (.ZN (n_0_1_342), .A1 (n_0_1_316), .A2 (drc_ipo_n47), .B1 (n_0_1_341), .B2 (n_0_1_326));
OR2_X1 i_0_1_526 (.ZN (n_0_1_341), .A1 (n_0_1_197), .A2 (n_0_1_8));
OAI22_X1 i_0_1_525 (.ZN (n_0_104), .A1 (n_0_1_334), .A2 (hfn_ipo_n36), .B1 (n_0_1_340), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_524 (.ZN (n_0_1_340), .A1 (n_0_1_339), .A2 (n_0_1_15), .B1 (n_0_1_327), .B2 (hfn_ipo_n41));
AOI22_X1 i_0_1_523 (.ZN (n_0_1_339), .A1 (n_0_1_313), .A2 (drc_ipo_n47), .B1 (n_0_1_338), .B2 (n_0_1_326));
NAND2_X1 i_0_1_522 (.ZN (n_0_1_338), .A1 (n_0_1_189), .A2 (\counter[4] ));
OAI22_X1 i_0_1_521 (.ZN (n_0_103), .A1 (n_0_1_331), .A2 (hfn_ipo_n36), .B1 (n_0_1_337), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_520 (.ZN (n_0_1_337), .A1 (n_0_1_336), .A2 (hfn_ipo_n40), .B1 (n_0_1_323), .B2 (hfn_ipo_n42));
AOI22_X1 i_0_1_519 (.ZN (n_0_1_336), .A1 (n_0_1_310), .A2 (drc_ipo_n47), .B1 (n_0_1_335), .B2 (n_0_1_326));
NAND2_X1 i_0_1_518 (.ZN (n_0_1_335), .A1 (n_0_1_181), .A2 (\counter[4] ));
OAI22_X1 i_0_1_517 (.ZN (n_0_102), .A1 (n_0_1_334), .A2 (hfn_ipo_n44), .B1 (n_0_1_328), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_516 (.ZN (n_0_1_334), .A1 (n_0_1_320), .A2 (hfn_ipo_n42), .B1 (n_0_1_333), .B2 (n_0_1_15));
AOI22_X1 i_0_1_515 (.ZN (n_0_1_333), .A1 (n_0_1_307), .A2 (drc_ipo_n47), .B1 (n_0_1_332), .B2 (n_0_1_326));
NAND2_X1 i_0_1_514 (.ZN (n_0_1_332), .A1 (n_0_1_173), .A2 (\counter[4] ));
OAI22_X1 i_0_1_513 (.ZN (n_0_101), .A1 (n_0_1_331), .A2 (hfn_ipo_n44), .B1 (n_0_1_324), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_512 (.ZN (n_0_1_331), .A1 (n_0_1_317), .A2 (hfn_ipo_n42), .B1 (n_0_1_330), .B2 (hfn_ipo_n40));
AOI22_X1 i_0_1_511 (.ZN (n_0_1_330), .A1 (n_0_1_304), .A2 (drc_ipo_n47), .B1 (n_0_1_329), .B2 (n_0_1_326));
OR2_X1 i_0_1_510 (.ZN (n_0_1_329), .A1 (n_0_1_164), .A2 (n_0_1_8));
OAI22_X1 i_0_1_509 (.ZN (n_0_100), .A1 (n_0_1_321), .A2 (hfn_ipo_n36), .B1 (n_0_1_328), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_508 (.ZN (n_0_1_328), .A1 (n_0_1_314), .A2 (hfn_ipo_n42), .B1 (n_0_1_327), .B2 (hfn_ipo_n40));
AOI22_X1 i_0_1_507 (.ZN (n_0_1_327), .A1 (n_0_1_301), .A2 (drc_ipo_n47), .B1 (n_0_1_325), .B2 (n_0_1_326));
NOR2_X2 i_0_1_506 (.ZN (n_0_1_326), .A1 (n_0_1_271), .A2 (drc_ipo_n47));
NAND2_X1 i_0_1_505 (.ZN (n_0_1_325), .A1 (n_0_1_157), .A2 (\counter[4] ));
OAI22_X1 i_0_1_504 (.ZN (n_0_99), .A1 (n_0_1_318), .A2 (hfn_ipo_n36), .B1 (n_0_1_324), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_503 (.ZN (n_0_1_324), .A1 (n_0_1_311), .A2 (hfn_ipo_n42), .B1 (n_0_1_323), .B2 (hfn_ipo_n40));
AOI22_X1 i_0_1_502 (.ZN (n_0_1_323), .A1 (n_0_1_298), .A2 (drc_ipo_n47), .B1 (n_0_1_7), .B2 (n_0_1_322));
AOI21_X1 i_0_1_501 (.ZN (n_0_1_322), .A (n_0_1_271), .B1 (n_0_1_14), .B2 (n_0_1_149));
OAI22_X1 i_0_1_500 (.ZN (n_0_98), .A1 (n_0_1_321), .A2 (hfn_ipo_n44), .B1 (n_0_1_315), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_499 (.ZN (n_0_1_321), .A1 (n_0_1_320), .A2 (hfn_ipo_n40), .B1 (n_0_1_308), .B2 (hfn_ipo_n42));
AOI22_X1 i_0_1_498 (.ZN (n_0_1_320), .A1 (n_0_1_295), .A2 (drc_ipo_n47), .B1 (n_0_1_319), .B2 (n_0_1_7));
AOI221_X2 i_0_1_497 (.ZN (n_0_1_319), .A (n_0_1_272), .B1 (n_0_1_262), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_141));
OAI22_X1 i_0_1_496 (.ZN (n_0_97), .A1 (n_0_1_318), .A2 (hfn_ipo_n44), .B1 (n_0_1_312), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_495 (.ZN (n_0_1_318), .A1 (n_0_1_305), .A2 (hfn_ipo_n42), .B1 (n_0_1_317), .B2 (hfn_ipo_n40));
AOI22_X1 i_0_1_494 (.ZN (n_0_1_317), .A1 (n_0_1_292), .A2 (drc_ipo_n47), .B1 (n_0_1_316), .B2 (n_0_1_7));
AOI221_X2 i_0_1_493 (.ZN (n_0_1_316), .A (n_0_1_272), .B1 (n_0_1_254), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_135));
OAI22_X1 i_0_1_492 (.ZN (n_0_96), .A1 (n_0_1_315), .A2 (hfn_ipo_n44), .B1 (n_0_1_309), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_491 (.ZN (n_0_1_315), .A1 (n_0_1_302), .A2 (hfn_ipo_n42), .B1 (n_0_1_314), .B2 (hfn_ipo_n40));
OAI22_X1 i_0_1_490 (.ZN (n_0_1_314), .A1 (n_0_1_289), .A2 (n_0_1_7), .B1 (n_0_1_313), .B2 (drc_ipo_n47));
AOI221_X2 i_0_1_489 (.ZN (n_0_1_313), .A (n_0_1_272), .B1 (n_0_1_246), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_128));
OAI22_X1 i_0_1_488 (.ZN (n_0_95), .A1 (n_0_1_306), .A2 (hfn_ipo_n36), .B1 (n_0_1_312), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_487 (.ZN (n_0_1_312), .A1 (n_0_1_311), .A2 (hfn_ipo_n40), .B1 (n_0_1_299), .B2 (hfn_ipo_n42));
OAI22_X1 i_0_1_486 (.ZN (n_0_1_311), .A1 (n_0_1_286), .A2 (n_0_1_7), .B1 (n_0_1_310), .B2 (drc_ipo_n47));
AOI221_X1 i_0_1_485 (.ZN (n_0_1_310), .A (n_0_1_272), .B1 (n_0_1_238), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_121));
OAI22_X1 i_0_1_484 (.ZN (n_0_94), .A1 (n_0_1_309), .A2 (hfn_ipo_n44), .B1 (n_0_1_303), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_483 (.ZN (n_0_1_309), .A1 (n_0_1_308), .A2 (hfn_ipo_n40), .B1 (n_0_1_296), .B2 (hfn_ipo_n42));
OAI22_X1 i_0_1_482 (.ZN (n_0_1_308), .A1 (n_0_1_283), .A2 (n_0_1_7), .B1 (n_0_1_307), .B2 (drc_ipo_n47));
AOI221_X1 i_0_1_481 (.ZN (n_0_1_307), .A (n_0_1_272), .B1 (n_0_1_230), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_115));
OAI22_X1 i_0_1_480 (.ZN (n_0_93), .A1 (n_0_1_306), .A2 (hfn_ipo_n44), .B1 (n_0_1_300), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_479 (.ZN (n_0_1_306), .A1 (n_0_1_305), .A2 (hfn_ipo_n40), .B1 (n_0_1_293), .B2 (hfn_ipo_n42));
AOI22_X1 i_0_1_478 (.ZN (n_0_1_305), .A1 (n_0_1_280), .A2 (drc_ipo_n47), .B1 (n_0_1_304), .B2 (n_0_1_7));
AOI221_X2 i_0_1_477 (.ZN (n_0_1_304), .A (n_0_1_272), .B1 (n_0_1_222), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_109));
OAI22_X1 i_0_1_476 (.ZN (n_0_92), .A1 (n_0_1_303), .A2 (hfn_ipo_n44), .B1 (n_0_1_297), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_475 (.ZN (n_0_1_303), .A1 (n_0_1_302), .A2 (hfn_ipo_n40), .B1 (n_0_1_290), .B2 (hfn_ipo_n42));
OAI22_X1 i_0_1_474 (.ZN (n_0_1_302), .A1 (n_0_1_277), .A2 (n_0_1_7), .B1 (n_0_1_301), .B2 (drc_ipo_n47));
AOI221_X1 i_0_1_473 (.ZN (n_0_1_301), .A (n_0_1_272), .B1 (n_0_1_214), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_101));
OAI22_X1 i_0_1_472 (.ZN (n_0_91), .A1 (n_0_1_294), .A2 (hfn_ipo_n36), .B1 (n_0_1_300), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_471 (.ZN (n_0_1_300), .A1 (n_0_1_287), .A2 (hfn_ipo_n42), .B1 (n_0_1_299), .B2 (hfn_ipo_n40));
OAI22_X1 i_0_1_470 (.ZN (n_0_1_299), .A1 (n_0_1_298), .A2 (drc_ipo_n47), .B1 (n_0_1_7), .B2 (n_0_1_274));
AOI221_X1 i_0_1_469 (.ZN (n_0_1_298), .A (n_0_1_272), .B1 (n_0_1_208), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_97));
OAI22_X1 i_0_1_468 (.ZN (n_0_90), .A1 (n_0_1_297), .A2 (hfn_ipo_n44), .B1 (n_0_1_291), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_467 (.ZN (n_0_1_297), .A1 (n_0_1_296), .A2 (hfn_ipo_n40), .B1 (n_0_1_284), .B2 (hfn_ipo_n42));
OAI22_X1 i_0_1_466 (.ZN (n_0_1_296), .A1 (n_0_1_295), .A2 (drc_ipo_n47), .B1 (n_0_1_265), .B2 (n_0_1_7));
AOI221_X1 i_0_1_465 (.ZN (n_0_1_295), .A (n_0_1_272), .B1 (n_0_1_202), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_93));
OAI22_X1 i_0_1_464 (.ZN (n_0_89), .A1 (n_0_1_294), .A2 (hfn_ipo_n43), .B1 (n_0_1_288), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_463 (.ZN (n_0_1_294), .A1 (n_0_1_281), .A2 (hfn_ipo_n42), .B1 (n_0_1_293), .B2 (hfn_ipo_n40));
OAI22_X1 i_0_1_462 (.ZN (n_0_1_293), .A1 (n_0_1_292), .A2 (drc_ipo_n47), .B1 (n_0_1_257), .B2 (n_0_1_7));
AOI221_X1 i_0_1_461 (.ZN (n_0_1_292), .A (n_0_1_272), .B1 (n_0_1_196), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_89));
OAI22_X1 i_0_1_460 (.ZN (n_0_88), .A1 (n_0_1_291), .A2 (hfn_ipo_n44), .B1 (n_0_1_285), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_459 (.ZN (n_0_1_291), .A1 (n_0_1_278), .A2 (hfn_ipo_n42), .B1 (n_0_1_290), .B2 (hfn_ipo_n40));
OAI22_X1 i_0_1_458 (.ZN (n_0_1_290), .A1 (n_0_1_289), .A2 (drc_ipo_n47), .B1 (n_0_1_249), .B2 (n_0_1_7));
AOI221_X1 i_0_1_457 (.ZN (n_0_1_289), .A (n_0_1_272), .B1 (n_0_1_187), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_82));
OAI22_X1 i_0_1_456 (.ZN (n_0_87), .A1 (n_0_1_282), .A2 (hfn_ipo_n35), .B1 (n_0_1_288), .B2 (hfn_ipo_n43));
AOI22_X1 i_0_1_455 (.ZN (n_0_1_288), .A1 (n_0_1_287), .A2 (hfn_ipo_n40), .B1 (n_0_1_275), .B2 (hfn_ipo_n42));
OAI22_X1 i_0_1_454 (.ZN (n_0_1_287), .A1 (n_0_1_286), .A2 (drc_ipo_n47), .B1 (n_0_1_241), .B2 (n_0_1_7));
AOI221_X1 i_0_1_453 (.ZN (n_0_1_286), .A (n_0_1_272), .B1 (n_0_1_179), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_78));
OAI22_X1 i_0_1_452 (.ZN (n_0_86), .A1 (n_0_1_279), .A2 (hfn_ipo_n35), .B1 (n_0_1_285), .B2 (hfn_ipo_n43));
AOI22_X1 i_0_1_451 (.ZN (n_0_1_285), .A1 (n_0_1_284), .A2 (hfn_ipo_n40), .B1 (hfn_ipo_n42), .B2 (n_0_1_266));
OAI22_X1 i_0_1_450 (.ZN (n_0_1_284), .A1 (n_0_1_283), .A2 (drc_ipo_n47), .B1 (n_0_1_233), .B2 (n_0_1_7));
AOI221_X1 i_0_1_449 (.ZN (n_0_1_283), .A (n_0_1_272), .B1 (n_0_1_171), .B2 (n_0_1_273)
    , .C1 (n_0_1_14), .C2 (n_0_1_73));
OAI22_X1 i_0_1_448 (.ZN (n_0_85), .A1 (n_0_1_282), .A2 (hfn_ipo_n43), .B1 (n_0_1_276), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_447 (.ZN (n_0_1_282), .A1 (n_0_1_281), .A2 (hfn_ipo_n40), .B1 (hfn_ipo_n42), .B2 (n_0_1_258));
OAI22_X1 i_0_1_446 (.ZN (n_0_1_281), .A1 (n_0_1_280), .A2 (drc_ipo_n47), .B1 (n_0_1_225), .B2 (n_0_1_7));
AOI221_X1 i_0_1_445 (.ZN (n_0_1_280), .A (n_0_1_272), .B1 (n_0_1_163), .B2 (n_0_1_273)
    , .C1 (n_0_1_86), .C2 (n_0_1_14));
OAI22_X1 i_0_1_444 (.ZN (n_0_84), .A1 (n_0_1_279), .A2 (hfn_ipo_n44), .B1 (n_0_1_267), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_443 (.ZN (n_0_1_279), .A1 (n_0_1_278), .A2 (hfn_ipo_n40), .B1 (n_0_1_250), .B2 (hfn_ipo_n42));
OAI22_X1 i_0_1_442 (.ZN (n_0_1_278), .A1 (n_0_1_277), .A2 (drc_ipo_n47), .B1 (n_0_1_217), .B2 (n_0_1_7));
AOI221_X1 i_0_1_441 (.ZN (n_0_1_277), .A (n_0_1_272), .B1 (n_0_1_14), .B2 (n_0_1_83)
    , .C1 (n_0_1_155), .C2 (n_0_1_273));
OAI22_X1 i_0_1_440 (.ZN (n_0_83), .A1 (n_0_1_276), .A2 (hfn_ipo_n44), .B1 (n_0_1_259), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_439 (.ZN (n_0_1_276), .A1 (n_0_1_275), .A2 (n_0_1_15), .B1 (n_0_1_242), .B2 (hfn_ipo_n41));
OAI22_X1 i_0_1_438 (.ZN (n_0_1_275), .A1 (n_0_1_274), .A2 (drc_ipo_n47), .B1 (n_0_1_103), .B2 (n_0_1_209));
AOI21_X1 i_0_1_437 (.ZN (n_0_1_274), .A (n_0_1_272), .B1 (n_0_1_149), .B2 (n_0_1_273));
NOR2_X2 i_0_1_436 (.ZN (n_0_1_273), .A1 (n_0_1_9), .A2 (\counter[4] ));
AND2_X1 i_0_1_435 (.ZN (n_0_1_272), .A1 (n_0_1_271), .A2 (n_0_1_9));
AND2_X1 i_0_1_434 (.ZN (n_0_1_271), .A1 (n_0_1_270), .A2 (n_0_1_8));
NAND2_X1 i_0_1_433 (.ZN (n_0_1_270), .A1 (n_0_1_268), .A2 (n_0_1_269));
AOI22_X1 i_0_1_432 (.ZN (n_0_1_269), .A1 (n_0_1_66), .A2 (\firstInputComplement[31] )
    , .B1 (\firstInputComplement[30] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_431 (.ZN (n_0_1_268), .A1 (n_0_1_68), .A2 (inputOne[31]), .B1 (n_0_1_70), .B2 (inputOne[30]));
OAI22_X1 i_0_1_430 (.ZN (n_0_82), .A1 (n_0_1_267), .A2 (hfn_ipo_n44), .B1 (n_0_1_251), .B2 (hfn_ipo_n36));
AOI22_X1 i_0_1_429 (.ZN (n_0_1_267), .A1 (n_0_1_234), .A2 (hfn_ipo_n42), .B1 (n_0_1_266), .B2 (n_0_1_15));
OAI22_X1 i_0_1_428 (.ZN (n_0_1_266), .A1 (n_0_1_265), .A2 (drc_ipo_n47), .B1 (n_0_1_203), .B2 (n_0_1_103));
NAND2_X1 i_0_1_427 (.ZN (n_0_1_265), .A1 (n_0_1_264), .A2 (n_0_1_8));
AOI22_X1 i_0_1_426 (.ZN (n_0_1_264), .A1 (n_0_1_263), .A2 (n_0_1_9), .B1 (n_0_1_142), .B2 (\counter[3] ));
INV_X1 i_0_1_425 (.ZN (n_0_1_263), .A (n_0_1_262));
NAND2_X1 i_0_1_424 (.ZN (n_0_1_262), .A1 (n_0_1_260), .A2 (n_0_1_261));
AOI22_X1 i_0_1_423 (.ZN (n_0_1_261), .A1 (n_0_1_66), .A2 (\firstInputComplement[30] )
    , .B1 (\firstInputComplement[29] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_422 (.ZN (n_0_1_260), .A1 (n_0_1_68), .A2 (inputOne[30]), .B1 (n_0_1_70), .B2 (inputOne[29]));
OAI22_X1 i_0_1_421 (.ZN (n_0_81), .A1 (n_0_1_243), .A2 (hfn_ipo_n35), .B1 (n_0_1_259), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_420 (.ZN (n_0_1_259), .A1 (n_0_1_226), .A2 (hfn_ipo_n41), .B1 (n_0_1_258), .B2 (n_0_1_15));
OAI22_X1 i_0_1_419 (.ZN (n_0_1_258), .A1 (n_0_1_257), .A2 (drc_ipo_n47), .B1 (n_0_1_197), .B2 (n_0_1_103));
NAND2_X1 i_0_1_418 (.ZN (n_0_1_257), .A1 (n_0_1_256), .A2 (n_0_1_8));
OAI22_X1 i_0_1_417 (.ZN (n_0_1_256), .A1 (n_0_1_255), .A2 (\counter[3] ), .B1 (n_0_1_136), .B2 (n_0_1_9));
INV_X1 i_0_1_416 (.ZN (n_0_1_255), .A (n_0_1_254));
NAND2_X1 i_0_1_415 (.ZN (n_0_1_254), .A1 (n_0_1_252), .A2 (n_0_1_253));
AOI22_X1 i_0_1_414 (.ZN (n_0_1_253), .A1 (n_0_1_68), .A2 (inputOne[29]), .B1 (\firstInputComplement[28] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_413 (.ZN (n_0_1_252), .A1 (n_0_1_66), .A2 (\firstInputComplement[29] )
    , .B1 (n_0_1_70), .B2 (inputOne[28]));
OAI22_X1 i_0_1_412 (.ZN (n_0_80), .A1 (n_0_1_235), .A2 (hfn_ipo_n36), .B1 (n_0_1_251), .B2 (hfn_ipo_n44));
AOI22_X1 i_0_1_411 (.ZN (n_0_1_251), .A1 (n_0_1_250), .A2 (n_0_1_15), .B1 (n_0_1_218), .B2 (hfn_ipo_n41));
OAI22_X1 i_0_1_410 (.ZN (n_0_1_250), .A1 (n_0_1_190), .A2 (n_0_1_7), .B1 (n_0_1_249), .B2 (drc_ipo_n47));
NAND2_X1 i_0_1_409 (.ZN (n_0_1_249), .A1 (n_0_1_248), .A2 (n_0_1_8));
AOI22_X1 i_0_1_408 (.ZN (n_0_1_248), .A1 (n_0_1_129), .A2 (\counter[3] ), .B1 (n_0_1_247), .B2 (n_0_1_9));
INV_X1 i_0_1_407 (.ZN (n_0_1_247), .A (n_0_1_246));
NAND2_X1 i_0_1_406 (.ZN (n_0_1_246), .A1 (n_0_1_244), .A2 (n_0_1_245));
AOI22_X1 i_0_1_405 (.ZN (n_0_1_245), .A1 (n_0_1_68), .A2 (inputOne[28]), .B1 (\firstInputComplement[27] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_404 (.ZN (n_0_1_244), .A1 (n_0_1_66), .A2 (\firstInputComplement[28] )
    , .B1 (n_0_1_70), .B2 (inputOne[27]));
OAI22_X1 i_0_1_403 (.ZN (n_0_79), .A1 (n_0_1_243), .A2 (hfn_ipo_n43), .B1 (n_0_1_227), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_402 (.ZN (n_0_1_243), .A1 (n_0_1_242), .A2 (n_0_1_15), .B1 (n_0_1_210), .B2 (n_0_1_193));
AOI22_X1 i_0_1_401 (.ZN (n_0_1_242), .A1 (n_0_1_182), .A2 (drc_ipo_n47), .B1 (n_0_1_241), .B2 (n_0_1_7));
NAND2_X1 i_0_1_400 (.ZN (n_0_1_241), .A1 (n_0_1_240), .A2 (n_0_1_8));
AOI22_X1 i_0_1_399 (.ZN (n_0_1_240), .A1 (n_0_1_122), .A2 (\counter[3] ), .B1 (n_0_1_239), .B2 (n_0_1_9));
INV_X1 i_0_1_398 (.ZN (n_0_1_239), .A (n_0_1_238));
NAND2_X1 i_0_1_397 (.ZN (n_0_1_238), .A1 (n_0_1_236), .A2 (n_0_1_237));
AOI22_X1 i_0_1_396 (.ZN (n_0_1_237), .A1 (n_0_1_68), .A2 (inputOne[27]), .B1 (\firstInputComplement[26] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_395 (.ZN (n_0_1_236), .A1 (n_0_1_66), .A2 (\firstInputComplement[27] )
    , .B1 (n_0_1_70), .B2 (inputOne[26]));
OAI22_X1 i_0_1_394 (.ZN (n_0_78), .A1 (n_0_1_235), .A2 (hfn_ipo_n44), .B1 (n_0_1_219), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_393 (.ZN (n_0_1_235), .A1 (n_0_1_234), .A2 (n_0_1_15), .B1 (n_0_1_204), .B2 (n_0_1_193));
AOI22_X1 i_0_1_392 (.ZN (n_0_1_234), .A1 (n_0_1_174), .A2 (drc_ipo_n47), .B1 (n_0_1_233), .B2 (n_0_1_7));
NAND2_X1 i_0_1_391 (.ZN (n_0_1_233), .A1 (n_0_1_232), .A2 (n_0_1_8));
AOI22_X1 i_0_1_390 (.ZN (n_0_1_232), .A1 (n_0_1_116), .A2 (\counter[3] ), .B1 (n_0_1_231), .B2 (n_0_1_9));
INV_X1 i_0_1_389 (.ZN (n_0_1_231), .A (n_0_1_230));
NAND2_X1 i_0_1_388 (.ZN (n_0_1_230), .A1 (n_0_1_228), .A2 (n_0_1_229));
AOI22_X1 i_0_1_387 (.ZN (n_0_1_229), .A1 (n_0_1_68), .A2 (inputOne[26]), .B1 (\firstInputComplement[25] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_386 (.ZN (n_0_1_228), .A1 (n_0_1_66), .A2 (\firstInputComplement[26] )
    , .B1 (n_0_1_70), .B2 (inputOne[25]));
OAI22_X1 i_0_1_385 (.ZN (n_0_77), .A1 (n_0_1_227), .A2 (hfn_ipo_n43), .B1 (n_0_1_211), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_384 (.ZN (n_0_1_227), .A1 (n_0_1_226), .A2 (n_0_1_15), .B1 (n_0_1_193), .B2 (n_0_1_198));
OAI22_X1 i_0_1_383 (.ZN (n_0_1_226), .A1 (n_0_1_225), .A2 (drc_ipo_n47), .B1 (n_0_1_164), .B2 (n_0_1_103));
NAND2_X1 i_0_1_382 (.ZN (n_0_1_225), .A1 (n_0_1_224), .A2 (n_0_1_8));
AOI22_X1 i_0_1_381 (.ZN (n_0_1_224), .A1 (n_0_1_110), .A2 (\counter[3] ), .B1 (n_0_1_223), .B2 (n_0_1_9));
INV_X1 i_0_1_380 (.ZN (n_0_1_223), .A (n_0_1_222));
NAND2_X1 i_0_1_379 (.ZN (n_0_1_222), .A1 (n_0_1_220), .A2 (n_0_1_221));
AOI22_X1 i_0_1_378 (.ZN (n_0_1_221), .A1 (n_0_1_66), .A2 (\firstInputComplement[25] )
    , .B1 (\firstInputComplement[24] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_377 (.ZN (n_0_1_220), .A1 (n_0_1_68), .A2 (inputOne[25]), .B1 (n_0_1_70), .B2 (inputOne[24]));
OAI22_X1 i_0_1_376 (.ZN (n_0_76), .A1 (n_0_1_219), .A2 (hfn_ipo_n44), .B1 (n_0_1_205), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_375 (.ZN (n_0_1_219), .A1 (n_0_1_191), .A2 (hfn_ipo_n41), .B1 (n_0_1_218), .B2 (n_0_1_15));
OAI22_X1 i_0_1_374 (.ZN (n_0_1_218), .A1 (n_0_1_217), .A2 (drc_ipo_n47), .B1 (n_0_1_158), .B2 (n_0_1_7));
NAND2_X1 i_0_1_373 (.ZN (n_0_1_217), .A1 (n_0_1_216), .A2 (n_0_1_8));
AOI22_X1 i_0_1_372 (.ZN (n_0_1_216), .A1 (n_0_1_102), .A2 (\counter[3] ), .B1 (n_0_1_215), .B2 (n_0_1_9));
INV_X1 i_0_1_371 (.ZN (n_0_1_215), .A (n_0_1_214));
NAND2_X1 i_0_1_370 (.ZN (n_0_1_214), .A1 (n_0_1_212), .A2 (n_0_1_213));
AOI22_X1 i_0_1_369 (.ZN (n_0_1_213), .A1 (n_0_1_66), .A2 (\firstInputComplement[24] )
    , .B1 (\firstInputComplement[23] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_368 (.ZN (n_0_1_212), .A1 (n_0_1_68), .A2 (inputOne[24]), .B1 (n_0_1_70), .B2 (inputOne[23]));
OAI22_X1 i_0_1_367 (.ZN (n_0_75), .A1 (n_0_1_211), .A2 (hfn_ipo_n43), .B1 (n_0_1_199), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_366 (.ZN (n_0_1_211), .A1 (n_0_1_183), .A2 (hfn_ipo_n41), .B1 (n_0_1_210), .B2 (n_0_1_167));
OAI22_X1 i_0_1_365 (.ZN (n_0_1_210), .A1 (n_0_1_209), .A2 (drc_ipo_n47), .B1 (n_0_1_150), .B2 (n_0_1_165));
OAI22_X1 i_0_1_364 (.ZN (n_0_1_209), .A1 (n_0_1_208), .A2 (\counter[3] ), .B1 (n_0_1_97), .B2 (n_0_1_9));
NAND2_X1 i_0_1_363 (.ZN (n_0_1_208), .A1 (n_0_1_206), .A2 (n_0_1_207));
AOI22_X1 i_0_1_362 (.ZN (n_0_1_207), .A1 (n_0_1_68), .A2 (inputOne[23]), .B1 (\firstInputComplement[22] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_361 (.ZN (n_0_1_206), .A1 (n_0_1_66), .A2 (\firstInputComplement[23] )
    , .B1 (n_0_1_70), .B2 (inputOne[22]));
OAI22_X1 i_0_1_360 (.ZN (n_0_74), .A1 (n_0_1_192), .A2 (hfn_ipo_n35), .B1 (n_0_1_205), .B2 (hfn_ipo_n43));
AOI22_X1 i_0_1_359 (.ZN (n_0_1_205), .A1 (n_0_1_175), .A2 (hfn_ipo_n41), .B1 (n_0_1_204), .B2 (n_0_1_167));
OAI22_X1 i_0_1_358 (.ZN (n_0_1_204), .A1 (n_0_1_203), .A2 (drc_ipo_n47), .B1 (n_0_1_142), .B2 (n_0_1_165));
OAI22_X1 i_0_1_357 (.ZN (n_0_1_203), .A1 (n_0_1_202), .A2 (\counter[3] ), .B1 (n_0_1_93), .B2 (n_0_1_9));
NAND2_X1 i_0_1_356 (.ZN (n_0_1_202), .A1 (n_0_1_200), .A2 (n_0_1_201));
AOI22_X1 i_0_1_355 (.ZN (n_0_1_201), .A1 (n_0_1_68), .A2 (inputOne[22]), .B1 (\firstInputComplement[21] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_354 (.ZN (n_0_1_200), .A1 (n_0_1_66), .A2 (\firstInputComplement[22] )
    , .B1 (n_0_1_70), .B2 (inputOne[21]));
OAI22_X1 i_0_1_353 (.ZN (n_0_73), .A1 (n_0_1_184), .A2 (hfn_ipo_n35), .B1 (n_0_1_199), .B2 (hfn_ipo_n43));
AOI22_X1 i_0_1_352 (.ZN (n_0_1_199), .A1 (n_0_1_166), .A2 (n_0_1_193), .B1 (n_0_1_167), .B2 (n_0_1_198));
OAI22_X1 i_0_1_351 (.ZN (n_0_1_198), .A1 (n_0_1_197), .A2 (drc_ipo_n47), .B1 (n_0_1_136), .B2 (n_0_1_165));
OAI22_X1 i_0_1_350 (.ZN (n_0_1_197), .A1 (n_0_1_196), .A2 (\counter[3] ), .B1 (n_0_1_89), .B2 (n_0_1_9));
NAND2_X1 i_0_1_349 (.ZN (n_0_1_196), .A1 (n_0_1_194), .A2 (n_0_1_195));
AOI22_X1 i_0_1_348 (.ZN (n_0_1_195), .A1 (n_0_1_68), .A2 (inputOne[21]), .B1 (\firstInputComplement[20] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_347 (.ZN (n_0_1_194), .A1 (n_0_1_66), .A2 (\firstInputComplement[21] )
    , .B1 (n_0_1_70), .B2 (inputOne[20]));
NOR2_X1 i_0_1_346 (.ZN (n_0_1_193), .A1 (n_0_1_15), .A2 (\counter[4] ));
OAI22_X1 i_0_1_345 (.ZN (n_0_72), .A1 (n_0_1_192), .A2 (hfn_ipo_n43), .B1 (n_0_1_176), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_344 (.ZN (n_0_1_192), .A1 (n_0_1_191), .A2 (n_0_1_15), .B1 (n_0_1_159), .B2 (hfn_ipo_n41));
OAI22_X1 i_0_1_343 (.ZN (n_0_1_191), .A1 (n_0_1_190), .A2 (drc_ipo_n47), .B1 (n_0_1_104), .B2 (n_0_1_129));
NAND2_X1 i_0_1_342 (.ZN (n_0_1_190), .A1 (n_0_1_189), .A2 (n_0_1_8));
AOI22_X1 i_0_1_341 (.ZN (n_0_1_189), .A1 (n_0_1_125), .A2 (\counter[3] ), .B1 (n_0_1_188), .B2 (n_0_1_9));
INV_X1 i_0_1_340 (.ZN (n_0_1_188), .A (n_0_1_187));
NAND2_X1 i_0_1_339 (.ZN (n_0_1_187), .A1 (n_0_1_185), .A2 (n_0_1_186));
AOI22_X1 i_0_1_338 (.ZN (n_0_1_186), .A1 (n_0_1_70), .A2 (inputOne[19]), .B1 (\firstInputComplement[19] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_337 (.ZN (n_0_1_185), .A1 (n_0_1_68), .A2 (inputOne[20]), .B1 (n_0_1_66), .B2 (\firstInputComplement[20] ));
OAI22_X1 i_0_1_336 (.ZN (n_0_71), .A1 (n_0_1_184), .A2 (hfn_ipo_n43), .B1 (n_0_1_168), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_335 (.ZN (n_0_1_184), .A1 (n_0_1_183), .A2 (n_0_1_15), .B1 (hfn_ipo_n41), .B2 (n_0_1_151));
OAI22_X1 i_0_1_334 (.ZN (n_0_1_183), .A1 (n_0_1_182), .A2 (drc_ipo_n47), .B1 (n_0_1_122), .B2 (n_0_1_104));
NAND2_X1 i_0_1_333 (.ZN (n_0_1_182), .A1 (n_0_1_181), .A2 (n_0_1_8));
AOI22_X1 i_0_1_332 (.ZN (n_0_1_181), .A1 (n_0_1_79), .A2 (\counter[3] ), .B1 (n_0_1_180), .B2 (n_0_1_9));
INV_X1 i_0_1_331 (.ZN (n_0_1_180), .A (n_0_1_179));
NAND2_X1 i_0_1_330 (.ZN (n_0_1_179), .A1 (n_0_1_177), .A2 (n_0_1_178));
AOI22_X1 i_0_1_329 (.ZN (n_0_1_178), .A1 (n_0_1_70), .A2 (inputOne[18]), .B1 (\firstInputComplement[18] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_328 (.ZN (n_0_1_177), .A1 (n_0_1_68), .A2 (inputOne[19]), .B1 (n_0_1_66), .B2 (\firstInputComplement[19] ));
OAI22_X1 i_0_1_327 (.ZN (n_0_70), .A1 (n_0_1_176), .A2 (hfn_ipo_n43), .B1 (n_0_1_160), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_326 (.ZN (n_0_1_176), .A1 (n_0_1_175), .A2 (n_0_1_15), .B1 (hfn_ipo_n41), .B2 (n_0_1_144));
OAI22_X1 i_0_1_325 (.ZN (n_0_1_175), .A1 (n_0_1_174), .A2 (drc_ipo_n47), .B1 (n_0_1_116), .B2 (n_0_1_104));
NAND2_X1 i_0_1_324 (.ZN (n_0_1_174), .A1 (n_0_1_173), .A2 (n_0_1_8));
AOI22_X1 i_0_1_323 (.ZN (n_0_1_173), .A1 (n_0_1_172), .A2 (n_0_1_9), .B1 (n_0_1_74), .B2 (\counter[3] ));
INV_X1 i_0_1_322 (.ZN (n_0_1_172), .A (n_0_1_171));
NAND2_X1 i_0_1_321 (.ZN (n_0_1_171), .A1 (n_0_1_169), .A2 (n_0_1_170));
AOI22_X1 i_0_1_320 (.ZN (n_0_1_170), .A1 (n_0_1_68), .A2 (inputOne[18]), .B1 (\firstInputComplement[17] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_319 (.ZN (n_0_1_169), .A1 (n_0_1_66), .A2 (\firstInputComplement[18] )
    , .B1 (n_0_1_70), .B2 (inputOne[17]));
OAI22_X1 i_0_1_318 (.ZN (n_0_69), .A1 (n_0_1_168), .A2 (hfn_ipo_n43), .B1 (n_0_1_152), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_317 (.ZN (n_0_1_168), .A1 (n_0_1_166), .A2 (n_0_1_167), .B1 (hfn_ipo_n41), .B2 (n_0_1_137));
NOR2_X1 i_0_1_316 (.ZN (n_0_1_167), .A1 (\counter[4] ), .A2 (hfn_ipo_n41));
OAI22_X1 i_0_1_315 (.ZN (n_0_1_166), .A1 (n_0_1_164), .A2 (drc_ipo_n47), .B1 (n_0_1_110), .B2 (n_0_1_165));
NAND2_X1 i_0_1_314 (.ZN (n_0_1_165), .A1 (n_0_1_9), .A2 (drc_ipo_n47));
OAI22_X1 i_0_1_313 (.ZN (n_0_1_164), .A1 (n_0_1_86), .A2 (n_0_1_9), .B1 (n_0_1_163), .B2 (\counter[3] ));
NAND2_X1 i_0_1_312 (.ZN (n_0_1_163), .A1 (n_0_1_161), .A2 (n_0_1_162));
AOI22_X1 i_0_1_311 (.ZN (n_0_1_162), .A1 (n_0_1_68), .A2 (inputOne[17]), .B1 (\firstInputComplement[16] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_310 (.ZN (n_0_1_161), .A1 (n_0_1_66), .A2 (\firstInputComplement[17] )
    , .B1 (n_0_1_70), .B2 (inputOne[16]));
OAI22_X1 i_0_1_309 (.ZN (n_0_68), .A1 (n_0_1_160), .A2 (hfn_ipo_n43), .B1 (hfn_ipo_n35), .B2 (n_0_1_145));
AOI22_X1 i_0_1_308 (.ZN (n_0_1_160), .A1 (n_0_1_159), .A2 (n_0_1_15), .B1 (hfn_ipo_n41), .B2 (n_0_1_130));
OAI22_X1 i_0_1_307 (.ZN (n_0_1_159), .A1 (n_0_1_158), .A2 (drc_ipo_n47), .B1 (n_0_1_102), .B2 (n_0_1_104));
NAND2_X1 i_0_1_306 (.ZN (n_0_1_158), .A1 (n_0_1_157), .A2 (n_0_1_8));
OAI22_X1 i_0_1_305 (.ZN (n_0_1_157), .A1 (n_0_1_156), .A2 (\counter[3] ), .B1 (n_0_1_9), .B2 (n_0_1_54));
INV_X1 i_0_1_304 (.ZN (n_0_1_156), .A (n_0_1_155));
NAND2_X1 i_0_1_303 (.ZN (n_0_1_155), .A1 (n_0_1_153), .A2 (n_0_1_154));
AOI22_X1 i_0_1_302 (.ZN (n_0_1_154), .A1 (n_0_1_68), .A2 (inputOne[16]), .B1 (\firstInputComplement[15] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_301 (.ZN (n_0_1_153), .A1 (n_0_1_66), .A2 (\firstInputComplement[16] )
    , .B1 (n_0_1_70), .B2 (inputOne[15]));
OAI22_X1 i_0_1_300 (.ZN (n_0_67), .A1 (n_0_1_138), .A2 (hfn_ipo_n35), .B1 (n_0_1_152), .B2 (hfn_ipo_n43));
AOI22_X1 i_0_1_299 (.ZN (n_0_1_152), .A1 (n_0_1_151), .A2 (hfn_ipo_n40), .B1 (n_0_1_123), .B2 (hfn_ipo_n42));
OAI22_X1 i_0_1_298 (.ZN (n_0_1_151), .A1 (n_0_1_146), .A2 (n_0_1_104), .B1 (n_0_1_150), .B2 (n_0_1_10));
INV_X1 i_0_1_297 (.ZN (n_0_1_150), .A (n_0_1_149));
NAND2_X1 i_0_1_296 (.ZN (n_0_1_149), .A1 (n_0_1_147), .A2 (n_0_1_148));
AOI22_X1 i_0_1_295 (.ZN (n_0_1_148), .A1 (n_0_1_68), .A2 (inputOne[15]), .B1 (drc_ipo_n48), .B2 (\firstInputComplement[14] ));
AOI22_X1 i_0_1_294 (.ZN (n_0_1_147), .A1 (n_0_1_66), .A2 (\firstInputComplement[15] )
    , .B1 (n_0_1_70), .B2 (inputOne[14]));
INV_X1 i_0_1_293 (.ZN (n_0_1_146), .A (n_0_1_97));
OAI22_X1 i_0_1_292 (.ZN (n_0_66), .A1 (n_0_1_145), .A2 (hfn_ipo_n43), .B1 (n_0_1_131), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_291 (.ZN (n_0_1_145), .A1 (n_0_1_144), .A2 (hfn_ipo_n40), .B1 (n_0_1_117), .B2 (hfn_ipo_n42));
OAI22_X1 i_0_1_290 (.ZN (n_0_1_144), .A1 (n_0_1_142), .A2 (n_0_1_10), .B1 (n_0_1_143), .B2 (n_0_1_104));
INV_X1 i_0_1_289 (.ZN (n_0_1_143), .A (n_0_1_93));
INV_X1 i_0_1_288 (.ZN (n_0_1_142), .A (n_0_1_141));
NAND2_X1 i_0_1_287 (.ZN (n_0_1_141), .A1 (n_0_1_139), .A2 (n_0_1_140));
AOI22_X1 i_0_1_286 (.ZN (n_0_1_140), .A1 (n_0_1_66), .A2 (\firstInputComplement[14] )
    , .B1 (\firstInputComplement[13] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_285 (.ZN (n_0_1_139), .A1 (n_0_1_68), .A2 (inputOne[14]), .B1 (n_0_1_70), .B2 (inputOne[13]));
OAI22_X1 i_0_1_284 (.ZN (n_0_65), .A1 (n_0_1_138), .A2 (hfn_ipo_n43), .B1 (n_0_1_124), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_283 (.ZN (n_0_1_138), .A1 (n_0_1_111), .A2 (hfn_ipo_n42), .B1 (n_0_1_137), .B2 (hfn_ipo_n40));
OAI22_X1 i_0_1_282 (.ZN (n_0_1_137), .A1 (n_0_1_132), .A2 (n_0_1_104), .B1 (n_0_1_136), .B2 (n_0_1_10));
INV_X1 i_0_1_281 (.ZN (n_0_1_136), .A (n_0_1_135));
NAND2_X1 i_0_1_280 (.ZN (n_0_1_135), .A1 (n_0_1_133), .A2 (n_0_1_134));
AOI22_X1 i_0_1_279 (.ZN (n_0_1_134), .A1 (n_0_1_68), .A2 (inputOne[13]), .B1 (\firstInputComplement[12] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_278 (.ZN (n_0_1_133), .A1 (n_0_1_66), .A2 (\firstInputComplement[13] )
    , .B1 (n_0_1_70), .B2 (inputOne[12]));
INV_X1 i_0_1_277 (.ZN (n_0_1_132), .A (n_0_1_89));
OAI22_X1 i_0_1_276 (.ZN (n_0_64), .A1 (n_0_1_131), .A2 (hfn_ipo_n43), .B1 (n_0_1_118), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_275 (.ZN (n_0_1_131), .A1 (n_0_1_130), .A2 (hfn_ipo_n40), .B1 (n_0_1_105), .B2 (hfn_ipo_n42));
OAI22_X1 i_0_1_274 (.ZN (n_0_1_130), .A1 (n_0_1_125), .A2 (n_0_1_104), .B1 (n_0_1_129), .B2 (n_0_1_10));
INV_X1 i_0_1_273 (.ZN (n_0_1_129), .A (n_0_1_128));
NAND2_X1 i_0_1_272 (.ZN (n_0_1_128), .A1 (n_0_1_126), .A2 (n_0_1_127));
AOI22_X1 i_0_1_271 (.ZN (n_0_1_127), .A1 (n_0_1_66), .A2 (\firstInputComplement[12] )
    , .B1 (\firstInputComplement[11] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_270 (.ZN (n_0_1_126), .A1 (n_0_1_68), .A2 (inputOne[12]), .B1 (n_0_1_70), .B2 (inputOne[11]));
INV_X1 i_0_1_269 (.ZN (n_0_1_125), .A (n_0_1_82));
OAI22_X1 i_0_1_268 (.ZN (n_0_63), .A1 (n_0_1_112), .A2 (hfn_ipo_n35), .B1 (n_0_1_124), .B2 (hfn_ipo_n43));
AOI22_X1 i_0_1_267 (.ZN (n_0_1_124), .A1 (n_0_1_123), .A2 (hfn_ipo_n40), .B1 (n_0_1_97), .B2 (n_0_1_84));
OAI22_X1 i_0_1_266 (.ZN (n_0_1_123), .A1 (n_0_1_79), .A2 (n_0_1_104), .B1 (n_0_1_122), .B2 (n_0_1_10));
INV_X1 i_0_1_265 (.ZN (n_0_1_122), .A (n_0_1_121));
NAND2_X1 i_0_1_264 (.ZN (n_0_1_121), .A1 (n_0_1_119), .A2 (n_0_1_120));
AOI22_X1 i_0_1_263 (.ZN (n_0_1_120), .A1 (n_0_1_66), .A2 (\firstInputComplement[11] )
    , .B1 (\firstInputComplement[10] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_262 (.ZN (n_0_1_119), .A1 (n_0_1_68), .A2 (inputOne[11]), .B1 (n_0_1_70), .B2 (inputOne[10]));
OAI22_X1 i_0_1_261 (.ZN (n_0_62), .A1 (n_0_1_118), .A2 (hfn_ipo_n43), .B1 (n_0_1_106), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_260 (.ZN (n_0_1_118), .A1 (n_0_1_117), .A2 (hfn_ipo_n40), .B1 (n_0_1_93), .B2 (n_0_1_84));
OAI22_X1 i_0_1_259 (.ZN (n_0_1_117), .A1 (n_0_1_116), .A2 (n_0_1_10), .B1 (n_0_1_74), .B2 (n_0_1_104));
INV_X1 i_0_1_258 (.ZN (n_0_1_116), .A (n_0_1_115));
NAND2_X1 i_0_1_257 (.ZN (n_0_1_115), .A1 (n_0_1_113), .A2 (n_0_1_114));
AOI22_X1 i_0_1_256 (.ZN (n_0_1_114), .A1 (n_0_1_66), .A2 (\firstInputComplement[10] )
    , .B1 (\firstInputComplement[9] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_255 (.ZN (n_0_1_113), .A1 (n_0_1_68), .A2 (inputOne[10]), .B1 (n_0_1_70), .B2 (inputOne[9]));
OAI22_X1 i_0_1_254 (.ZN (n_0_61), .A1 (n_0_1_112), .A2 (hfn_ipo_n43), .B1 (hfn_ipo_n35), .B2 (n_0_1_98));
AOI22_X1 i_0_1_253 (.ZN (n_0_1_112), .A1 (n_0_1_111), .A2 (hfn_ipo_n40), .B1 (n_0_1_89), .B2 (n_0_1_84));
OAI22_X1 i_0_1_252 (.ZN (n_0_1_111), .A1 (n_0_1_69), .A2 (n_0_1_104), .B1 (n_0_1_110), .B2 (n_0_1_10));
INV_X1 i_0_1_251 (.ZN (n_0_1_110), .A (n_0_1_109));
NAND2_X1 i_0_1_250 (.ZN (n_0_1_109), .A1 (n_0_1_107), .A2 (n_0_1_108));
AOI22_X1 i_0_1_249 (.ZN (n_0_1_108), .A1 (n_0_1_68), .A2 (inputOne[9]), .B1 (\firstInputComplement[8] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_248 (.ZN (n_0_1_107), .A1 (n_0_1_66), .A2 (\firstInputComplement[9] )
    , .B1 (n_0_1_70), .B2 (inputOne[8]));
OAI22_X1 i_0_1_247 (.ZN (n_0_60), .A1 (n_0_1_106), .A2 (hfn_ipo_n43), .B1 (hfn_ipo_n35), .B2 (n_0_1_94));
AOI22_X1 i_0_1_246 (.ZN (n_0_1_106), .A1 (n_0_1_105), .A2 (hfn_ipo_n40), .B1 (n_0_1_82), .B2 (n_0_1_84));
OAI22_X1 i_0_1_245 (.ZN (n_0_1_105), .A1 (n_0_1_102), .A2 (n_0_1_10), .B1 (n_0_1_54), .B2 (n_0_1_104));
OR2_X1 i_0_1_244 (.ZN (n_0_1_104), .A1 (n_0_1_103), .A2 (\counter[3] ));
NAND2_X1 i_0_1_243 (.ZN (n_0_1_103), .A1 (n_0_1_8), .A2 (drc_ipo_n47));
INV_X1 i_0_1_242 (.ZN (n_0_1_102), .A (n_0_1_101));
NAND2_X1 i_0_1_241 (.ZN (n_0_1_101), .A1 (n_0_1_99), .A2 (n_0_1_100));
AOI22_X1 i_0_1_240 (.ZN (n_0_1_100), .A1 (n_0_1_66), .A2 (\firstInputComplement[8] )
    , .B1 (\firstInputComplement[7] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_239 (.ZN (n_0_1_99), .A1 (n_0_1_68), .A2 (inputOne[8]), .B1 (n_0_1_70), .B2 (inputOne[7]));
OAI22_X1 i_0_1_238 (.ZN (n_0_59), .A1 (n_0_1_90), .A2 (hfn_ipo_n35), .B1 (n_0_1_98), .B2 (hfn_ipo_n43));
AOI22_X1 i_0_1_237 (.ZN (n_0_1_98), .A1 (n_0_1_78), .A2 (n_0_1_84), .B1 (n_0_1_97), .B2 (n_0_1_11));
NAND2_X1 i_0_1_236 (.ZN (n_0_1_97), .A1 (n_0_1_95), .A2 (n_0_1_96));
AOI22_X1 i_0_1_235 (.ZN (n_0_1_96), .A1 (n_0_1_66), .A2 (\firstInputComplement[7] )
    , .B1 (\firstInputComplement[6] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_234 (.ZN (n_0_1_95), .A1 (n_0_1_68), .A2 (inputOne[7]), .B1 (n_0_1_70), .B2 (inputOne[6]));
OAI22_X1 i_0_1_233 (.ZN (n_0_58), .A1 (n_0_1_94), .A2 (hfn_ipo_n43), .B1 (n_0_1_85), .B2 (hfn_ipo_n35));
AOI22_X1 i_0_1_232 (.ZN (n_0_1_94), .A1 (n_0_1_93), .A2 (n_0_1_11), .B1 (n_0_1_73), .B2 (n_0_1_84));
NAND2_X1 i_0_1_231 (.ZN (n_0_1_93), .A1 (n_0_1_91), .A2 (n_0_1_92));
AOI22_X1 i_0_1_230 (.ZN (n_0_1_92), .A1 (n_0_1_66), .A2 (\firstInputComplement[6] )
    , .B1 (\firstInputComplement[5] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_229 (.ZN (n_0_1_91), .A1 (n_0_1_68), .A2 (inputOne[6]), .B1 (n_0_1_70), .B2 (inputOne[5]));
OAI22_X2 i_0_1_228 (.ZN (n_0_57), .A1 (n_0_1_90), .A2 (hfn_ipo_n43), .B1 (n_0_1_79), .B2 (n_0_1_75));
AOI22_X2 i_0_1_227 (.ZN (n_0_1_90), .A1 (n_0_1_86), .A2 (n_0_1_84), .B1 (n_0_1_11), .B2 (n_0_1_89));
NAND2_X1 i_0_1_226 (.ZN (n_0_1_89), .A1 (n_0_1_87), .A2 (n_0_1_88));
AOI22_X1 i_0_1_225 (.ZN (n_0_1_88), .A1 (n_0_1_68), .A2 (inputOne[5]), .B1 (\firstInputComplement[4] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_224 (.ZN (n_0_1_87), .A1 (n_0_1_66), .A2 (\firstInputComplement[5] )
    , .B1 (n_0_1_70), .B2 (inputOne[4]));
INV_X1 i_0_1_223 (.ZN (n_0_1_86), .A (n_0_1_69));
OAI22_X1 i_0_1_222 (.ZN (n_0_56), .A1 (n_0_1_85), .A2 (hfn_ipo_n43), .B1 (n_0_1_74), .B2 (n_0_1_75));
AOI22_X1 i_0_1_221 (.ZN (n_0_1_85), .A1 (n_0_1_82), .A2 (n_0_1_11), .B1 (n_0_1_83), .B2 (n_0_1_84));
NOR2_X1 i_0_1_220 (.ZN (n_0_1_84), .A1 (n_0_1_10), .A2 (hfn_ipo_n40));
INV_X1 i_0_1_219 (.ZN (n_0_1_83), .A (n_0_1_54));
NAND2_X1 i_0_1_218 (.ZN (n_0_1_82), .A1 (n_0_1_80), .A2 (n_0_1_81));
AOI22_X1 i_0_1_217 (.ZN (n_0_1_81), .A1 (n_0_1_70), .A2 (inputOne[3]), .B1 (\firstInputComplement[3] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_216 (.ZN (n_0_1_80), .A1 (n_0_1_66), .A2 (\firstInputComplement[4] )
    , .B1 (n_0_1_68), .B2 (inputOne[4]));
OAI22_X1 i_0_1_215 (.ZN (n_0_55), .A1 (n_0_1_69), .A2 (n_0_1_75), .B1 (n_0_1_79), .B2 (hfn_ipo_n37));
INV_X1 i_0_1_214 (.ZN (n_0_1_79), .A (n_0_1_78));
NAND2_X1 i_0_1_213 (.ZN (n_0_1_78), .A1 (n_0_1_76), .A2 (n_0_1_77));
AOI22_X1 i_0_1_212 (.ZN (n_0_1_77), .A1 (n_0_1_70), .A2 (inputOne[2]), .B1 (\firstInputComplement[2] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_211 (.ZN (n_0_1_76), .A1 (n_0_1_66), .A2 (\firstInputComplement[3] )
    , .B1 (n_0_1_68), .B2 (inputOne[3]));
OAI22_X1 i_0_1_210 (.ZN (n_0_54), .A1 (n_0_1_74), .A2 (hfn_ipo_n37), .B1 (n_0_1_54), .B2 (n_0_1_75));
NAND2_X1 i_0_1_209 (.ZN (n_0_1_75), .A1 (n_0_1_11), .A2 (hfn_ipo_n43));
INV_X1 i_0_1_208 (.ZN (n_0_1_74), .A (n_0_1_73));
NAND2_X1 i_0_1_207 (.ZN (n_0_1_73), .A1 (n_0_1_71), .A2 (n_0_1_72));
AOI22_X1 i_0_1_206 (.ZN (n_0_1_72), .A1 (n_0_1_66), .A2 (\firstInputComplement[2] )
    , .B1 (\firstInputComplement[1] ), .B2 (drc_ipo_n48));
AOI22_X1 i_0_1_205 (.ZN (n_0_1_71), .A1 (n_0_1_68), .A2 (inputOne[2]), .B1 (n_0_1_70), .B2 (inputOne[1]));
INV_X2 i_0_1_204 (.ZN (n_0_1_70), .A (n_0_1_64));
NOR2_X2 i_0_1_203 (.ZN (n_0_53), .A1 (n_0_1_69), .A2 (hfn_ipo_n37));
AOI221_X1 i_0_1_202 (.ZN (n_0_1_69), .A (n_0_1_65), .B1 (n_0_1_66), .B2 (\firstInputComplement[1] )
    , .C1 (inputOne[1]), .C2 (n_0_1_68));
NOR2_X4 i_0_1_201 (.ZN (n_0_1_68), .A1 (n_0_1_52), .A2 (n_0_1_67));
INV_X1 i_0_1_200 (.ZN (n_0_1_67), .A (n_0_1_61));
NOR2_X4 i_0_1_199 (.ZN (n_0_1_66), .A1 (n_0_1_52), .A2 (n_0_1_61));
AOI21_X1 i_0_1_198 (.ZN (n_0_1_65), .A (n_0_1_53), .B1 (n_0_1_63), .B2 (n_0_1_64));
NAND3_X1 i_0_1_197 (.ZN (n_0_1_64), .A1 (n_0_1_36), .A2 (n_0_1_50), .A3 (n_0_1_61));
INV_X1 i_0_1_196 (.ZN (n_0_1_63), .A (drc_ipo_n48));
NOR3_X1 i_0_1_195 (.ZN (n_0_1_62), .A1 (n_0_1_36), .A2 (n_0_1_50), .A3 (n_0_1_61));
OAI222_X1 i_0_1_194 (.ZN (n_0_1_61), .A1 (n_0_1_59), .A2 (hfn_ipo_n35), .B1 (n_0_1_48)
    , .B2 (n_0_1_60), .C1 (n_0_1_17), .C2 (n_0_1_40));
NAND2_X1 i_0_1_193 (.ZN (n_0_1_60), .A1 (hfn_ipo_n35), .A2 (drc_ipo_n47));
AOI22_X1 i_0_1_192 (.ZN (n_0_1_59), .A1 (n_0_1_55), .A2 (n_0_1_56), .B1 (n_0_1_57), .B2 (n_0_1_58));
AOI22_X1 i_0_1_191 (.ZN (n_0_1_58), .A1 (n_0_1_22), .A2 (inputTwo[7]), .B1 (n_0_1_25), .B2 (inputTwo[19]));
AOI221_X1 i_0_1_190 (.ZN (n_0_1_57), .A (drc_ipo_n47), .B1 (n_0_1_21), .B2 (inputTwo[3])
    , .C1 (inputTwo[23]), .C2 (n_0_1_24));
AOI21_X1 i_0_1_189 (.ZN (n_0_1_56), .A (n_0_1_7), .B1 (n_0_1_24), .B2 (inputTwo[31]));
AOI222_X1 i_0_1_188 (.ZN (n_0_1_55), .A1 (inputTwo[27]), .A2 (n_0_1_25), .B1 (n_0_1_22)
    , .B2 (inputTwo[15]), .C1 (n_0_1_21), .C2 (inputTwo[11]));
NOR2_X1 i_0_1_187 (.ZN (n_0_52), .A1 (n_0_1_54), .A2 (hfn_ipo_n37));
OR2_X1 i_0_1_186 (.ZN (n_0_1_54), .A1 (n_0_1_52), .A2 (n_0_1_53));
INV_X1 i_0_1_185 (.ZN (n_0_1_53), .A (inputOne[0]));
OAI22_X1 i_0_1_184 (.ZN (n_0_1_52), .A1 (n_0_1_37), .A2 (n_0_1_51), .B1 (n_0_1_36), .B2 (n_0_1_50));
INV_X1 i_0_1_183 (.ZN (n_0_1_51), .A (n_0_1_50));
OAI221_X1 i_0_1_182 (.ZN (n_0_1_50), .A (n_0_1_41), .B1 (n_0_1_42), .B2 (n_0_1_17)
    , .C1 (n_0_1_49), .C2 (n_0_1_7));
AOI21_X1 i_0_1_181 (.ZN (n_0_1_49), .A (n_0_1_45), .B1 (hfn_ipo_n43), .B2 (n_0_1_48));
NAND2_X1 i_0_1_180 (.ZN (n_0_1_48), .A1 (n_0_1_46), .A2 (n_0_1_47));
AOI22_X1 i_0_1_179 (.ZN (n_0_1_47), .A1 (inputTwo[13]), .A2 (n_0_1_22), .B1 (n_0_1_21), .B2 (inputTwo[9]));
AOI22_X1 i_0_1_178 (.ZN (n_0_1_46), .A1 (n_0_1_24), .A2 (inputTwo[29]), .B1 (n_0_1_25), .B2 (inputTwo[25]));
AOI21_X1 i_0_1_177 (.ZN (n_0_1_45), .A (hfn_ipo_n43), .B1 (n_0_1_43), .B2 (n_0_1_44));
AOI22_X1 i_0_1_176 (.ZN (n_0_1_44), .A1 (n_0_1_22), .A2 (inputTwo[11]), .B1 (n_0_1_21), .B2 (inputTwo[7]));
AOI22_X1 i_0_1_175 (.ZN (n_0_1_43), .A1 (inputTwo[27]), .A2 (n_0_1_24), .B1 (n_0_1_25), .B2 (inputTwo[23]));
AOI222_X1 i_0_1_174 (.ZN (n_0_1_42), .A1 (n_0_1_24), .A2 (inputTwo[19]), .B1 (n_0_1_22)
    , .B2 (inputTwo[3]), .C1 (n_0_1_25), .C2 (inputTwo[15]));
NAND3_X1 i_0_1_173 (.ZN (n_0_1_41), .A1 (n_0_1_40), .A2 (n_0_1_7), .A3 (hfn_ipo_n43));
NAND2_X1 i_0_1_172 (.ZN (n_0_1_40), .A1 (n_0_1_38), .A2 (n_0_1_39));
AOI22_X1 i_0_1_171 (.ZN (n_0_1_39), .A1 (n_0_1_24), .A2 (inputTwo[21]), .B1 (n_0_1_21), .B2 (inputTwo[1]));
AOI22_X1 i_0_1_170 (.ZN (n_0_1_38), .A1 (n_0_1_25), .A2 (inputTwo[17]), .B1 (n_0_1_22), .B2 (inputTwo[5]));
INV_X2 i_0_1_169 (.ZN (n_0_1_37), .A (n_0_1_36));
AOI221_X2 i_0_1_168 (.ZN (n_0_1_36), .A (n_0_1_31), .B1 (n_0_1_32), .B2 (n_0_1_33)
    , .C1 (n_0_1_34), .C2 (n_0_1_35));
AOI222_X1 i_0_1_167 (.ZN (n_0_1_35), .A1 (n_0_1_25), .A2 (inputTwo[16]), .B1 (n_0_1_22)
    , .B2 (inputTwo[4]), .C1 (n_0_1_21), .C2 (inputTwo[0]));
AOI21_X1 i_0_1_166 (.ZN (n_0_1_34), .A (n_0_1_17), .B1 (n_0_1_24), .B2 (inputTwo[20]));
AOI222_X1 i_0_1_165 (.ZN (n_0_1_33), .A1 (n_0_1_25), .A2 (inputTwo[18]), .B1 (n_0_1_22)
    , .B2 (inputTwo[6]), .C1 (n_0_1_21), .C2 (inputTwo[2]));
AOI211_X1 i_0_1_164 (.ZN (n_0_1_32), .A (drc_ipo_n47), .B (hfn_ipo_n35), .C1 (n_0_1_24), .C2 (inputTwo[22]));
AOI21_X2 i_0_1_163 (.ZN (n_0_1_31), .A (n_0_1_7), .B1 (n_0_1_27), .B2 (n_0_1_30));
NAND3_X1 i_0_1_162 (.ZN (n_0_1_30), .A1 (n_0_1_28), .A2 (n_0_1_29), .A3 (hfn_ipo_n43));
AOI22_X1 i_0_1_161 (.ZN (n_0_1_29), .A1 (n_0_1_22), .A2 (inputTwo[14]), .B1 (n_0_1_21), .B2 (inputTwo[10]));
AOI22_X1 i_0_1_160 (.ZN (n_0_1_28), .A1 (inputTwo[30]), .A2 (n_0_1_24), .B1 (n_0_1_25), .B2 (inputTwo[26]));
NAND2_X1 i_0_1_159 (.ZN (n_0_1_27), .A1 (n_0_1_23), .A2 (n_0_1_26));
AOI22_X1 i_0_1_158 (.ZN (n_0_1_26), .A1 (inputTwo[28]), .A2 (n_0_1_24), .B1 (n_0_1_25), .B2 (inputTwo[24]));
NOR2_X1 i_0_1_157 (.ZN (n_0_1_25), .A1 (n_0_1_9), .A2 (hfn_ipo_n41));
NOR2_X1 i_0_1_156 (.ZN (n_0_1_24), .A1 (n_0_1_9), .A2 (n_0_1_15));
AOI221_X1 i_0_1_155 (.ZN (n_0_1_23), .A (hfn_ipo_n43), .B1 (n_0_1_21), .B2 (inputTwo[8])
    , .C1 (n_0_1_22), .C2 (inputTwo[12]));
NOR2_X1 i_0_1_154 (.ZN (n_0_1_22), .A1 (n_0_1_15), .A2 (\counter[3] ));
NOR2_X1 i_0_1_153 (.ZN (n_0_1_21), .A1 (\counter[3] ), .A2 (hfn_ipo_n41));
AND2_X1 i_0_1_152 (.ZN (n_0_129), .A1 (enable), .A2 (reset));
INV_X1 i_0_1_151 (.ZN (n_0_130), .A (hfn_ipo_n33));
AOI221_X1 i_0_1_150 (.ZN (n_0_263), .A (n_0_1_18), .B1 (n_0_1_20), .B2 (n_0_1_8), .C1 (n_0_1_2), .C2 (\counter[4] ));
INV_X1 i_0_1_149 (.ZN (n_0_1_20), .A (n_0_1_2));
AND2_X1 i_0_1_148 (.ZN (n_0_262), .A1 (n_0_1_19), .A2 (n_0_1_5));
AND2_X1 i_0_1_147 (.ZN (n_0_261), .A1 (n_0_1_19), .A2 (n_0_1_4));
AND2_X1 i_0_1_146 (.ZN (n_0_260), .A1 (n_0_1_19), .A2 (n_0_1_3));
INV_X1 i_0_1_145 (.ZN (n_0_1_19), .A (n_0_1_18));
NOR2_X1 i_0_1_144 (.ZN (n_0_259), .A1 (n_0_1_18), .A2 (hfn_ipo_n43));
OAI21_X1 i_0_1_143 (.ZN (n_0_1_18), .A (hfn_ipo_n33), .B1 (n_0_1_16), .B2 (n_0_1_17));
NAND2_X1 i_0_1_142 (.ZN (n_0_1_17), .A1 (n_0_1_7), .A2 (hfn_ipo_n35));
NAND3_X1 i_0_1_141 (.ZN (n_0_1_16), .A1 (n_0_1_14), .A2 (enable), .A3 (n_0_1_15));
INV_X2 i_0_1_140 (.ZN (n_0_1_15), .A (hfn_ipo_n42));
NOR2_X2 i_0_1_139 (.ZN (n_0_1_14), .A1 (n_0_1_8), .A2 (\counter[3] ));
AND2_X1 i_0_1_138 (.ZN (n_0_258), .A1 (n_0_1_13), .A2 (finalResult[63]));
AND2_X1 i_0_1_137 (.ZN (n_0_257), .A1 (n_0_1_13), .A2 (finalResult[62]));
AND2_X1 i_0_1_136 (.ZN (n_0_256), .A1 (n_0_1_13), .A2 (finalResult[61]));
AND2_X1 i_0_1_135 (.ZN (n_0_255), .A1 (n_0_1_13), .A2 (finalResult[60]));
AND2_X1 i_0_1_134 (.ZN (n_0_254), .A1 (n_0_1_13), .A2 (finalResult[59]));
AND2_X1 i_0_1_133 (.ZN (n_0_253), .A1 (n_0_1_13), .A2 (finalResult[58]));
AND2_X1 i_0_1_132 (.ZN (n_0_252), .A1 (n_0_1_13), .A2 (finalResult[57]));
AND2_X1 i_0_1_131 (.ZN (n_0_251), .A1 (n_0_1_13), .A2 (finalResult[56]));
AND2_X1 i_0_1_130 (.ZN (n_0_250), .A1 (n_0_1_13), .A2 (finalResult[55]));
AND2_X1 i_0_1_129 (.ZN (n_0_249), .A1 (n_0_1_13), .A2 (finalResult[54]));
AND2_X1 i_0_1_128 (.ZN (n_0_248), .A1 (hfn_ipo_n37), .A2 (finalResult[53]));
AND2_X1 i_0_1_127 (.ZN (n_0_247), .A1 (n_0_1_13), .A2 (finalResult[52]));
AND2_X1 i_0_1_126 (.ZN (n_0_246), .A1 (hfn_ipo_n37), .A2 (finalResult[51]));
AND2_X1 i_0_1_125 (.ZN (n_0_245), .A1 (hfn_ipo_n37), .A2 (finalResult[50]));
AND2_X1 i_0_1_124 (.ZN (n_0_244), .A1 (hfn_ipo_n37), .A2 (finalResult[49]));
AND2_X1 i_0_1_123 (.ZN (n_0_243), .A1 (hfn_ipo_n37), .A2 (finalResult[48]));
AND2_X1 i_0_1_122 (.ZN (n_0_242), .A1 (hfn_ipo_n37), .A2 (finalResult[47]));
AND2_X1 i_0_1_121 (.ZN (n_0_241), .A1 (hfn_ipo_n37), .A2 (finalResult[46]));
AND2_X1 i_0_1_120 (.ZN (n_0_240), .A1 (hfn_ipo_n37), .A2 (finalResult[45]));
AND2_X1 i_0_1_119 (.ZN (n_0_239), .A1 (hfn_ipo_n37), .A2 (finalResult[44]));
AND2_X1 i_0_1_118 (.ZN (n_0_238), .A1 (hfn_ipo_n37), .A2 (finalResult[43]));
AND2_X1 i_0_1_117 (.ZN (n_0_237), .A1 (hfn_ipo_n37), .A2 (finalResult[42]));
AND2_X1 i_0_1_116 (.ZN (n_0_236), .A1 (hfn_ipo_n37), .A2 (finalResult[41]));
AND2_X1 i_0_1_115 (.ZN (n_0_235), .A1 (hfn_ipo_n37), .A2 (finalResult[40]));
AND2_X1 i_0_1_114 (.ZN (n_0_234), .A1 (hfn_ipo_n37), .A2 (finalResult[39]));
AND2_X1 i_0_1_113 (.ZN (n_0_233), .A1 (hfn_ipo_n37), .A2 (finalResult[38]));
AND2_X1 i_0_1_112 (.ZN (n_0_232), .A1 (hfn_ipo_n37), .A2 (finalResult[37]));
AND2_X1 i_0_1_111 (.ZN (n_0_231), .A1 (hfn_ipo_n37), .A2 (finalResult[36]));
AND2_X1 i_0_1_110 (.ZN (n_0_230), .A1 (hfn_ipo_n37), .A2 (finalResult[35]));
AND2_X1 i_0_1_109 (.ZN (n_0_229), .A1 (hfn_ipo_n37), .A2 (finalResult[34]));
AND2_X1 i_0_1_108 (.ZN (n_0_228), .A1 (hfn_ipo_n37), .A2 (finalResult[33]));
AND2_X1 i_0_1_107 (.ZN (n_0_227), .A1 (hfn_ipo_n37), .A2 (finalResult[32]));
AND2_X1 i_0_1_106 (.ZN (n_0_226), .A1 (n_0_1_13), .A2 (finalResult[31]));
AND2_X1 i_0_1_105 (.ZN (n_0_225), .A1 (n_0_1_13), .A2 (finalResult[30]));
AND2_X1 i_0_1_104 (.ZN (n_0_224), .A1 (n_0_1_13), .A2 (finalResult[29]));
AND2_X1 i_0_1_103 (.ZN (n_0_223), .A1 (n_0_1_13), .A2 (finalResult[28]));
AND2_X1 i_0_1_102 (.ZN (n_0_222), .A1 (n_0_1_13), .A2 (finalResult[27]));
AND2_X1 i_0_1_101 (.ZN (n_0_221), .A1 (n_0_1_13), .A2 (finalResult[26]));
AND2_X1 i_0_1_100 (.ZN (n_0_220), .A1 (n_0_1_13), .A2 (finalResult[25]));
AND2_X1 i_0_1_99 (.ZN (n_0_219), .A1 (n_0_1_13), .A2 (finalResult[24]));
AND2_X1 i_0_1_98 (.ZN (n_0_218), .A1 (n_0_1_13), .A2 (finalResult[23]));
AND2_X1 i_0_1_97 (.ZN (n_0_217), .A1 (n_0_1_13), .A2 (finalResult[22]));
AND2_X1 i_0_1_96 (.ZN (n_0_216), .A1 (hfn_ipo_n37), .A2 (finalResult[21]));
AND2_X1 i_0_1_95 (.ZN (n_0_215), .A1 (hfn_ipo_n37), .A2 (finalResult[20]));
AND2_X1 i_0_1_94 (.ZN (n_0_214), .A1 (hfn_ipo_n37), .A2 (finalResult[19]));
AND2_X1 i_0_1_93 (.ZN (n_0_213), .A1 (hfn_ipo_n37), .A2 (finalResult[18]));
AND2_X1 i_0_1_92 (.ZN (n_0_212), .A1 (hfn_ipo_n37), .A2 (finalResult[17]));
AND2_X1 i_0_1_91 (.ZN (n_0_211), .A1 (n_0_1_13), .A2 (finalResult[16]));
AND2_X1 i_0_1_90 (.ZN (n_0_210), .A1 (hfn_ipo_n37), .A2 (finalResult[15]));
AND2_X1 i_0_1_89 (.ZN (n_0_209), .A1 (hfn_ipo_n37), .A2 (finalResult[14]));
AND2_X1 i_0_1_88 (.ZN (n_0_208), .A1 (hfn_ipo_n37), .A2 (finalResult[13]));
AND2_X1 i_0_1_87 (.ZN (n_0_207), .A1 (hfn_ipo_n37), .A2 (finalResult[12]));
AND2_X1 i_0_1_86 (.ZN (n_0_206), .A1 (hfn_ipo_n37), .A2 (finalResult[11]));
AND2_X1 i_0_1_85 (.ZN (n_0_205), .A1 (hfn_ipo_n37), .A2 (finalResult[10]));
AND2_X1 i_0_1_84 (.ZN (n_0_204), .A1 (hfn_ipo_n37), .A2 (finalResult[9]));
AND2_X1 i_0_1_83 (.ZN (n_0_203), .A1 (hfn_ipo_n37), .A2 (finalResult[8]));
AND2_X1 i_0_1_82 (.ZN (n_0_202), .A1 (hfn_ipo_n37), .A2 (finalResult[7]));
AND2_X1 i_0_1_81 (.ZN (n_0_201), .A1 (hfn_ipo_n37), .A2 (finalResult[6]));
AND2_X1 i_0_1_80 (.ZN (n_0_200), .A1 (hfn_ipo_n37), .A2 (finalResult[5]));
AND2_X1 i_0_1_79 (.ZN (n_0_199), .A1 (hfn_ipo_n37), .A2 (finalResult[4]));
AND2_X1 i_0_1_78 (.ZN (n_0_198), .A1 (hfn_ipo_n37), .A2 (finalResult[3]));
AND2_X1 i_0_1_77 (.ZN (n_0_197), .A1 (hfn_ipo_n37), .A2 (finalResult[2]));
AND2_X1 i_0_1_76 (.ZN (n_0_196), .A1 (hfn_ipo_n37), .A2 (finalResult[1]));
AND2_X1 i_0_1_75 (.ZN (n_0_195), .A1 (hfn_ipo_n37), .A2 (finalResult[0]));
NAND2_X1 i_0_1_74 (.ZN (n_0_1_13), .A1 (n_0_1_11), .A2 (hfn_ipo_n35));
INV_X1 i_0_1_73 (.ZN (n_0_1_12), .A (hfn_ipo_n44));
NOR2_X1 i_0_1_72 (.ZN (n_0_1_11), .A1 (n_0_1_10), .A2 (hfn_ipo_n42));
NAND3_X1 i_0_1_71 (.ZN (n_0_1_10), .A1 (n_0_1_7), .A2 (n_0_1_8), .A3 (n_0_1_9));
INV_X1 i_0_1_70 (.ZN (n_0_1_9), .A (\counter[3] ));
INV_X1 i_0_1_69 (.ZN (n_0_1_8), .A (\counter[4] ));
INV_X2 i_0_1_68 (.ZN (n_0_1_7), .A (drc_ipo_n47));
AND2_X1 i_0_1_67 (.ZN (n_0_194), .A1 (hfn_ipo_n33), .A2 (n_0_128));
AND2_X1 i_0_1_66 (.ZN (n_0_193), .A1 (hfn_ipo_n33), .A2 (n_0_127));
AND2_X1 i_0_1_65 (.ZN (n_0_192), .A1 (hfn_ipo_n33), .A2 (n_0_126));
AND2_X1 i_0_1_64 (.ZN (n_0_191), .A1 (hfn_ipo_n33), .A2 (n_0_125));
AND2_X1 i_0_1_63 (.ZN (n_0_190), .A1 (hfn_ipo_n33), .A2 (n_0_124));
AND2_X1 i_0_1_62 (.ZN (n_0_189), .A1 (hfn_ipo_n33), .A2 (n_0_123));
AND2_X1 i_0_1_61 (.ZN (n_0_188), .A1 (hfn_ipo_n33), .A2 (n_0_122));
AND2_X1 i_0_1_60 (.ZN (n_0_187), .A1 (hfn_ipo_n33), .A2 (n_0_121));
AND2_X1 i_0_1_59 (.ZN (n_0_186), .A1 (hfn_ipo_n33), .A2 (n_0_120));
AND2_X1 i_0_1_58 (.ZN (n_0_185), .A1 (hfn_ipo_n33), .A2 (n_0_119));
AND2_X1 i_0_1_57 (.ZN (n_0_184), .A1 (hfn_ipo_n34), .A2 (n_0_118));
AND2_X1 i_0_1_56 (.ZN (n_0_183), .A1 (hfn_ipo_n33), .A2 (n_0_117));
AND2_X1 i_0_1_55 (.ZN (n_0_182), .A1 (hfn_ipo_n34), .A2 (n_0_116));
AND2_X1 i_0_1_54 (.ZN (n_0_181), .A1 (hfn_ipo_n34), .A2 (n_0_51));
AND2_X1 i_0_1_53 (.ZN (n_0_180), .A1 (hfn_ipo_n34), .A2 (n_0_50));
AND2_X1 i_0_1_52 (.ZN (n_0_179), .A1 (hfn_ipo_n34), .A2 (n_0_49));
AND2_X1 i_0_1_51 (.ZN (n_0_178), .A1 (hfn_ipo_n34), .A2 (n_0_48));
AND2_X1 i_0_1_50 (.ZN (n_0_177), .A1 (hfn_ipo_n34), .A2 (n_0_47));
AND2_X1 i_0_1_49 (.ZN (n_0_176), .A1 (hfn_ipo_n34), .A2 (n_0_46));
AND2_X1 i_0_1_48 (.ZN (n_0_175), .A1 (hfn_ipo_n34), .A2 (n_0_45));
AND2_X1 i_0_1_47 (.ZN (n_0_174), .A1 (hfn_ipo_n34), .A2 (n_0_44));
AND2_X1 i_0_1_46 (.ZN (n_0_173), .A1 (hfn_ipo_n34), .A2 (n_0_43));
AND2_X1 i_0_1_45 (.ZN (n_0_172), .A1 (hfn_ipo_n34), .A2 (n_0_42));
AND2_X1 i_0_1_44 (.ZN (n_0_171), .A1 (hfn_ipo_n34), .A2 (n_0_41));
AND2_X1 i_0_1_43 (.ZN (n_0_170), .A1 (hfn_ipo_n34), .A2 (n_0_40));
AND2_X1 i_0_1_42 (.ZN (n_0_169), .A1 (hfn_ipo_n34), .A2 (n_0_39));
AND2_X1 i_0_1_41 (.ZN (n_0_168), .A1 (hfn_ipo_n34), .A2 (n_0_38));
AND2_X1 i_0_1_40 (.ZN (n_0_167), .A1 (hfn_ipo_n34), .A2 (n_0_37));
AND2_X1 i_0_1_39 (.ZN (n_0_166), .A1 (hfn_ipo_n34), .A2 (n_0_36));
AND2_X1 i_0_1_38 (.ZN (n_0_165), .A1 (hfn_ipo_n34), .A2 (n_0_35));
AND2_X1 i_0_1_37 (.ZN (n_0_164), .A1 (hfn_ipo_n34), .A2 (n_0_34));
AND2_X1 i_0_1_36 (.ZN (n_0_163), .A1 (hfn_ipo_n33), .A2 (n_0_33));
AND2_X1 i_0_1_35 (.ZN (n_0_162), .A1 (hfn_ipo_n33), .A2 (n_0_32));
AND2_X1 i_0_1_34 (.ZN (n_0_161), .A1 (hfn_ipo_n33), .A2 (n_0_31));
AND2_X1 i_0_1_33 (.ZN (n_0_160), .A1 (hfn_ipo_n33), .A2 (n_0_30));
AND2_X1 i_0_1_32 (.ZN (n_0_159), .A1 (hfn_ipo_n33), .A2 (n_0_29));
AND2_X1 i_0_1_31 (.ZN (n_0_158), .A1 (hfn_ipo_n33), .A2 (n_0_28));
AND2_X1 i_0_1_30 (.ZN (n_0_157), .A1 (hfn_ipo_n33), .A2 (n_0_27));
AND2_X1 i_0_1_29 (.ZN (n_0_156), .A1 (hfn_ipo_n33), .A2 (n_0_26));
AND2_X1 i_0_1_28 (.ZN (n_0_155), .A1 (hfn_ipo_n33), .A2 (n_0_25));
AND2_X1 i_0_1_27 (.ZN (n_0_154), .A1 (hfn_ipo_n33), .A2 (n_0_24));
AND2_X1 i_0_1_26 (.ZN (n_0_153), .A1 (hfn_ipo_n33), .A2 (n_0_23));
AND2_X1 i_0_1_25 (.ZN (n_0_152), .A1 (hfn_ipo_n33), .A2 (n_0_22));
AND2_X1 i_0_1_24 (.ZN (n_0_151), .A1 (hfn_ipo_n33), .A2 (n_0_21));
AND2_X1 i_0_1_23 (.ZN (n_0_150), .A1 (hfn_ipo_n33), .A2 (n_0_20));
AND2_X1 i_0_1_22 (.ZN (n_0_149), .A1 (hfn_ipo_n33), .A2 (n_0_19));
AND2_X1 i_0_1_21 (.ZN (n_0_148), .A1 (hfn_ipo_n33), .A2 (n_0_18));
AND2_X1 i_0_1_20 (.ZN (n_0_147), .A1 (hfn_ipo_n33), .A2 (n_0_17));
AND2_X1 i_0_1_19 (.ZN (n_0_146), .A1 (hfn_ipo_n33), .A2 (n_0_16));
AND2_X1 i_0_1_18 (.ZN (n_0_145), .A1 (hfn_ipo_n33), .A2 (n_0_15));
AND2_X1 i_0_1_17 (.ZN (n_0_144), .A1 (hfn_ipo_n33), .A2 (n_0_14));
AND2_X1 i_0_1_16 (.ZN (n_0_143), .A1 (hfn_ipo_n33), .A2 (n_0_13));
AND2_X1 i_0_1_15 (.ZN (n_0_142), .A1 (hfn_ipo_n33), .A2 (n_0_12));
AND2_X1 i_0_1_14 (.ZN (n_0_141), .A1 (hfn_ipo_n33), .A2 (n_0_11));
AND2_X1 i_0_1_13 (.ZN (n_0_140), .A1 (hfn_ipo_n33), .A2 (n_0_10));
AND2_X1 i_0_1_12 (.ZN (n_0_139), .A1 (hfn_ipo_n33), .A2 (n_0_9));
AND2_X1 i_0_1_11 (.ZN (n_0_138), .A1 (hfn_ipo_n33), .A2 (n_0_8));
AND2_X1 i_0_1_10 (.ZN (n_0_137), .A1 (hfn_ipo_n33), .A2 (n_0_7));
AND2_X1 i_0_1_9 (.ZN (n_0_136), .A1 (hfn_ipo_n33), .A2 (n_0_6));
AND2_X1 i_0_1_8 (.ZN (n_0_135), .A1 (hfn_ipo_n33), .A2 (n_0_5));
AND2_X1 i_0_1_7 (.ZN (n_0_134), .A1 (hfn_ipo_n33), .A2 (n_0_4));
AND2_X1 i_0_1_6 (.ZN (n_0_133), .A1 (hfn_ipo_n33), .A2 (n_0_3));
AND2_X1 i_0_1_5 (.ZN (n_0_132), .A1 (hfn_ipo_n33), .A2 (n_0_2));
AND2_X1 i_0_1_4 (.ZN (n_0_131), .A1 (hfn_ipo_n33), .A2 (n_0_1));
OAI21_X1 i_0_1_3 (.ZN (n_0_1_6), .A (enable), .B1 (resetReg), .B2 (reset));
HA_X1 i_0_1_2 (.CO (n_0_1_2), .S (n_0_1_5), .A (\counter[3] ), .B (n_0_1_1));
HA_X1 i_0_1_1 (.CO (n_0_1_1), .S (n_0_1_4), .A (drc_ipo_n47), .B (n_0_1_0));
HA_X1 i_0_1_0 (.CO (n_0_1_0), .S (n_0_1_3), .A (hfn_ipo_n41), .B (hfn_ipo_n43));
datapath__0_10 i_0_200 (.p_1 ({n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, 
    n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_51, n_0_50, 
    n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, 
    n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, 
    n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, 
    n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, 
    n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1}), .finalResult ({
    n_0_258, n_0_257, n_0_256, n_0_255, n_0_254, n_0_253, n_0_252, n_0_251, n_0_250, 
    n_0_249, n_0_248, n_0_247, n_0_246, n_0_245, n_0_244, n_0_243, n_0_242, n_0_241, 
    n_0_240, n_0_239, n_0_238, n_0_237, n_0_236, n_0_235, n_0_234, n_0_233, n_0_232, 
    n_0_231, n_0_230, n_0_229, n_0_228, n_0_227, n_0_226, n_0_225, n_0_224, n_0_223, 
    n_0_222, n_0_221, n_0_220, n_0_219, n_0_218, n_0_217, n_0_216, n_0_215, n_0_214, 
    n_0_213, n_0_212, n_0_211, n_0_210, n_0_209, n_0_208, n_0_207, n_0_206, n_0_205, 
    n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, n_0_199, n_0_198, n_0_197, n_0_196, 
    n_0_195}), .p_0 ({n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, 
    n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, 
    n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, 
    n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, 
    n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, 
    n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, 
    n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52}));
DFF_X1 \finalResult_reg[0]  (.Q (n_64), .CK (CTS_n_tid0_64), .D (n_0_131));
DFF_X1 \finalResult_reg[1]  (.Q (n_63), .CK (CTS_n_tid0_64), .D (n_0_132));
DFF_X1 \finalResult_reg[2]  (.Q (n_62), .CK (CTS_n_tid0_64), .D (n_0_133));
DFF_X1 \finalResult_reg[3]  (.Q (n_61), .CK (CTS_n_tid0_64), .D (n_0_134));
DFF_X1 \finalResult_reg[4]  (.Q (n_60), .CK (CTS_n_tid0_64), .D (n_0_135));
DFF_X1 \finalResult_reg[5]  (.Q (n_59), .CK (CTS_n_tid0_64), .D (n_0_136));
DFF_X1 \finalResult_reg[6]  (.Q (n_58), .CK (CTS_n_tid0_64), .D (n_0_137));
DFF_X1 \finalResult_reg[7]  (.Q (n_57), .CK (CTS_n_tid0_64), .D (n_0_138));
DFF_X1 \finalResult_reg[8]  (.Q (n_56), .CK (CTS_n_tid0_64), .D (n_0_139));
DFF_X1 \finalResult_reg[9]  (.Q (n_55), .CK (CTS_n_tid0_64), .D (n_0_140));
DFF_X1 \finalResult_reg[10]  (.Q (n_54), .CK (CTS_n_tid0_64), .D (n_0_141));
DFF_X1 \finalResult_reg[11]  (.Q (n_53), .CK (CTS_n_tid0_64), .D (n_0_142));
DFF_X1 \finalResult_reg[12]  (.Q (n_52), .CK (CTS_n_tid0_64), .D (n_0_143));
DFF_X1 \finalResult_reg[13]  (.Q (n_51), .CK (CTS_n_tid0_64), .D (n_0_144));
DFF_X1 \finalResult_reg[14]  (.Q (n_50), .CK (CTS_n_tid0_64), .D (n_0_145));
DFF_X1 \finalResult_reg[15]  (.Q (n_49), .CK (CTS_n_tid0_64), .D (n_0_146));
DFF_X1 \finalResult_reg[16]  (.Q (n_48), .CK (CTS_n_tid0_63), .D (n_0_147));
DFF_X1 \finalResult_reg[17]  (.Q (n_47), .CK (CTS_n_tid0_63), .D (n_0_148));
DFF_X1 \finalResult_reg[18]  (.Q (n_46), .CK (CTS_n_tid0_63), .D (n_0_149));
DFF_X1 \finalResult_reg[19]  (.Q (n_45), .CK (CTS_n_tid0_63), .D (n_0_150));
DFF_X1 \finalResult_reg[20]  (.Q (n_44), .CK (CTS_n_tid0_63), .D (n_0_151));
DFF_X1 \finalResult_reg[21]  (.Q (n_43), .CK (CTS_n_tid0_63), .D (n_0_152));
DFF_X1 \finalResult_reg[22]  (.Q (n_42), .CK (CTS_n_tid0_63), .D (n_0_153));
DFF_X1 \finalResult_reg[23]  (.Q (n_41), .CK (CTS_n_tid0_63), .D (n_0_154));
DFF_X1 \finalResult_reg[24]  (.Q (n_40), .CK (CTS_n_tid0_63), .D (n_0_155));
DFF_X1 \finalResult_reg[25]  (.Q (n_39), .CK (CTS_n_tid0_63), .D (n_0_156));
DFF_X1 \finalResult_reg[26]  (.Q (n_38), .CK (CTS_n_tid0_63), .D (n_0_157));
DFF_X1 \finalResult_reg[27]  (.Q (n_37), .CK (CTS_n_tid0_63), .D (n_0_158));
DFF_X1 \finalResult_reg[28]  (.Q (n_36), .CK (CTS_n_tid0_63), .D (n_0_159));
DFF_X1 \finalResult_reg[29]  (.Q (n_35), .CK (CTS_n_tid0_63), .D (n_0_160));
DFF_X1 \finalResult_reg[30]  (.Q (n_34), .CK (CTS_n_tid0_63), .D (n_0_161));
DFF_X1 \finalResult_reg[31]  (.Q (n_33), .CK (CTS_n_tid0_63), .D (n_0_162));
DFF_X1 \finalResult_reg[32]  (.Q (n_32), .CK (CTS_n_tid0_63), .D (n_0_163));
DFF_X1 \finalResult_reg[33]  (.Q (n_31), .CK (CTS_n_tid0_64), .D (n_0_164));
DFF_X1 \finalResult_reg[34]  (.Q (n_30), .CK (CTS_n_tid0_64), .D (n_0_165));
DFF_X1 \finalResult_reg[35]  (.Q (n_29), .CK (CTS_n_tid0_64), .D (n_0_166));
DFF_X1 \finalResult_reg[36]  (.Q (n_28), .CK (CTS_n_tid0_64), .D (n_0_167));
DFF_X1 \finalResult_reg[37]  (.Q (n_27), .CK (CTS_n_tid0_64), .D (n_0_168));
DFF_X1 \finalResult_reg[38]  (.Q (n_26), .CK (CTS_n_tid0_64), .D (n_0_169));
DFF_X1 \finalResult_reg[39]  (.Q (n_25), .CK (CTS_n_tid0_64), .D (n_0_170));
DFF_X1 \finalResult_reg[40]  (.Q (n_24), .CK (CTS_n_tid0_64), .D (n_0_171));
DFF_X1 \finalResult_reg[41]  (.Q (n_23), .CK (CTS_n_tid0_64), .D (n_0_172));
DFF_X1 \finalResult_reg[42]  (.Q (n_22), .CK (CTS_n_tid0_64), .D (n_0_173));
DFF_X1 \finalResult_reg[43]  (.Q (n_21), .CK (CTS_n_tid0_64), .D (n_0_174));
DFF_X1 \finalResult_reg[44]  (.Q (n_20), .CK (CTS_n_tid0_64), .D (n_0_175));
DFF_X1 \finalResult_reg[45]  (.Q (n_19), .CK (CTS_n_tid0_64), .D (n_0_176));
DFF_X1 \finalResult_reg[46]  (.Q (n_18), .CK (CTS_n_tid0_64), .D (n_0_177));
DFF_X1 \finalResult_reg[47]  (.Q (n_17), .CK (CTS_n_tid0_64), .D (n_0_178));
DFF_X1 \finalResult_reg[48]  (.Q (n_16), .CK (CTS_n_tid0_64), .D (n_0_179));
DFF_X1 \finalResult_reg[49]  (.Q (n_15), .CK (CTS_n_tid0_64), .D (n_0_180));
DFF_X1 \finalResult_reg[50]  (.Q (n_14), .CK (CTS_n_tid0_64), .D (n_0_181));
DFF_X1 \finalResult_reg[51]  (.Q (n_13), .CK (CTS_n_tid0_64), .D (n_0_182));
DFF_X1 \finalResult_reg[52]  (.Q (n_12), .CK (CTS_n_tid0_63), .D (n_0_183));
DFF_X1 \finalResult_reg[53]  (.Q (n_11), .CK (CTS_n_tid0_63), .D (n_0_184));
DFF_X1 \finalResult_reg[54]  (.Q (n_10), .CK (CTS_n_tid0_63), .D (n_0_185));
DFF_X1 \finalResult_reg[55]  (.Q (n_9), .CK (CTS_n_tid0_63), .D (n_0_186));
DFF_X1 \finalResult_reg[56]  (.Q (n_8), .CK (CTS_n_tid0_63), .D (n_0_187));
DFF_X1 \finalResult_reg[57]  (.Q (n_7), .CK (CTS_n_tid0_63), .D (n_0_188));
DFF_X1 \finalResult_reg[58]  (.Q (n_6), .CK (CTS_n_tid0_63), .D (n_0_189));
DFF_X1 \finalResult_reg[59]  (.Q (n_5), .CK (CTS_n_tid0_63), .D (n_0_190));
DFF_X1 \finalResult_reg[60]  (.Q (n_4), .CK (CTS_n_tid0_63), .D (n_0_191));
DFF_X1 \finalResult_reg[61]  (.Q (n_3), .CK (CTS_n_tid0_63), .D (n_0_192));
DFF_X1 \finalResult_reg[62]  (.Q (n_2), .CK (CTS_n_tid0_63), .D (n_0_193));
DFF_X1 \finalResult_reg[63]  (.Q (n_1), .CK (CTS_n_tid0_63), .D (n_0_194));
INV_X1 i_0_128 (.ZN (n_0), .A (enableRegisterOutput));
DFF_X1 enableRegisterOutput_reg (.Q (enableRegisterOutput), .CK (CTS_n_tid0_64), .D (enable));
datapath i_0_0 (.firstInputComplement ({\firstInputComplement[31] , \firstInputComplement[30] , 
    \firstInputComplement[29] , \firstInputComplement[28] , \firstInputComplement[27] , 
    \firstInputComplement[26] , \firstInputComplement[25] , \firstInputComplement[24] , 
    \firstInputComplement[23] , \firstInputComplement[22] , \firstInputComplement[21] , 
    \firstInputComplement[20] , \firstInputComplement[19] , \firstInputComplement[18] , 
    \firstInputComplement[17] , \firstInputComplement[16] , \firstInputComplement[15] , 
    \firstInputComplement[14] , \firstInputComplement[13] , \firstInputComplement[12] , 
    \firstInputComplement[11] , \firstInputComplement[10] , \firstInputComplement[9] , 
    \firstInputComplement[8] , \firstInputComplement[7] , \firstInputComplement[6] , 
    \firstInputComplement[5] , \firstInputComplement[4] , \firstInputComplement[3] , 
    \firstInputComplement[2] , \firstInputComplement[1] , uc_0}), .inputOne ({inputOne[31], 
    inputOne[30], inputOne[29], inputOne[28], inputOne[27], inputOne[26], inputOne[25], 
    inputOne[24], inputOne[23], inputOne[22], inputOne[21], inputOne[20], inputOne[19], 
    inputOne[18], inputOne[17], inputOne[16], inputOne[15], inputOne[14], inputOne[13], 
    inputOne[12], inputOne[11], inputOne[10], inputOne[9], inputOne[8], inputOne[7], 
    inputOne[6], inputOne[5], inputOne[4], inputOne[3], inputOne[2], inputOne[1], 
    inputOne[0]}));
TBUF_X1 i_127 (.Z (finalResult[63]), .A (n_1), .EN (hfn_ipo_n46));
TBUF_X1 i_125 (.Z (finalResult[62]), .A (n_2), .EN (hfn_ipo_n46));
TBUF_X1 i_123 (.Z (finalResult[61]), .A (n_3), .EN (hfn_ipo_n46));
TBUF_X1 i_121 (.Z (finalResult[60]), .A (n_4), .EN (hfn_ipo_n46));
TBUF_X1 i_119 (.Z (finalResult[59]), .A (n_5), .EN (hfn_ipo_n46));
TBUF_X1 i_117 (.Z (finalResult[58]), .A (n_6), .EN (hfn_ipo_n46));
TBUF_X1 i_115 (.Z (finalResult[57]), .A (n_7), .EN (hfn_ipo_n46));
TBUF_X1 i_113 (.Z (finalResult[56]), .A (n_8), .EN (hfn_ipo_n46));
TBUF_X1 i_111 (.Z (finalResult[55]), .A (n_9), .EN (hfn_ipo_n46));
TBUF_X1 i_109 (.Z (finalResult[54]), .A (n_10), .EN (hfn_ipo_n45));
TBUF_X1 i_107 (.Z (finalResult[53]), .A (n_11), .EN (hfn_ipo_n45));
TBUF_X1 i_105 (.Z (finalResult[52]), .A (n_12), .EN (hfn_ipo_n46));
TBUF_X1 i_103 (.Z (finalResult[51]), .A (n_13), .EN (hfn_ipo_n45));
TBUF_X1 i_101 (.Z (finalResult[50]), .A (n_14), .EN (hfn_ipo_n45));
TBUF_X1 i_99 (.Z (finalResult[49]), .A (n_15), .EN (hfn_ipo_n45));
TBUF_X1 i_97 (.Z (finalResult[48]), .A (n_16), .EN (hfn_ipo_n45));
TBUF_X1 i_95 (.Z (finalResult[47]), .A (n_17), .EN (hfn_ipo_n45));
TBUF_X1 i_93 (.Z (finalResult[46]), .A (n_18), .EN (hfn_ipo_n45));
TBUF_X1 i_91 (.Z (finalResult[45]), .A (n_19), .EN (hfn_ipo_n45));
TBUF_X1 i_89 (.Z (finalResult[44]), .A (n_20), .EN (hfn_ipo_n45));
TBUF_X1 i_87 (.Z (finalResult[43]), .A (n_21), .EN (hfn_ipo_n45));
TBUF_X1 i_85 (.Z (finalResult[42]), .A (n_22), .EN (hfn_ipo_n45));
TBUF_X1 i_83 (.Z (finalResult[41]), .A (n_23), .EN (hfn_ipo_n45));
TBUF_X1 i_81 (.Z (finalResult[40]), .A (n_24), .EN (hfn_ipo_n45));
TBUF_X1 i_79 (.Z (finalResult[39]), .A (n_25), .EN (hfn_ipo_n45));
TBUF_X1 i_77 (.Z (finalResult[38]), .A (n_26), .EN (hfn_ipo_n45));
TBUF_X1 i_75 (.Z (finalResult[37]), .A (n_27), .EN (hfn_ipo_n45));
TBUF_X1 i_73 (.Z (finalResult[36]), .A (n_28), .EN (hfn_ipo_n45));
TBUF_X1 i_71 (.Z (finalResult[35]), .A (n_29), .EN (hfn_ipo_n45));
TBUF_X1 i_69 (.Z (finalResult[34]), .A (n_30), .EN (hfn_ipo_n45));
TBUF_X1 i_67 (.Z (finalResult[33]), .A (n_31), .EN (hfn_ipo_n45));
TBUF_X1 i_65 (.Z (finalResult[32]), .A (n_32), .EN (hfn_ipo_n45));
TBUF_X1 i_63 (.Z (finalResult[31]), .A (n_33), .EN (hfn_ipo_n46));
TBUF_X1 i_61 (.Z (finalResult[30]), .A (n_34), .EN (hfn_ipo_n46));
TBUF_X1 i_59 (.Z (finalResult[29]), .A (n_35), .EN (hfn_ipo_n46));
TBUF_X1 i_57 (.Z (finalResult[28]), .A (n_36), .EN (hfn_ipo_n46));
TBUF_X1 i_55 (.Z (finalResult[27]), .A (n_37), .EN (hfn_ipo_n46));
TBUF_X1 i_53 (.Z (finalResult[26]), .A (n_38), .EN (hfn_ipo_n46));
TBUF_X1 i_51 (.Z (finalResult[25]), .A (n_39), .EN (hfn_ipo_n46));
TBUF_X1 i_49 (.Z (finalResult[24]), .A (n_40), .EN (hfn_ipo_n46));
TBUF_X1 i_47 (.Z (finalResult[23]), .A (n_41), .EN (hfn_ipo_n46));
TBUF_X1 i_45 (.Z (finalResult[22]), .A (n_42), .EN (hfn_ipo_n46));
TBUF_X1 i_43 (.Z (finalResult[21]), .A (n_43), .EN (hfn_ipo_n46));
TBUF_X1 i_41 (.Z (finalResult[20]), .A (n_44), .EN (hfn_ipo_n45));
TBUF_X1 i_39 (.Z (finalResult[19]), .A (n_45), .EN (hfn_ipo_n45));
TBUF_X1 i_37 (.Z (finalResult[18]), .A (n_46), .EN (hfn_ipo_n45));
TBUF_X1 i_35 (.Z (finalResult[17]), .A (n_47), .EN (hfn_ipo_n45));
TBUF_X1 i_33 (.Z (finalResult[16]), .A (n_48), .EN (hfn_ipo_n46));
TBUF_X1 i_31 (.Z (finalResult[15]), .A (n_49), .EN (hfn_ipo_n45));
TBUF_X1 i_29 (.Z (finalResult[14]), .A (n_50), .EN (hfn_ipo_n45));
TBUF_X1 i_27 (.Z (finalResult[13]), .A (n_51), .EN (hfn_ipo_n45));
TBUF_X1 i_25 (.Z (finalResult[12]), .A (n_52), .EN (hfn_ipo_n45));
TBUF_X1 i_23 (.Z (finalResult[11]), .A (n_53), .EN (hfn_ipo_n45));
TBUF_X1 i_21 (.Z (finalResult[10]), .A (n_54), .EN (hfn_ipo_n45));
TBUF_X1 i_19 (.Z (finalResult[9]), .A (n_55), .EN (hfn_ipo_n45));
TBUF_X1 i_17 (.Z (finalResult[8]), .A (n_56), .EN (hfn_ipo_n45));
TBUF_X1 i_15 (.Z (finalResult[7]), .A (n_57), .EN (hfn_ipo_n45));
TBUF_X1 i_13 (.Z (finalResult[6]), .A (n_58), .EN (hfn_ipo_n45));
TBUF_X1 i_11 (.Z (finalResult[5]), .A (n_59), .EN (hfn_ipo_n45));
TBUF_X1 i_9 (.Z (finalResult[4]), .A (n_60), .EN (hfn_ipo_n45));
TBUF_X1 i_7 (.Z (finalResult[3]), .A (n_61), .EN (hfn_ipo_n45));
TBUF_X1 i_5 (.Z (finalResult[2]), .A (n_62), .EN (hfn_ipo_n45));
TBUF_X1 i_3 (.Z (finalResult[1]), .A (n_63), .EN (hfn_ipo_n45));
TBUF_X1 i_1 (.Z (finalResult[0]), .A (n_64), .EN (hfn_ipo_n45));
CLKBUF_X2 hfn_ipo_c35 (.Z (hfn_ipo_n35), .A (n_0_1_12));
CLKBUF_X2 hfn_ipo_c36 (.Z (hfn_ipo_n36), .A (n_0_1_12));
BUF_X4 drc_ipo_c47 (.Z (drc_ipo_n47), .A (\counter[2] ));
CLKBUF_X3 drc_ipo_c48 (.Z (drc_ipo_n48), .A (n_0_1_62));
BUF_X4 hfn_ipo_c37 (.Z (hfn_ipo_n37), .A (n_0_1_13));
CLKBUF_X2 CTS_L3_c_tid0_65 (.Z (CTS_n_tid0_63), .A (clk_CTS_0_PP_10));
CLKBUF_X2 hfn_ipo_c42 (.Z (hfn_ipo_n42), .A (\counter[1] ));
CLKBUF_X3 hfn_ipo_c43 (.Z (hfn_ipo_n43), .A (\counter[0] ));
CLKBUF_X1 hfn_ipo_c41 (.Z (hfn_ipo_n41), .A (\counter[1] ));
BUF_X4 hfn_ipo_c44 (.Z (hfn_ipo_n44), .A (\counter[0] ));
BUF_X4 hfn_ipo_c45 (.Z (hfn_ipo_n45), .A (n_0));
CLKBUF_X1 hfn_ipo_c46 (.Z (hfn_ipo_n46), .A (n_0));
BUF_X4 hfn_ipo_c33 (.Z (hfn_ipo_n33), .A (n_0_1_6));
CLKBUF_X1 hfn_ipo_c34 (.Z (hfn_ipo_n34), .A (n_0_1_6));
CLKBUF_X1 hfn_ipo_c40 (.Z (hfn_ipo_n40), .A (n_0_1_15));
CLKBUF_X2 CTS_L2_c_tid0_66 (.Z (CTS_n_tid0_64), .A (clk_CTS_0_PP_11));

endmodule //RadixNoaman

module finalRadix4 (inputA, inputB, clk, reset, en, result);

output [63:0] result;
input clk;
input en;
input [31:0] inputA;
input [31:0] inputB;
input reset;
wire CLOCK_slh_n174;
wire CLOCK_slh_n249;
wire CLOCK_slh_n144;
wire CLOCK_slh_n124;
wire CLOCK_slh_n219;
wire CLOCK_slh_n244;
wire CLOCK_slh_n209;
wire CLOCK_slh_n214;
wire CLOCK_slh_n149;
wire CLOCK_slh_n89;
wire CLOCK_slh_n114;
wire CLOCK_slh_n94;
wire CLOCK_slh_n169;
wire CLOCK_slh_n189;
wire CLOCK_slh_n154;
wire CLOCK_slh_n119;
wire CLOCK_slh_n129;
wire CLOCK_slh_n104;
wire CLOCK_slh_n99;
wire CLOCK_slh_n164;
wire CLOCK_slh_n179;
wire CLOCK_slh_n139;
wire CLOCK_slh_n134;
wire CLOCK_slh_n84;
wire CLOCK_slh_n194;
wire CLOCK_slh_n159;
wire CLOCK_slh_n109;
wire CLOCK_slh_n204;
wire CLOCK_slh_n264;
wire CLOCK_slh_n199;
wire CLOCK_slh_n234;
wire CLOCK_slh_n229;
wire CLOCK_slh_n259;
wire CLOCK_slh_n184;
wire CLOCK_slh_n254;
wire CLOCK_slh_n274;
wire CLOCK_slh_n224;
wire CLOCK_slh_n239;
wire CLOCK_slh_n269;
wire enableOutput;
wire \result_out[63] ;
wire \result_out[62] ;
wire \result_out[61] ;
wire \result_out[60] ;
wire \result_out[59] ;
wire \result_out[58] ;
wire \result_out[57] ;
wire \result_out[56] ;
wire \result_out[55] ;
wire \result_out[54] ;
wire \result_out[53] ;
wire \result_out[52] ;
wire \result_out[51] ;
wire \result_out[50] ;
wire \result_out[49] ;
wire \result_out[48] ;
wire \result_out[47] ;
wire \result_out[46] ;
wire \result_out[45] ;
wire \result_out[44] ;
wire \result_out[43] ;
wire \result_out[42] ;
wire \result_out[41] ;
wire \result_out[40] ;
wire \result_out[39] ;
wire \result_out[38] ;
wire \result_out[37] ;
wire \result_out[36] ;
wire \result_out[35] ;
wire \result_out[34] ;
wire \result_out[33] ;
wire \result_out[32] ;
wire \result_out[31] ;
wire \result_out[30] ;
wire \result_out[29] ;
wire \result_out[28] ;
wire \result_out[27] ;
wire \result_out[26] ;
wire \result_out[25] ;
wire \result_out[24] ;
wire \result_out[23] ;
wire \result_out[22] ;
wire \result_out[21] ;
wire \result_out[20] ;
wire \result_out[19] ;
wire \result_out[18] ;
wire \result_out[17] ;
wire \result_out[16] ;
wire \result_out[15] ;
wire \result_out[14] ;
wire \result_out[13] ;
wire \result_out[12] ;
wire \result_out[11] ;
wire \result_out[10] ;
wire \result_out[9] ;
wire \result_out[8] ;
wire \result_out[7] ;
wire \result_out[6] ;
wire \result_out[5] ;
wire \result_out[4] ;
wire \result_out[3] ;
wire \result_out[2] ;
wire \result_out[1] ;
wire \result_out[0] ;
wire \A_reg[31] ;
wire \A_reg[30] ;
wire \A_reg[29] ;
wire \A_reg[28] ;
wire \A_reg[27] ;
wire \A_reg[26] ;
wire \A_reg[25] ;
wire \A_reg[24] ;
wire \A_reg[23] ;
wire \A_reg[22] ;
wire \A_reg[21] ;
wire \A_reg[20] ;
wire \A_reg[19] ;
wire \A_reg[18] ;
wire \A_reg[17] ;
wire \A_reg[16] ;
wire \A_reg[15] ;
wire \A_reg[14] ;
wire \A_reg[13] ;
wire \A_reg[12] ;
wire \A_reg[11] ;
wire \A_reg[10] ;
wire \A_reg[9] ;
wire \A_reg[8] ;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire \B_reg[31] ;
wire \B_reg[30] ;
wire \B_reg[29] ;
wire \B_reg[28] ;
wire \B_reg[27] ;
wire \B_reg[26] ;
wire \B_reg[25] ;
wire \B_reg[24] ;
wire \B_reg[23] ;
wire \B_reg[22] ;
wire \B_reg[21] ;
wire \B_reg[20] ;
wire \B_reg[19] ;
wire \B_reg[18] ;
wire \B_reg[17] ;
wire \B_reg[16] ;
wire \B_reg[15] ;
wire \B_reg[14] ;
wire \B_reg[13] ;
wire \B_reg[12] ;
wire \B_reg[11] ;
wire \B_reg[10] ;
wire \B_reg[9] ;
wire \B_reg[8] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;
wire drc_ipo_n1;
wire drc_ipo_n2;
wire CTS_n_tid0_72;
wire CTS_n_tid0_73;


buffer__parameterized0 out (.Q ({result[63], result[62], result[61], result[60], 
    result[59], result[58], result[57], result[56], result[55], result[54], result[53], 
    result[52], result[51], result[50], result[49], result[48], result[47], result[46], 
    result[45], result[44], result[43], result[42], result[41], result[40], result[39], 
    result[38], result[37], result[36], result[35], result[34], result[33], result[32], 
    result[31], result[30], result[29], result[28], result[27], result[26], result[25], 
    result[24], result[23], result[22], result[21], result[20], result[19], result[18], 
    result[17], result[16], result[15], result[14], result[13], result[12], result[11], 
    result[10], result[9], result[8], result[7], result[6], result[5], result[4], 
    result[3], result[2], result[1], result[0]}), .D ({\result_out[63] , \result_out[62] , 
    \result_out[61] , \result_out[60] , \result_out[59] , \result_out[58] , \result_out[57] , 
    \result_out[56] , \result_out[55] , \result_out[54] , \result_out[53] , \result_out[52] , 
    \result_out[51] , \result_out[50] , \result_out[49] , \result_out[48] , \result_out[47] , 
    \result_out[46] , \result_out[45] , \result_out[44] , \result_out[43] , \result_out[42] , 
    \result_out[41] , \result_out[40] , \result_out[39] , \result_out[38] , \result_out[37] , 
    \result_out[36] , \result_out[35] , \result_out[34] , \result_out[33] , \result_out[32] , 
    \result_out[31] , \result_out[30] , \result_out[29] , \result_out[28] , \result_out[27] , 
    \result_out[26] , \result_out[25] , \result_out[24] , \result_out[23] , \result_out[22] , 
    \result_out[21] , \result_out[20] , \result_out[19] , \result_out[18] , \result_out[17] , 
    \result_out[16] , \result_out[15] , \result_out[14] , \result_out[13] , \result_out[12] , 
    \result_out[11] , \result_out[10] , \result_out[9] , \result_out[8] , \result_out[7] , 
    \result_out[6] , \result_out[5] , \result_out[4] , \result_out[3] , \result_out[2] , 
    \result_out[1] , \result_out[0] }), .en (enableOutput), .rst (drc_ipo_n2), .clk_CTS_0_PP_10 (CTS_n_tid0_73));
buffer regB (.Q ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , \B_reg[27] , 
    \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , \B_reg[21] , 
    \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , \B_reg[15] , 
    \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , \B_reg[9] , 
    \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , \B_reg[2] , 
    \B_reg[1] , \B_reg[0] }), .D ({CLOCK_slh_n204, inputB[30], inputB[29], inputB[28], 
    CLOCK_slh_n264, CLOCK_slh_n199, inputB[25], inputB[24], inputB[23], inputB[22], 
    inputB[21], CLOCK_slh_n234, inputB[19], CLOCK_slh_n229, inputB[17], CLOCK_slh_n259, 
    CLOCK_slh_n184, inputB[14], inputB[13], CLOCK_slh_n254, CLOCK_slh_n274, inputB[10], 
    inputB[9], inputB[8], CLOCK_slh_n224, inputB[6], inputB[5], CLOCK_slh_n239, CLOCK_slh_n269, 
    inputB[2], inputB[1], inputB[0]}), .en (drc_ipo_n1), .rst (drc_ipo_n2), .clk_CTS_0_PP_11 (CTS_n_tid0_73));
buffer__0_18 regA (.Q ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , \A_reg[27] , 
    \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , \A_reg[21] , 
    \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , \A_reg[15] , 
    \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , \A_reg[9] , 
    \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , \A_reg[2] , 
    \A_reg[1] , \A_reg[0] }), .D ({inputA[31], CLOCK_slh_n174, inputA[29], inputA[28], 
    inputA[27], CLOCK_slh_n249, CLOCK_slh_n144, CLOCK_slh_n124, CLOCK_slh_n219, CLOCK_slh_n244, 
    CLOCK_slh_n209, CLOCK_slh_n214, CLOCK_slh_n149, CLOCK_slh_n89, CLOCK_slh_n114, 
    CLOCK_slh_n94, CLOCK_slh_n169, CLOCK_slh_n189, inputA[13], CLOCK_slh_n154, CLOCK_slh_n119, 
    CLOCK_slh_n129, CLOCK_slh_n104, CLOCK_slh_n99, CLOCK_slh_n164, CLOCK_slh_n179, 
    CLOCK_slh_n139, CLOCK_slh_n134, CLOCK_slh_n84, CLOCK_slh_n194, CLOCK_slh_n159, 
    CLOCK_slh_n109}), .en (drc_ipo_n1), .rst (drc_ipo_n2), .clk_CTS_0_PP_10 (CTS_n_tid0_73));
RadixNoaman radixNoamanMult (.enableRegisterOutput (enableOutput), .finalResult ({
    \result_out[63] , \result_out[62] , \result_out[61] , \result_out[60] , \result_out[59] , 
    \result_out[58] , \result_out[57] , \result_out[56] , \result_out[55] , \result_out[54] , 
    \result_out[53] , \result_out[52] , \result_out[51] , \result_out[50] , \result_out[49] , 
    \result_out[48] , \result_out[47] , \result_out[46] , \result_out[45] , \result_out[44] , 
    \result_out[43] , \result_out[42] , \result_out[41] , \result_out[40] , \result_out[39] , 
    \result_out[38] , \result_out[37] , \result_out[36] , \result_out[35] , \result_out[34] , 
    \result_out[33] , \result_out[32] , \result_out[31] , \result_out[30] , \result_out[29] , 
    \result_out[28] , \result_out[27] , \result_out[26] , \result_out[25] , \result_out[24] , 
    \result_out[23] , \result_out[22] , \result_out[21] , \result_out[20] , \result_out[19] , 
    \result_out[18] , \result_out[17] , \result_out[16] , \result_out[15] , \result_out[14] , 
    \result_out[13] , \result_out[12] , \result_out[11] , \result_out[10] , \result_out[9] , 
    \result_out[8] , \result_out[7] , \result_out[6] , \result_out[5] , \result_out[4] , 
    \result_out[3] , \result_out[2] , \result_out[1] , \result_out[0] }), .enable (drc_ipo_n1)
    , .inputOne ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , \A_reg[27] , 
    \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , \A_reg[21] , 
    \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , \A_reg[15] , 
    \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , \A_reg[9] , 
    \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , \A_reg[2] , 
    \A_reg[1] , \A_reg[0] }), .inputTwo ({\B_reg[31] , \B_reg[30] , \B_reg[29] , 
    \B_reg[28] , \B_reg[27] , \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , 
    \B_reg[22] , \B_reg[21] , \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , 
    \B_reg[16] , \B_reg[15] , \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , 
    \B_reg[10] , \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , 
    \B_reg[3] , \B_reg[2] , \B_reg[1] , \B_reg[0] }), .reset (drc_ipo_n2), .clk_CTS_0_PP_10 (CTS_n_tid0_72)
    , .clk_CTS_0_PP_11 (CTS_n_tid0_73));
CLKBUF_X1 drc_ipo_c1 (.Z (drc_ipo_n1), .A (en));
CLKBUF_X1 drc_ipo_c2 (.Z (drc_ipo_n2), .A (reset));
CLKBUF_X2 CTS_L1_tid0__c1_tid0__c3 (.Z (CTS_n_tid0_73), .A (clk));
CLKBUF_X1 CLOCK_slh__c33 (.Z (CLOCK_slh_n84), .A (inputA[3]));
CLKBUF_X1 CLOCK_slh__c35 (.Z (CLOCK_slh_n89), .A (inputA[18]));
CLKBUF_X1 CLOCK_slh__c37 (.Z (CLOCK_slh_n94), .A (inputA[16]));
CLKBUF_X1 CLOCK_slh__c39 (.Z (CLOCK_slh_n99), .A (inputA[8]));
CLKBUF_X1 CTS_L2_c_tid0_32 (.Z (CTS_n_tid0_72), .A (CTS_n_tid0_73));
CLKBUF_X1 CLOCK_slh__c41 (.Z (CLOCK_slh_n104), .A (inputA[9]));
CLKBUF_X1 CLOCK_slh__c43 (.Z (CLOCK_slh_n109), .A (inputA[0]));
CLKBUF_X1 CLOCK_slh__c45 (.Z (CLOCK_slh_n114), .A (inputA[17]));
CLKBUF_X1 CLOCK_slh__c47 (.Z (CLOCK_slh_n119), .A (inputA[11]));
CLKBUF_X1 CLOCK_slh__c49 (.Z (CLOCK_slh_n124), .A (inputA[24]));
CLKBUF_X1 CLOCK_slh__c51 (.Z (CLOCK_slh_n129), .A (inputA[10]));
CLKBUF_X1 CLOCK_slh__c53 (.Z (CLOCK_slh_n134), .A (inputA[4]));
CLKBUF_X1 CLOCK_slh__c55 (.Z (CLOCK_slh_n139), .A (inputA[5]));
CLKBUF_X1 CLOCK_slh__c57 (.Z (CLOCK_slh_n144), .A (inputA[25]));
CLKBUF_X1 CLOCK_slh__c59 (.Z (CLOCK_slh_n149), .A (inputA[19]));
CLKBUF_X1 CLOCK_slh__c61 (.Z (CLOCK_slh_n154), .A (inputA[12]));
CLKBUF_X1 CLOCK_slh__c63 (.Z (CLOCK_slh_n159), .A (inputA[1]));
CLKBUF_X1 CLOCK_slh__c65 (.Z (CLOCK_slh_n164), .A (inputA[7]));
CLKBUF_X1 CLOCK_slh__c67 (.Z (CLOCK_slh_n169), .A (inputA[15]));
CLKBUF_X1 CLOCK_slh__c69 (.Z (CLOCK_slh_n174), .A (inputA[30]));
CLKBUF_X1 CLOCK_slh__c71 (.Z (CLOCK_slh_n179), .A (inputA[6]));
CLKBUF_X1 CLOCK_slh__c73 (.Z (CLOCK_slh_n184), .A (inputB[15]));
CLKBUF_X1 CLOCK_slh__c75 (.Z (CLOCK_slh_n189), .A (inputA[14]));
CLKBUF_X1 CLOCK_slh__c77 (.Z (CLOCK_slh_n194), .A (inputA[2]));
CLKBUF_X1 CLOCK_slh__c79 (.Z (CLOCK_slh_n199), .A (inputB[26]));
CLKBUF_X1 CLOCK_slh__c81 (.Z (CLOCK_slh_n204), .A (inputB[31]));
CLKBUF_X1 CLOCK_slh__c83 (.Z (CLOCK_slh_n209), .A (inputA[21]));
CLKBUF_X1 CLOCK_slh__c85 (.Z (CLOCK_slh_n214), .A (inputA[20]));
CLKBUF_X1 CLOCK_slh__c87 (.Z (CLOCK_slh_n219), .A (inputA[23]));
CLKBUF_X1 CLOCK_slh__c89 (.Z (CLOCK_slh_n224), .A (inputB[7]));
CLKBUF_X1 CLOCK_slh__c91 (.Z (CLOCK_slh_n229), .A (inputB[18]));
CLKBUF_X1 CLOCK_slh__c93 (.Z (CLOCK_slh_n234), .A (inputB[20]));
CLKBUF_X1 CLOCK_slh__c95 (.Z (CLOCK_slh_n239), .A (inputB[4]));
CLKBUF_X1 CLOCK_slh__c97 (.Z (CLOCK_slh_n244), .A (inputA[22]));
CLKBUF_X1 CLOCK_slh__c99 (.Z (CLOCK_slh_n249), .A (inputA[26]));
CLKBUF_X1 CLOCK_slh__c101 (.Z (CLOCK_slh_n254), .A (inputB[12]));
CLKBUF_X1 CLOCK_slh__c103 (.Z (CLOCK_slh_n259), .A (inputB[16]));
CLKBUF_X1 CLOCK_slh__c105 (.Z (CLOCK_slh_n264), .A (inputB[27]));
CLKBUF_X1 CLOCK_slh__c107 (.Z (CLOCK_slh_n269), .A (inputB[3]));
CLKBUF_X1 CLOCK_slh__c109 (.Z (CLOCK_slh_n274), .A (inputB[11]));

endmodule //finalRadix4


