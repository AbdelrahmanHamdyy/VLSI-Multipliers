/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Jan  4 05:56:05 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 808492695 */

module datapath__0_0(p_0, p_1);
   output [32:0]p_0;
   input [32:0]p_1;

   XOR2_X1 i_0 (.A(p_1[2]), .B(p_1[1]), .Z(p_0[2]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[3]));
   OAI21_X1 i_2 (.A(p_1[3]), .B1(p_1[2]), .B2(p_1[1]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_1[4]), .B(n_29), .Z(p_0[4]));
   XOR2_X1 i_4 (.A(p_1[5]), .B(n_28), .Z(p_0[5]));
   XOR2_X1 i_5 (.A(p_1[6]), .B(n_27), .Z(p_0[6]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[7]));
   OAI21_X1 i_7 (.A(p_1[7]), .B1(n_27), .B2(p_1[6]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_1[8]), .B(n_26), .Z(p_0[8]));
   XOR2_X1 i_9 (.A(p_1[9]), .B(n_25), .Z(p_0[9]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[10]));
   OAI21_X1 i_11 (.A(p_1[10]), .B1(n_25), .B2(p_1[9]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_1[11]), .B(n_24), .Z(p_0[11]));
   XNOR2_X1 i_13 (.A(p_1[12]), .B(n_23), .ZN(p_0[12]));
   XOR2_X1 i_14 (.A(p_1[13]), .B(n_22), .Z(p_0[13]));
   XNOR2_X1 i_15 (.A(p_1[14]), .B(n_21), .ZN(p_0[14]));
   XNOR2_X1 i_16 (.A(p_1[15]), .B(n_20), .ZN(p_0[15]));
   XOR2_X1 i_17 (.A(p_1[16]), .B(n_19), .Z(p_0[16]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[17]));
   OAI21_X1 i_19 (.A(p_1[17]), .B1(n_19), .B2(p_1[16]), .ZN(n_3));
   XOR2_X1 i_20 (.A(p_1[18]), .B(n_18), .Z(p_0[18]));
   XOR2_X1 i_21 (.A(p_1[19]), .B(n_17), .Z(p_0[19]));
   XNOR2_X1 i_22 (.A(p_1[20]), .B(n_16), .ZN(p_0[20]));
   XNOR2_X1 i_23 (.A(p_1[21]), .B(n_15), .ZN(p_0[21]));
   XNOR2_X1 i_24 (.A(p_1[22]), .B(n_14), .ZN(p_0[22]));
   XOR2_X1 i_25 (.A(p_1[23]), .B(n_13), .Z(p_0[23]));
   XOR2_X1 i_26 (.A(p_1[24]), .B(n_12), .Z(p_0[24]));
   XNOR2_X1 i_27 (.A(p_1[25]), .B(n_11), .ZN(p_0[25]));
   XNOR2_X1 i_28 (.A(p_1[26]), .B(n_10), .ZN(p_0[26]));
   XOR2_X1 i_29 (.A(p_1[27]), .B(n_9), .Z(p_0[27]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[28]));
   OAI21_X1 i_31 (.A(p_1[28]), .B1(n_9), .B2(p_1[27]), .ZN(n_4));
   XOR2_X1 i_32 (.A(p_1[29]), .B(n_8), .Z(p_0[29]));
   XNOR2_X1 i_33 (.A(p_1[30]), .B(n_7), .ZN(p_0[30]));
   XNOR2_X1 i_34 (.A(p_1[31]), .B(n_6), .ZN(p_0[31]));
   XNOR2_X1 i_35 (.A(p_1[32]), .B(n_5), .ZN(p_0[32]));
   NOR4_X1 i_36 (.A1(n_8), .A2(p_1[29]), .A3(p_1[30]), .A4(p_1[31]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(p_1[29]), .A3(p_1[30]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(p_1[29]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(p_1[27]), .A3(p_1[28]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(p_1[24]), .A3(p_1[25]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(p_1[24]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(p_1[23]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(p_1[19]), .A3(p_1[20]), .A4(p_1[21]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(p_1[19]), .A3(p_1[20]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(p_1[19]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(p_1[18]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(p_1[16]), .A3(p_1[17]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(p_1[13]), .A3(p_1[14]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(p_1[13]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(p_1[11]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(p_1[9]), .A3(p_1[10]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(p_1[8]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(p_1[6]), .A3(p_1[7]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(p_1[5]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(p_1[4]), .ZN(n_28));
   OR3_X1 i_60 (.A1(p_1[3]), .A2(p_1[2]), .A3(p_1[1]), .ZN(n_29));
   INV_X1 i_61 (.A(p_1[12]), .ZN(n_30));
   INV_X1 i_62 (.A(p_1[15]), .ZN(n_31));
   INV_X1 i_63 (.A(p_1[22]), .ZN(n_32));
   INV_X1 i_64 (.A(p_1[26]), .ZN(n_33));
endmodule

module datapath__0_12(p_0, tempResult, p_1);
   input [63:0]p_0;
   input [63:0]tempResult;
   output [63:0]p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1[0]));
   OAI21_X1 i_1 (.A(n_366), .B1(p_0[0]), .B2(tempResult[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_366), .B(n_1), .Z(p_1[1]));
   OAI21_X1 i_3 (.A(n_365), .B1(p_0[1]), .B2(tempResult[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_364), .B(n_2), .ZN(p_1[2]));
   OAI21_X1 i_5 (.A(n_369), .B1(p_0[2]), .B2(tempResult[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_363), .B(n_3), .Z(p_1[3]));
   OAI21_X1 i_7 (.A(n_370), .B1(n_376), .B2(n_372), .ZN(n_3));
   XOR2_X1 i_8 (.A(n_361), .B(n_10), .Z(p_1[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_1[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_1[6]));
   NOR2_X1 i_11 (.A1(n_358), .A2(n_349), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_1[7]));
   OAI22_X1 i_13 (.A1(p_0[6]), .A2(tempResult[6]), .B1(n_349), .B2(n_7), 
      .ZN(n_5));
   AOI21_X1 i_14 (.A(n_359), .B1(p_0[5]), .B2(tempResult[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_359), .B1(n_353), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_356), .B1(n_361), .B2(n_354), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_354), .B1(p_0[4]), .B2(tempResult[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_360), .A2(n_351), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_347), .B(n_18), .ZN(p_1[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_1[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_1[10]));
   NOR2_X1 i_23 (.A1(n_344), .A2(n_335), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_1[11]));
   OAI22_X1 i_25 (.A1(p_0[10]), .A2(tempResult[10]), .B1(n_335), .B2(n_15), 
      .ZN(n_13));
   AOI21_X1 i_26 (.A(n_345), .B1(p_0[9]), .B2(tempResult[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_345), .B1(n_339), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_342), .B1(n_347), .B2(n_340), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_342), .B1(p_0[8]), .B2(tempResult[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_346), .A2(n_337), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_333), .B(n_26), .Z(p_1[12]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(p_1[13]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(p_1[14]));
   NOR2_X1 i_35 (.A1(n_330), .A2(n_321), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(p_1[15]));
   OAI22_X1 i_37 (.A1(p_0[14]), .A2(tempResult[14]), .B1(n_321), .B2(n_23), 
      .ZN(n_21));
   AOI21_X1 i_38 (.A(n_331), .B1(p_0[13]), .B2(tempResult[13]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_331), .B1(n_325), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_328), .B1(n_333), .B2(n_326), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_326), .B1(p_0[12]), .B2(tempResult[12]), .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_332), .A2(n_323), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_319), .B(n_34), .Z(p_1[16]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(p_1[17]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(p_1[18]));
   NOR2_X1 i_47 (.A1(n_285), .A2(n_275), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(p_1[19]));
   OAI21_X1 i_49 (.A(n_284), .B1(n_275), .B2(n_31), .ZN(n_29));
   NOR2_X1 i_50 (.A1(n_287), .A2(n_277), .ZN(n_30));
   INV_X1 i_51 (.A(n_32), .ZN(n_31));
   OAI21_X1 i_52 (.A(n_286), .B1(n_277), .B2(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_282), .B1(n_319), .B2(n_279), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_279), .B1(p_0[16]), .B2(tempResult[16]), .ZN(n_34));
   AOI21_X1 i_55 (.A(n_289), .B1(p_0[19]), .B2(tempResult[19]), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_63), .B(n_42), .Z(p_1[20]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(p_1[21]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(p_1[22]));
   NOR2_X1 i_59 (.A1(n_313), .A2(n_257), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(p_1[23]));
   OAI21_X1 i_61 (.A(n_312), .B1(n_257), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_315), .A2(n_259), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_314), .B1(n_259), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_318), .B1(n_261), .B2(n_63), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_261), .B1(p_0[20]), .B2(tempResult[20]), .ZN(n_42));
   AOI21_X1 i_67 (.A(n_317), .B1(p_0[23]), .B2(tempResult[23]), .ZN(n_43));
   XOR2_X1 i_68 (.A(n_61), .B(n_50), .Z(p_1[24]));
   XOR2_X1 i_69 (.A(n_49), .B(n_46), .Z(p_1[25]));
   XOR2_X1 i_70 (.A(n_47), .B(n_44), .Z(p_1[26]));
   NOR2_X1 i_71 (.A1(n_296), .A2(n_269), .ZN(n_44));
   XNOR2_X1 i_72 (.A(n_51), .B(n_45), .ZN(p_1[27]));
   OAI21_X1 i_73 (.A(n_295), .B1(n_269), .B2(n_47), .ZN(n_45));
   NOR2_X1 i_74 (.A1(n_298), .A2(n_271), .ZN(n_46));
   INV_X1 i_75 (.A(n_48), .ZN(n_47));
   OAI21_X1 i_76 (.A(n_297), .B1(n_271), .B2(n_49), .ZN(n_48));
   AOI21_X1 i_77 (.A(n_293), .B1(n_273), .B2(n_61), .ZN(n_49));
   OAI21_X1 i_78 (.A(n_273), .B1(p_0[24]), .B2(tempResult[24]), .ZN(n_50));
   AOI21_X1 i_79 (.A(n_300), .B1(p_0[27]), .B2(tempResult[27]), .ZN(n_51));
   XOR2_X1 i_80 (.A(n_59), .B(n_58), .Z(p_1[28]));
   XOR2_X1 i_81 (.A(n_57), .B(n_54), .Z(p_1[29]));
   XOR2_X1 i_82 (.A(n_55), .B(n_52), .Z(p_1[30]));
   NOR2_X1 i_83 (.A1(n_305), .A2(n_263), .ZN(n_52));
   XOR2_X1 i_84 (.A(n_65), .B(n_53), .Z(p_1[31]));
   OAI21_X1 i_85 (.A(n_304), .B1(n_263), .B2(n_55), .ZN(n_53));
   NOR2_X1 i_86 (.A1(n_307), .A2(n_266), .ZN(n_54));
   INV_X1 i_87 (.A(n_56), .ZN(n_55));
   OAI21_X1 i_88 (.A(n_306), .B1(n_266), .B2(n_57), .ZN(n_56));
   AOI21_X1 i_89 (.A(n_302), .B1(n_267), .B2(n_59), .ZN(n_57));
   OAI21_X1 i_90 (.A(n_267), .B1(p_0[28]), .B2(tempResult[28]), .ZN(n_58));
   INV_X1 i_91 (.A(n_60), .ZN(n_59));
   OAI21_X1 i_92 (.A(n_268), .B1(n_292), .B2(n_61), .ZN(n_60));
   INV_X1 i_93 (.A(n_62), .ZN(n_61));
   OAI21_X1 i_94 (.A(n_256), .B1(n_310), .B2(n_63), .ZN(n_62));
   INV_X1 i_95 (.A(n_64), .ZN(n_63));
   OAI21_X1 i_96 (.A(n_274), .B1(n_319), .B2(n_281), .ZN(n_64));
   OAI21_X1 i_97 (.A(n_308), .B1(n_377), .B2(n_373), .ZN(n_65));
   XOR2_X1 i_98 (.A(n_254), .B(n_72), .Z(p_1[32]));
   XOR2_X1 i_99 (.A(n_71), .B(n_68), .Z(p_1[33]));
   XOR2_X1 i_100 (.A(n_69), .B(n_66), .Z(p_1[34]));
   NOR2_X1 i_101 (.A1(n_223), .A2(n_213), .ZN(n_66));
   XNOR2_X1 i_102 (.A(n_73), .B(n_67), .ZN(p_1[35]));
   OAI21_X1 i_103 (.A(n_222), .B1(n_213), .B2(n_69), .ZN(n_67));
   NOR2_X1 i_104 (.A1(n_225), .A2(n_215), .ZN(n_68));
   INV_X1 i_105 (.A(n_70), .ZN(n_69));
   OAI21_X1 i_106 (.A(n_224), .B1(n_215), .B2(n_71), .ZN(n_70));
   AOI21_X1 i_107 (.A(n_220), .B1(n_254), .B2(n_217), .ZN(n_71));
   OAI21_X1 i_108 (.A(n_217), .B1(p_0[32]), .B2(tempResult[32]), .ZN(n_72));
   AOI21_X1 i_109 (.A(n_227), .B1(p_0[35]), .B2(tempResult[35]), .ZN(n_73));
   XOR2_X1 i_110 (.A(n_101), .B(n_80), .Z(p_1[36]));
   XOR2_X1 i_111 (.A(n_79), .B(n_76), .Z(p_1[37]));
   XOR2_X1 i_112 (.A(n_77), .B(n_74), .Z(p_1[38]));
   NOR2_X1 i_113 (.A1(n_248), .A2(n_206), .ZN(n_74));
   XNOR2_X1 i_114 (.A(n_81), .B(n_75), .ZN(p_1[39]));
   OAI21_X1 i_115 (.A(n_247), .B1(n_206), .B2(n_77), .ZN(n_75));
   NOR2_X1 i_116 (.A1(n_250), .A2(n_208), .ZN(n_76));
   INV_X1 i_117 (.A(n_78), .ZN(n_77));
   OAI21_X1 i_118 (.A(n_249), .B1(n_208), .B2(n_79), .ZN(n_78));
   AOI21_X1 i_119 (.A(n_253), .B1(n_210), .B2(n_101), .ZN(n_79));
   OAI21_X1 i_120 (.A(n_210), .B1(p_0[36]), .B2(tempResult[36]), .ZN(n_80));
   AOI21_X1 i_121 (.A(n_252), .B1(p_0[39]), .B2(tempResult[39]), .ZN(n_81));
   XOR2_X1 i_122 (.A(n_99), .B(n_88), .Z(p_1[40]));
   XOR2_X1 i_123 (.A(n_87), .B(n_84), .Z(p_1[41]));
   XOR2_X1 i_124 (.A(n_85), .B(n_82), .Z(p_1[42]));
   NOR2_X1 i_125 (.A1(n_234), .A2(n_192), .ZN(n_82));
   XNOR2_X1 i_126 (.A(n_89), .B(n_83), .ZN(p_1[43]));
   OAI21_X1 i_127 (.A(n_233), .B1(n_192), .B2(n_85), .ZN(n_83));
   NOR2_X1 i_128 (.A1(n_236), .A2(n_194), .ZN(n_84));
   INV_X1 i_129 (.A(n_86), .ZN(n_85));
   OAI21_X1 i_130 (.A(n_235), .B1(n_194), .B2(n_87), .ZN(n_86));
   AOI21_X1 i_131 (.A(n_231), .B1(n_196), .B2(n_99), .ZN(n_87));
   OAI21_X1 i_132 (.A(n_196), .B1(p_0[40]), .B2(tempResult[40]), .ZN(n_88));
   AOI21_X1 i_133 (.A(n_238), .B1(p_0[43]), .B2(tempResult[43]), .ZN(n_89));
   XNOR2_X1 i_134 (.A(n_98), .B(n_97), .ZN(p_1[44]));
   XOR2_X1 i_135 (.A(n_95), .B(n_94), .Z(p_1[45]));
   XNOR2_X1 i_136 (.A(n_91), .B(n_90), .ZN(p_1[46]));
   OAI22_X1 i_137 (.A1(p_0[45]), .A2(tempResult[45]), .B1(n_202), .B2(n_95), 
      .ZN(n_90));
   NOR2_X1 i_138 (.A1(n_242), .A2(n_199), .ZN(n_91));
   XNOR2_X1 i_139 (.A(n_103), .B(n_92), .ZN(p_1[47]));
   OAI21_X1 i_140 (.A(n_93), .B1(n_241), .B2(n_199), .ZN(n_92));
   NAND3_X1 i_141 (.A1(n_200), .A2(n_94), .A3(n_96), .ZN(n_93));
   NOR2_X1 i_142 (.A1(n_243), .A2(n_202), .ZN(n_94));
   INV_X1 i_143 (.A(n_96), .ZN(n_95));
   OAI22_X1 i_144 (.A1(p_0[44]), .A2(tempResult[44]), .B1(n_203), .B2(n_98), 
      .ZN(n_96));
   OAI21_X1 i_145 (.A(n_204), .B1(p_0[44]), .B2(tempResult[44]), .ZN(n_97));
   OAI21_X1 i_146 (.A(n_191), .B1(n_230), .B2(n_99), .ZN(n_98));
   INV_X1 i_147 (.A(n_100), .ZN(n_99));
   OAI21_X1 i_148 (.A(n_205), .B1(n_245), .B2(n_101), .ZN(n_100));
   INV_X1 i_149 (.A(n_102), .ZN(n_101));
   OAI21_X1 i_150 (.A(n_212), .B1(n_254), .B2(n_219), .ZN(n_102));
   AOI21_X1 i_151 (.A(n_244), .B1(p_0[47]), .B2(tempResult[47]), .ZN(n_103));
   XOR2_X1 i_152 (.A(n_189), .B(n_110), .Z(p_1[48]));
   XOR2_X1 i_153 (.A(n_109), .B(n_106), .Z(p_1[49]));
   XOR2_X1 i_154 (.A(n_107), .B(n_104), .Z(p_1[50]));
   NOR2_X1 i_155 (.A1(n_186), .A2(n_177), .ZN(n_104));
   XNOR2_X1 i_156 (.A(n_111), .B(n_105), .ZN(p_1[51]));
   OAI22_X1 i_157 (.A1(p_0[50]), .A2(tempResult[50]), .B1(n_177), .B2(n_107), 
      .ZN(n_105));
   AOI21_X1 i_158 (.A(n_187), .B1(p_0[49]), .B2(tempResult[49]), .ZN(n_106));
   AOI21_X1 i_159 (.A(n_187), .B1(n_181), .B2(n_108), .ZN(n_107));
   INV_X1 i_160 (.A(n_109), .ZN(n_108));
   AOI21_X1 i_161 (.A(n_184), .B1(n_189), .B2(n_182), .ZN(n_109));
   OAI21_X1 i_162 (.A(n_182), .B1(p_0[48]), .B2(tempResult[48]), .ZN(n_110));
   NOR2_X1 i_163 (.A1(n_188), .A2(n_179), .ZN(n_111));
   XOR2_X1 i_164 (.A(n_175), .B(n_118), .Z(p_1[52]));
   XOR2_X1 i_165 (.A(n_117), .B(n_114), .Z(p_1[53]));
   XOR2_X1 i_166 (.A(n_115), .B(n_112), .Z(p_1[54]));
   NOR2_X1 i_167 (.A1(n_164), .A2(n_154), .ZN(n_112));
   XNOR2_X1 i_168 (.A(n_119), .B(n_113), .ZN(p_1[55]));
   OAI21_X1 i_169 (.A(n_163), .B1(n_154), .B2(n_115), .ZN(n_113));
   NOR2_X1 i_170 (.A1(n_166), .A2(n_156), .ZN(n_114));
   INV_X1 i_171 (.A(n_116), .ZN(n_115));
   OAI21_X1 i_172 (.A(n_165), .B1(n_156), .B2(n_117), .ZN(n_116));
   AOI21_X1 i_173 (.A(n_161), .B1(n_175), .B2(n_158), .ZN(n_117));
   OAI21_X1 i_174 (.A(n_158), .B1(p_0[52]), .B2(tempResult[52]), .ZN(n_118));
   AOI21_X1 i_175 (.A(n_168), .B1(p_0[55]), .B2(tempResult[55]), .ZN(n_119));
   XNOR2_X1 i_176 (.A(n_128), .B(n_127), .ZN(p_1[56]));
   XOR2_X1 i_177 (.A(n_125), .B(n_124), .Z(p_1[57]));
   XNOR2_X1 i_178 (.A(n_121), .B(n_120), .ZN(p_1[58]));
   OAI22_X1 i_179 (.A1(p_0[57]), .A2(tempResult[57]), .B1(n_149), .B2(n_125), 
      .ZN(n_120));
   NOR2_X1 i_180 (.A1(n_172), .A2(n_145), .ZN(n_121));
   XNOR2_X1 i_181 (.A(n_129), .B(n_122), .ZN(p_1[59]));
   OAI21_X1 i_182 (.A(n_123), .B1(n_171), .B2(n_145), .ZN(n_122));
   NAND3_X1 i_183 (.A1(n_146), .A2(n_124), .A3(n_126), .ZN(n_123));
   NOR2_X1 i_184 (.A1(n_173), .A2(n_149), .ZN(n_124));
   INV_X1 i_185 (.A(n_126), .ZN(n_125));
   OAI22_X1 i_186 (.A1(p_0[56]), .A2(tempResult[56]), .B1(n_150), .B2(n_128), 
      .ZN(n_126));
   OAI21_X1 i_187 (.A(n_151), .B1(p_0[56]), .B2(tempResult[56]), .ZN(n_127));
   OAI21_X1 i_188 (.A(n_153), .B1(n_175), .B2(n_160), .ZN(n_128));
   AOI21_X1 i_189 (.A(n_174), .B1(p_0[59]), .B2(tempResult[59]), .ZN(n_129));
   XNOR2_X1 i_190 (.A(n_143), .B(n_142), .ZN(p_1[60]));
   AOI22_X1 i_191 (.A1(n_140), .A2(n_136), .B1(n_141), .B2(n_135), .ZN(p_1[61]));
   XOR2_X1 i_192 (.A(n_131), .B(n_130), .Z(p_1[62]));
   AOI22_X1 i_193 (.A1(p_0[61]), .A2(tempResult[61]), .B1(n_141), .B2(n_137), 
      .ZN(n_130));
   OAI21_X1 i_194 (.A(n_139), .B1(p_0[62]), .B2(tempResult[62]), .ZN(n_131));
   XOR2_X1 i_195 (.A(n_133), .B(n_132), .Z(p_1[63]));
   XNOR2_X1 i_196 (.A(p_0[63]), .B(tempResult[63]), .ZN(n_132));
   OAI221_X1 i_197 (.A(n_134), .B1(p_0[62]), .B2(tempResult[62]), .C1(n_138), 
      .C2(n_137), .ZN(n_133));
   NAND3_X1 i_198 (.A1(n_139), .A2(n_135), .A3(n_140), .ZN(n_134));
   INV_X1 i_199 (.A(n_136), .ZN(n_135));
   OAI21_X1 i_200 (.A(n_137), .B1(n_379), .B2(n_375), .ZN(n_136));
   NAND2_X1 i_201 (.A1(n_379), .A2(n_375), .ZN(n_137));
   INV_X1 i_202 (.A(n_139), .ZN(n_138));
   NAND2_X1 i_203 (.A1(p_0[62]), .A2(tempResult[62]), .ZN(n_139));
   INV_X1 i_204 (.A(n_141), .ZN(n_140));
   AOI21_X1 i_205 (.A(n_371), .B1(n_143), .B2(n_142), .ZN(n_141));
   AOI21_X1 i_206 (.A(n_371), .B1(p_0[60]), .B2(tempResult[60]), .ZN(n_142));
   NOR4_X1 i_207 (.A1(n_147), .A2(n_144), .A3(n_152), .A4(n_159), .ZN(n_143));
   OAI22_X1 i_208 (.A1(n_378), .A2(n_374), .B1(n_174), .B2(n_146), .ZN(n_144));
   INV_X1 i_209 (.A(n_146), .ZN(n_145));
   NAND2_X1 i_210 (.A1(p_0[58]), .A2(tempResult[58]), .ZN(n_146));
   INV_X1 i_211 (.A(n_148), .ZN(n_147));
   OAI21_X1 i_212 (.A(n_170), .B1(n_150), .B2(n_149), .ZN(n_148));
   AND2_X1 i_213 (.A1(p_0[57]), .A2(tempResult[57]), .ZN(n_149));
   INV_X1 i_214 (.A(n_151), .ZN(n_150));
   NAND2_X1 i_215 (.A1(p_0[56]), .A2(tempResult[56]), .ZN(n_151));
   NOR2_X1 i_216 (.A1(n_169), .A2(n_153), .ZN(n_152));
   AOI221_X1 i_217 (.A(n_155), .B1(p_0[55]), .B2(tempResult[55]), .C1(n_167), 
      .C2(n_154), .ZN(n_153));
   AND2_X1 i_218 (.A1(p_0[54]), .A2(tempResult[54]), .ZN(n_154));
   AOI21_X1 i_219 (.A(n_162), .B1(n_158), .B2(n_157), .ZN(n_155));
   INV_X1 i_220 (.A(n_157), .ZN(n_156));
   NAND2_X1 i_221 (.A1(p_0[53]), .A2(tempResult[53]), .ZN(n_157));
   NAND2_X1 i_222 (.A1(p_0[52]), .A2(tempResult[52]), .ZN(n_158));
   NOR3_X1 i_223 (.A1(n_169), .A2(n_160), .A3(n_175), .ZN(n_159));
   OR2_X1 i_224 (.A1(n_162), .A2(n_161), .ZN(n_160));
   NOR2_X1 i_225 (.A1(p_0[52]), .A2(tempResult[52]), .ZN(n_161));
   NAND3_X1 i_226 (.A1(n_167), .A2(n_163), .A3(n_165), .ZN(n_162));
   INV_X1 i_227 (.A(n_164), .ZN(n_163));
   NOR2_X1 i_228 (.A1(p_0[54]), .A2(tempResult[54]), .ZN(n_164));
   INV_X1 i_229 (.A(n_166), .ZN(n_165));
   NOR2_X1 i_230 (.A1(p_0[53]), .A2(tempResult[53]), .ZN(n_166));
   INV_X1 i_231 (.A(n_168), .ZN(n_167));
   NOR2_X1 i_232 (.A1(p_0[55]), .A2(tempResult[55]), .ZN(n_168));
   OAI21_X1 i_233 (.A(n_170), .B1(p_0[56]), .B2(tempResult[56]), .ZN(n_169));
   NOR3_X1 i_234 (.A1(n_174), .A2(n_172), .A3(n_173), .ZN(n_170));
   NOR2_X1 i_235 (.A1(n_173), .A2(n_172), .ZN(n_171));
   NOR2_X1 i_236 (.A1(p_0[58]), .A2(tempResult[58]), .ZN(n_172));
   NOR2_X1 i_237 (.A1(p_0[57]), .A2(tempResult[57]), .ZN(n_173));
   NOR2_X1 i_238 (.A1(p_0[59]), .A2(tempResult[59]), .ZN(n_174));
   NOR4_X1 i_239 (.A1(n_179), .A2(n_176), .A3(n_180), .A4(n_183), .ZN(n_175));
   NOR2_X1 i_240 (.A1(n_188), .A2(n_178), .ZN(n_176));
   INV_X1 i_241 (.A(n_178), .ZN(n_177));
   NAND2_X1 i_242 (.A1(p_0[50]), .A2(tempResult[50]), .ZN(n_178));
   AND2_X1 i_243 (.A1(p_0[51]), .A2(tempResult[51]), .ZN(n_179));
   AOI21_X1 i_244 (.A(n_185), .B1(n_182), .B2(n_181), .ZN(n_180));
   NAND2_X1 i_245 (.A1(p_0[49]), .A2(tempResult[49]), .ZN(n_181));
   NAND2_X1 i_246 (.A1(p_0[48]), .A2(tempResult[48]), .ZN(n_182));
   NOR3_X1 i_247 (.A1(n_185), .A2(n_184), .A3(n_189), .ZN(n_183));
   NOR2_X1 i_248 (.A1(p_0[48]), .A2(tempResult[48]), .ZN(n_184));
   OR3_X1 i_249 (.A1(n_188), .A2(n_186), .A3(n_187), .ZN(n_185));
   NOR2_X1 i_250 (.A1(p_0[50]), .A2(tempResult[50]), .ZN(n_186));
   NOR2_X1 i_251 (.A1(p_0[49]), .A2(tempResult[49]), .ZN(n_187));
   NOR2_X1 i_252 (.A1(p_0[51]), .A2(tempResult[51]), .ZN(n_188));
   NOR3_X1 i_253 (.A1(n_211), .A2(n_190), .A3(n_218), .ZN(n_189));
   OAI221_X1 i_254 (.A(n_197), .B1(n_239), .B2(n_191), .C1(n_229), .C2(n_205), 
      .ZN(n_190));
   AOI221_X1 i_255 (.A(n_193), .B1(p_0[43]), .B2(tempResult[43]), .C1(n_237), 
      .C2(n_192), .ZN(n_191));
   AND2_X1 i_256 (.A1(p_0[42]), .A2(tempResult[42]), .ZN(n_192));
   AOI21_X1 i_257 (.A(n_232), .B1(n_196), .B2(n_195), .ZN(n_193));
   INV_X1 i_258 (.A(n_195), .ZN(n_194));
   NAND2_X1 i_259 (.A1(p_0[41]), .A2(tempResult[41]), .ZN(n_195));
   NAND2_X1 i_260 (.A1(p_0[40]), .A2(tempResult[40]), .ZN(n_196));
   AOI21_X1 i_261 (.A(n_198), .B1(p_0[47]), .B2(tempResult[47]), .ZN(n_197));
   OAI21_X1 i_262 (.A(n_201), .B1(n_244), .B2(n_200), .ZN(n_198));
   INV_X1 i_263 (.A(n_200), .ZN(n_199));
   NAND2_X1 i_264 (.A1(p_0[46]), .A2(tempResult[46]), .ZN(n_200));
   OAI21_X1 i_265 (.A(n_240), .B1(n_203), .B2(n_202), .ZN(n_201));
   AND2_X1 i_266 (.A1(p_0[45]), .A2(tempResult[45]), .ZN(n_202));
   INV_X1 i_267 (.A(n_204), .ZN(n_203));
   NAND2_X1 i_268 (.A1(p_0[44]), .A2(tempResult[44]), .ZN(n_204));
   AOI221_X1 i_269 (.A(n_207), .B1(p_0[39]), .B2(tempResult[39]), .C1(n_251), 
      .C2(n_206), .ZN(n_205));
   AND2_X1 i_270 (.A1(p_0[38]), .A2(tempResult[38]), .ZN(n_206));
   AOI21_X1 i_271 (.A(n_246), .B1(n_210), .B2(n_209), .ZN(n_207));
   INV_X1 i_272 (.A(n_209), .ZN(n_208));
   NAND2_X1 i_273 (.A1(p_0[37]), .A2(tempResult[37]), .ZN(n_209));
   NAND2_X1 i_274 (.A1(p_0[36]), .A2(tempResult[36]), .ZN(n_210));
   NOR2_X1 i_275 (.A1(n_228), .A2(n_212), .ZN(n_211));
   AOI221_X1 i_276 (.A(n_214), .B1(p_0[35]), .B2(tempResult[35]), .C1(n_226), 
      .C2(n_213), .ZN(n_212));
   AND2_X1 i_277 (.A1(p_0[34]), .A2(tempResult[34]), .ZN(n_213));
   AOI21_X1 i_278 (.A(n_221), .B1(n_217), .B2(n_216), .ZN(n_214));
   INV_X1 i_279 (.A(n_216), .ZN(n_215));
   NAND2_X1 i_280 (.A1(p_0[33]), .A2(tempResult[33]), .ZN(n_216));
   NAND2_X1 i_281 (.A1(p_0[32]), .A2(tempResult[32]), .ZN(n_217));
   NOR3_X1 i_282 (.A1(n_228), .A2(n_219), .A3(n_254), .ZN(n_218));
   OR2_X1 i_283 (.A1(n_221), .A2(n_220), .ZN(n_219));
   NOR2_X1 i_284 (.A1(p_0[32]), .A2(tempResult[32]), .ZN(n_220));
   NAND3_X1 i_285 (.A1(n_226), .A2(n_222), .A3(n_224), .ZN(n_221));
   INV_X1 i_286 (.A(n_223), .ZN(n_222));
   NOR2_X1 i_287 (.A1(p_0[34]), .A2(tempResult[34]), .ZN(n_223));
   INV_X1 i_288 (.A(n_225), .ZN(n_224));
   NOR2_X1 i_289 (.A1(p_0[33]), .A2(tempResult[33]), .ZN(n_225));
   INV_X1 i_290 (.A(n_227), .ZN(n_226));
   NOR2_X1 i_291 (.A1(p_0[35]), .A2(tempResult[35]), .ZN(n_227));
   OR2_X1 i_292 (.A1(n_245), .A2(n_229), .ZN(n_228));
   OR2_X1 i_293 (.A1(n_239), .A2(n_230), .ZN(n_229));
   OR2_X1 i_294 (.A1(n_232), .A2(n_231), .ZN(n_230));
   NOR2_X1 i_295 (.A1(p_0[40]), .A2(tempResult[40]), .ZN(n_231));
   NAND3_X1 i_296 (.A1(n_237), .A2(n_233), .A3(n_235), .ZN(n_232));
   INV_X1 i_297 (.A(n_234), .ZN(n_233));
   NOR2_X1 i_298 (.A1(p_0[42]), .A2(tempResult[42]), .ZN(n_234));
   INV_X1 i_299 (.A(n_236), .ZN(n_235));
   NOR2_X1 i_300 (.A1(p_0[41]), .A2(tempResult[41]), .ZN(n_236));
   INV_X1 i_301 (.A(n_238), .ZN(n_237));
   NOR2_X1 i_302 (.A1(p_0[43]), .A2(tempResult[43]), .ZN(n_238));
   OAI21_X1 i_303 (.A(n_240), .B1(p_0[44]), .B2(tempResult[44]), .ZN(n_239));
   NOR3_X1 i_304 (.A1(n_244), .A2(n_242), .A3(n_243), .ZN(n_240));
   NOR2_X1 i_305 (.A1(n_243), .A2(n_242), .ZN(n_241));
   NOR2_X1 i_306 (.A1(p_0[46]), .A2(tempResult[46]), .ZN(n_242));
   NOR2_X1 i_307 (.A1(p_0[45]), .A2(tempResult[45]), .ZN(n_243));
   NOR2_X1 i_308 (.A1(p_0[47]), .A2(tempResult[47]), .ZN(n_244));
   OR2_X1 i_309 (.A1(n_253), .A2(n_246), .ZN(n_245));
   NAND3_X1 i_310 (.A1(n_251), .A2(n_247), .A3(n_249), .ZN(n_246));
   INV_X1 i_311 (.A(n_248), .ZN(n_247));
   NOR2_X1 i_312 (.A1(p_0[38]), .A2(tempResult[38]), .ZN(n_248));
   INV_X1 i_313 (.A(n_250), .ZN(n_249));
   NOR2_X1 i_314 (.A1(p_0[37]), .A2(tempResult[37]), .ZN(n_250));
   INV_X1 i_315 (.A(n_252), .ZN(n_251));
   NOR2_X1 i_316 (.A1(p_0[39]), .A2(tempResult[39]), .ZN(n_252));
   NOR2_X1 i_317 (.A1(p_0[36]), .A2(tempResult[36]), .ZN(n_253));
   NOR3_X1 i_318 (.A1(n_262), .A2(n_255), .A3(n_280), .ZN(n_254));
   OAI222_X1 i_319 (.A1(n_290), .A2(n_274), .B1(n_291), .B2(n_256), .C1(n_301), 
      .C2(n_268), .ZN(n_255));
   AOI221_X1 i_320 (.A(n_258), .B1(p_0[23]), .B2(tempResult[23]), .C1(n_316), 
      .C2(n_257), .ZN(n_256));
   AND2_X1 i_321 (.A1(p_0[22]), .A2(tempResult[22]), .ZN(n_257));
   AOI21_X1 i_322 (.A(n_311), .B1(n_261), .B2(n_260), .ZN(n_258));
   INV_X1 i_323 (.A(n_260), .ZN(n_259));
   NAND2_X1 i_324 (.A1(p_0[21]), .A2(tempResult[21]), .ZN(n_260));
   NAND2_X1 i_325 (.A1(p_0[20]), .A2(tempResult[20]), .ZN(n_261));
   OAI222_X1 i_326 (.A1(n_303), .A2(n_265), .B1(n_309), .B2(n_264), .C1(n_377), 
      .C2(n_373), .ZN(n_262));
   INV_X1 i_327 (.A(n_264), .ZN(n_263));
   NAND2_X1 i_328 (.A1(p_0[30]), .A2(tempResult[30]), .ZN(n_264));
   AOI21_X1 i_329 (.A(n_266), .B1(p_0[28]), .B2(tempResult[28]), .ZN(n_265));
   AND2_X1 i_330 (.A1(p_0[29]), .A2(tempResult[29]), .ZN(n_266));
   NAND2_X1 i_331 (.A1(p_0[28]), .A2(tempResult[28]), .ZN(n_267));
   AOI221_X1 i_332 (.A(n_270), .B1(p_0[27]), .B2(tempResult[27]), .C1(n_299), 
      .C2(n_269), .ZN(n_268));
   AND2_X1 i_333 (.A1(p_0[26]), .A2(tempResult[26]), .ZN(n_269));
   AOI21_X1 i_334 (.A(n_294), .B1(n_273), .B2(n_272), .ZN(n_270));
   INV_X1 i_335 (.A(n_272), .ZN(n_271));
   NAND2_X1 i_336 (.A1(p_0[25]), .A2(tempResult[25]), .ZN(n_272));
   NAND2_X1 i_337 (.A1(p_0[24]), .A2(tempResult[24]), .ZN(n_273));
   AOI221_X1 i_338 (.A(n_276), .B1(p_0[19]), .B2(tempResult[19]), .C1(n_288), 
      .C2(n_275), .ZN(n_274));
   AND2_X1 i_339 (.A1(p_0[18]), .A2(tempResult[18]), .ZN(n_275));
   AOI21_X1 i_340 (.A(n_283), .B1(n_279), .B2(n_278), .ZN(n_276));
   INV_X1 i_341 (.A(n_278), .ZN(n_277));
   NAND2_X1 i_342 (.A1(p_0[17]), .A2(tempResult[17]), .ZN(n_278));
   NAND2_X1 i_343 (.A1(p_0[16]), .A2(tempResult[16]), .ZN(n_279));
   NOR3_X1 i_344 (.A1(n_290), .A2(n_281), .A3(n_319), .ZN(n_280));
   OR2_X1 i_345 (.A1(n_283), .A2(n_282), .ZN(n_281));
   NOR2_X1 i_346 (.A1(p_0[16]), .A2(tempResult[16]), .ZN(n_282));
   NAND3_X1 i_347 (.A1(n_288), .A2(n_284), .A3(n_286), .ZN(n_283));
   INV_X1 i_348 (.A(n_285), .ZN(n_284));
   NOR2_X1 i_349 (.A1(p_0[18]), .A2(tempResult[18]), .ZN(n_285));
   INV_X1 i_350 (.A(n_287), .ZN(n_286));
   NOR2_X1 i_351 (.A1(p_0[17]), .A2(tempResult[17]), .ZN(n_287));
   INV_X1 i_352 (.A(n_289), .ZN(n_288));
   NOR2_X1 i_353 (.A1(p_0[19]), .A2(tempResult[19]), .ZN(n_289));
   OR2_X1 i_354 (.A1(n_310), .A2(n_291), .ZN(n_290));
   OR2_X1 i_355 (.A1(n_301), .A2(n_292), .ZN(n_291));
   OR2_X1 i_356 (.A1(n_294), .A2(n_293), .ZN(n_292));
   NOR2_X1 i_357 (.A1(p_0[24]), .A2(tempResult[24]), .ZN(n_293));
   NAND3_X1 i_358 (.A1(n_299), .A2(n_295), .A3(n_297), .ZN(n_294));
   INV_X1 i_359 (.A(n_296), .ZN(n_295));
   NOR2_X1 i_360 (.A1(p_0[26]), .A2(tempResult[26]), .ZN(n_296));
   INV_X1 i_361 (.A(n_298), .ZN(n_297));
   NOR2_X1 i_362 (.A1(p_0[25]), .A2(tempResult[25]), .ZN(n_298));
   INV_X1 i_363 (.A(n_300), .ZN(n_299));
   NOR2_X1 i_364 (.A1(p_0[27]), .A2(tempResult[27]), .ZN(n_300));
   OR2_X1 i_365 (.A1(n_303), .A2(n_302), .ZN(n_301));
   NOR2_X1 i_366 (.A1(p_0[28]), .A2(tempResult[28]), .ZN(n_302));
   NAND3_X1 i_367 (.A1(n_308), .A2(n_304), .A3(n_306), .ZN(n_303));
   INV_X1 i_368 (.A(n_305), .ZN(n_304));
   NOR2_X1 i_369 (.A1(p_0[30]), .A2(tempResult[30]), .ZN(n_305));
   INV_X1 i_370 (.A(n_307), .ZN(n_306));
   NOR2_X1 i_371 (.A1(p_0[29]), .A2(tempResult[29]), .ZN(n_307));
   INV_X1 i_372 (.A(n_309), .ZN(n_308));
   NOR2_X1 i_373 (.A1(p_0[31]), .A2(tempResult[31]), .ZN(n_309));
   OR2_X1 i_374 (.A1(n_318), .A2(n_311), .ZN(n_310));
   NAND3_X1 i_375 (.A1(n_316), .A2(n_312), .A3(n_314), .ZN(n_311));
   INV_X1 i_376 (.A(n_313), .ZN(n_312));
   NOR2_X1 i_377 (.A1(p_0[22]), .A2(tempResult[22]), .ZN(n_313));
   INV_X1 i_378 (.A(n_315), .ZN(n_314));
   NOR2_X1 i_379 (.A1(p_0[21]), .A2(tempResult[21]), .ZN(n_315));
   INV_X1 i_380 (.A(n_317), .ZN(n_316));
   NOR2_X1 i_381 (.A1(p_0[23]), .A2(tempResult[23]), .ZN(n_317));
   NOR2_X1 i_382 (.A1(p_0[20]), .A2(tempResult[20]), .ZN(n_318));
   NOR4_X1 i_383 (.A1(n_323), .A2(n_320), .A3(n_324), .A4(n_327), .ZN(n_319));
   NOR2_X1 i_384 (.A1(n_332), .A2(n_322), .ZN(n_320));
   INV_X1 i_385 (.A(n_322), .ZN(n_321));
   NAND2_X1 i_386 (.A1(p_0[14]), .A2(tempResult[14]), .ZN(n_322));
   AND2_X1 i_387 (.A1(p_0[15]), .A2(tempResult[15]), .ZN(n_323));
   AOI21_X1 i_388 (.A(n_329), .B1(n_326), .B2(n_325), .ZN(n_324));
   NAND2_X1 i_389 (.A1(p_0[13]), .A2(tempResult[13]), .ZN(n_325));
   NAND2_X1 i_390 (.A1(p_0[12]), .A2(tempResult[12]), .ZN(n_326));
   NOR3_X1 i_391 (.A1(n_329), .A2(n_328), .A3(n_333), .ZN(n_327));
   NOR2_X1 i_392 (.A1(p_0[12]), .A2(tempResult[12]), .ZN(n_328));
   OR3_X1 i_393 (.A1(n_332), .A2(n_330), .A3(n_331), .ZN(n_329));
   NOR2_X1 i_394 (.A1(p_0[14]), .A2(tempResult[14]), .ZN(n_330));
   NOR2_X1 i_395 (.A1(p_0[13]), .A2(tempResult[13]), .ZN(n_331));
   NOR2_X1 i_396 (.A1(p_0[15]), .A2(tempResult[15]), .ZN(n_332));
   NOR4_X1 i_397 (.A1(n_337), .A2(n_334), .A3(n_338), .A4(n_341), .ZN(n_333));
   NOR2_X1 i_398 (.A1(n_346), .A2(n_336), .ZN(n_334));
   INV_X1 i_399 (.A(n_336), .ZN(n_335));
   NAND2_X1 i_400 (.A1(p_0[10]), .A2(tempResult[10]), .ZN(n_336));
   AND2_X1 i_401 (.A1(p_0[11]), .A2(tempResult[11]), .ZN(n_337));
   AOI21_X1 i_402 (.A(n_343), .B1(n_340), .B2(n_339), .ZN(n_338));
   NAND2_X1 i_403 (.A1(p_0[9]), .A2(tempResult[9]), .ZN(n_339));
   NAND2_X1 i_404 (.A1(p_0[8]), .A2(tempResult[8]), .ZN(n_340));
   NOR3_X1 i_405 (.A1(n_343), .A2(n_342), .A3(n_347), .ZN(n_341));
   NOR2_X1 i_406 (.A1(p_0[8]), .A2(tempResult[8]), .ZN(n_342));
   OR3_X1 i_407 (.A1(n_346), .A2(n_344), .A3(n_345), .ZN(n_343));
   NOR2_X1 i_408 (.A1(p_0[10]), .A2(tempResult[10]), .ZN(n_344));
   NOR2_X1 i_409 (.A1(p_0[9]), .A2(tempResult[9]), .ZN(n_345));
   NOR2_X1 i_410 (.A1(p_0[11]), .A2(tempResult[11]), .ZN(n_346));
   NOR4_X1 i_411 (.A1(n_351), .A2(n_348), .A3(n_352), .A4(n_355), .ZN(n_347));
   NOR2_X1 i_412 (.A1(n_360), .A2(n_350), .ZN(n_348));
   INV_X1 i_413 (.A(n_350), .ZN(n_349));
   NAND2_X1 i_414 (.A1(p_0[6]), .A2(tempResult[6]), .ZN(n_350));
   AND2_X1 i_415 (.A1(p_0[7]), .A2(tempResult[7]), .ZN(n_351));
   AOI21_X1 i_416 (.A(n_357), .B1(n_354), .B2(n_353), .ZN(n_352));
   NAND2_X1 i_417 (.A1(p_0[5]), .A2(tempResult[5]), .ZN(n_353));
   NAND2_X1 i_418 (.A1(p_0[4]), .A2(tempResult[4]), .ZN(n_354));
   NOR3_X1 i_419 (.A1(n_357), .A2(n_356), .A3(n_361), .ZN(n_355));
   NOR2_X1 i_420 (.A1(p_0[4]), .A2(tempResult[4]), .ZN(n_356));
   OR3_X1 i_421 (.A1(n_360), .A2(n_358), .A3(n_359), .ZN(n_357));
   NOR2_X1 i_422 (.A1(p_0[6]), .A2(tempResult[6]), .ZN(n_358));
   NOR2_X1 i_423 (.A1(p_0[5]), .A2(tempResult[5]), .ZN(n_359));
   NOR2_X1 i_424 (.A1(p_0[7]), .A2(tempResult[7]), .ZN(n_360));
   NAND2_X1 i_425 (.A1(n_370), .A2(n_362), .ZN(n_361));
   OAI21_X1 i_426 (.A(n_363), .B1(n_376), .B2(n_372), .ZN(n_362));
   OAI22_X1 i_427 (.A1(p_0[2]), .A2(tempResult[2]), .B1(n_368), .B2(n_364), 
      .ZN(n_363));
   AOI21_X1 i_428 (.A(n_367), .B1(n_366), .B2(n_365), .ZN(n_364));
   NAND2_X1 i_429 (.A1(p_0[1]), .A2(tempResult[1]), .ZN(n_365));
   NAND2_X1 i_430 (.A1(p_0[0]), .A2(tempResult[0]), .ZN(n_366));
   NOR2_X1 i_431 (.A1(p_0[1]), .A2(tempResult[1]), .ZN(n_367));
   INV_X1 i_432 (.A(n_369), .ZN(n_368));
   NAND2_X1 i_433 (.A1(p_0[2]), .A2(tempResult[2]), .ZN(n_369));
   NAND2_X1 i_434 (.A1(n_376), .A2(n_372), .ZN(n_370));
   NOR2_X1 i_435 (.A1(p_0[60]), .A2(tempResult[60]), .ZN(n_371));
   INV_X1 i_436 (.A(tempResult[3]), .ZN(n_372));
   INV_X1 i_437 (.A(tempResult[31]), .ZN(n_373));
   INV_X1 i_438 (.A(tempResult[59]), .ZN(n_374));
   INV_X1 i_439 (.A(tempResult[61]), .ZN(n_375));
   INV_X1 i_440 (.A(p_0[3]), .ZN(n_376));
   INV_X1 i_441 (.A(p_0[31]), .ZN(n_377));
   INV_X1 i_442 (.A(p_0[59]), .ZN(n_378));
   INV_X1 i_443 (.A(p_0[61]), .ZN(n_379));
endmodule

module Noaman_4_Booth(start, clk, in1, in2, result);
   input start;
   input clk;
   input [31:0]in1;
   input [31:0]in2;
   output [63:0]result;

   wire n_0_3;
   wire n_0_0;
   wire n_0_4;
   wire n_0_1;
   wire n_0_5;
   wire n_0_2;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_316__0;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_318__0;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_320__0;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_321__0;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_322__0;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_323__0;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_324__0;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_325__0;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_326__0;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_327__0;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_328__0;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_329__0;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_330__0;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_331__0;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_332__0;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_333__0;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_334__0;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_335__0;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_336__0;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_337__0;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_338__0;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_339__0;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_340__0;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_341__0;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_342__0;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_343__0;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_344__0;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_345__0;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_346__0;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_347__0;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_348__0;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_349__0;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_350__0;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_351__0;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_352__0;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_353__0;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_354__0;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_355__0;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_356__0;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_357__0;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_358__0;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_359__0;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_360__0;
   wire n_0_316__1;
   wire n_0_317;
   wire n_0_318__1;
   wire n_0_361__0;
   wire n_0_319;
   wire n_0_320__1;
   wire n_0_321__1;
   wire n_0_362__0;
   wire n_0_322__1;
   wire n_0_323__1;
   wire n_0_324__1;
   wire n_0_363__0;
   wire n_0_325__1;
   wire n_0_326__1;
   wire n_0_327__1;
   wire n_0_364__0;
   wire n_0_328__1;
   wire n_0_329__1;
   wire n_0_330__1;
   wire n_0_365__0;
   wire n_0_331__1;
   wire n_0_332__1;
   wire n_0_333__1;
   wire n_0_334__1;
   wire n_0_335__1;
   wire n_0_366__0;
   wire n_0_336__1;
   wire n_0_337__1;
   wire n_0_338__1;
   wire n_0_367__0;
   wire n_0_339__1;
   wire n_0_340__1;
   wire n_0_341__1;
   wire n_0_368__0;
   wire n_0_342__1;
   wire n_0_343__1;
   wire n_0_344__1;
   wire n_0_369__0;
   wire n_0_345__1;
   wire n_0_346__1;
   wire n_0_347__1;
   wire n_0_370__0;
   wire n_0_348__1;
   wire n_0_349__1;
   wire n_0_350__1;
   wire n_0_371__0;
   wire n_0_351__1;
   wire n_0_352__1;
   wire n_0_353__1;
   wire n_0_372;
   wire n_0_354__1;
   wire n_0_355__1;
   wire n_0_356__1;
   wire n_0_373;
   wire n_0_357__1;
   wire n_0_358__1;
   wire n_0_359__1;
   wire n_0_374;
   wire n_0_360__1;
   wire n_0_361__1;
   wire n_0_362__1;
   wire n_0_375;
   wire n_0_363__1;
   wire n_0_364__1;
   wire n_0_365__1;
   wire n_0_376;
   wire n_0_366__1;
   wire n_0_367__1;
   wire n_0_368__1;
   wire n_0_377;
   wire n_0_369__1;
   wire n_0_381;
   wire n_0_370__1;
   wire n_0_378;
   wire n_0_379;
   wire n_0_371__1;
   wire n_0_380;
   wire [63:0]tempResult;
   wire [5:0]shiftingAmount;
   wire [34:0]newB;
   wire [63:0]Input1_1_Negative;
   wire [63:0]Input1_1_Positive;
   wire [63:0]Input1_2_Negative;
   wire [63:0]Input1_2_Positive;

   CLKGATETST_X1 clk_gate_result_reg (.CK(clk), .E(n_168), .SE(1'b0), .GCK(n_0));
   DFF_X1 \result_reg[63]  (.D(tempResult[63]), .CK(n_0), .Q(result[63]), .QN());
   DFF_X1 \result_reg[62]  (.D(tempResult[62]), .CK(n_0), .Q(result[62]), .QN());
   DFF_X1 \result_reg[61]  (.D(tempResult[61]), .CK(n_0), .Q(result[61]), .QN());
   DFF_X1 \result_reg[60]  (.D(tempResult[60]), .CK(n_0), .Q(result[60]), .QN());
   DFF_X1 \result_reg[59]  (.D(tempResult[59]), .CK(n_0), .Q(result[59]), .QN());
   DFF_X1 \result_reg[58]  (.D(tempResult[58]), .CK(n_0), .Q(result[58]), .QN());
   DFF_X1 \result_reg[57]  (.D(tempResult[57]), .CK(n_0), .Q(result[57]), .QN());
   DFF_X1 \result_reg[56]  (.D(tempResult[56]), .CK(n_0), .Q(result[56]), .QN());
   DFF_X1 \result_reg[55]  (.D(tempResult[55]), .CK(n_0), .Q(result[55]), .QN());
   DFF_X1 \result_reg[54]  (.D(tempResult[54]), .CK(n_0), .Q(result[54]), .QN());
   DFF_X1 \result_reg[53]  (.D(tempResult[53]), .CK(n_0), .Q(result[53]), .QN());
   DFF_X1 \result_reg[52]  (.D(tempResult[52]), .CK(n_0), .Q(result[52]), .QN());
   DFF_X1 \result_reg[51]  (.D(tempResult[51]), .CK(n_0), .Q(result[51]), .QN());
   DFF_X1 \result_reg[50]  (.D(tempResult[50]), .CK(n_0), .Q(result[50]), .QN());
   DFF_X1 \result_reg[49]  (.D(tempResult[49]), .CK(n_0), .Q(result[49]), .QN());
   DFF_X1 \result_reg[48]  (.D(tempResult[48]), .CK(n_0), .Q(result[48]), .QN());
   DFF_X1 \result_reg[47]  (.D(tempResult[47]), .CK(n_0), .Q(result[47]), .QN());
   DFF_X1 \result_reg[46]  (.D(tempResult[46]), .CK(n_0), .Q(result[46]), .QN());
   DFF_X1 \result_reg[45]  (.D(tempResult[45]), .CK(n_0), .Q(result[45]), .QN());
   DFF_X1 \result_reg[44]  (.D(tempResult[44]), .CK(n_0), .Q(result[44]), .QN());
   DFF_X1 \result_reg[43]  (.D(tempResult[43]), .CK(n_0), .Q(result[43]), .QN());
   DFF_X1 \result_reg[42]  (.D(tempResult[42]), .CK(n_0), .Q(result[42]), .QN());
   DFF_X1 \result_reg[41]  (.D(tempResult[41]), .CK(n_0), .Q(result[41]), .QN());
   DFF_X1 \result_reg[40]  (.D(tempResult[40]), .CK(n_0), .Q(result[40]), .QN());
   DFF_X1 \result_reg[39]  (.D(tempResult[39]), .CK(n_0), .Q(result[39]), .QN());
   DFF_X1 \result_reg[38]  (.D(tempResult[38]), .CK(n_0), .Q(result[38]), .QN());
   DFF_X1 \result_reg[37]  (.D(tempResult[37]), .CK(n_0), .Q(result[37]), .QN());
   DFF_X1 \result_reg[36]  (.D(tempResult[36]), .CK(n_0), .Q(result[36]), .QN());
   DFF_X1 \result_reg[35]  (.D(tempResult[35]), .CK(n_0), .Q(result[35]), .QN());
   DFF_X1 \result_reg[34]  (.D(tempResult[34]), .CK(n_0), .Q(result[34]), .QN());
   DFF_X1 \result_reg[33]  (.D(tempResult[33]), .CK(n_0), .Q(result[33]), .QN());
   DFF_X1 \result_reg[32]  (.D(tempResult[32]), .CK(n_0), .Q(result[32]), .QN());
   DFF_X1 \result_reg[31]  (.D(tempResult[31]), .CK(n_0), .Q(result[31]), .QN());
   DFF_X1 \result_reg[30]  (.D(tempResult[30]), .CK(n_0), .Q(result[30]), .QN());
   DFF_X1 \result_reg[29]  (.D(tempResult[29]), .CK(n_0), .Q(result[29]), .QN());
   DFF_X1 \result_reg[28]  (.D(tempResult[28]), .CK(n_0), .Q(result[28]), .QN());
   DFF_X1 \result_reg[27]  (.D(tempResult[27]), .CK(n_0), .Q(result[27]), .QN());
   DFF_X1 \result_reg[26]  (.D(tempResult[26]), .CK(n_0), .Q(result[26]), .QN());
   DFF_X1 \result_reg[25]  (.D(tempResult[25]), .CK(n_0), .Q(result[25]), .QN());
   DFF_X1 \result_reg[24]  (.D(tempResult[24]), .CK(n_0), .Q(result[24]), .QN());
   DFF_X1 \result_reg[23]  (.D(tempResult[23]), .CK(n_0), .Q(result[23]), .QN());
   DFF_X1 \result_reg[22]  (.D(tempResult[22]), .CK(n_0), .Q(result[22]), .QN());
   DFF_X1 \result_reg[21]  (.D(tempResult[21]), .CK(n_0), .Q(result[21]), .QN());
   DFF_X1 \result_reg[20]  (.D(tempResult[20]), .CK(n_0), .Q(result[20]), .QN());
   DFF_X1 \result_reg[19]  (.D(tempResult[19]), .CK(n_0), .Q(result[19]), .QN());
   DFF_X1 \result_reg[18]  (.D(tempResult[18]), .CK(n_0), .Q(result[18]), .QN());
   DFF_X1 \result_reg[17]  (.D(tempResult[17]), .CK(n_0), .Q(result[17]), .QN());
   DFF_X1 \result_reg[16]  (.D(tempResult[16]), .CK(n_0), .Q(result[16]), .QN());
   DFF_X1 \result_reg[15]  (.D(tempResult[15]), .CK(n_0), .Q(result[15]), .QN());
   DFF_X1 \result_reg[14]  (.D(tempResult[14]), .CK(n_0), .Q(result[14]), .QN());
   DFF_X1 \result_reg[13]  (.D(tempResult[13]), .CK(n_0), .Q(result[13]), .QN());
   DFF_X1 \result_reg[12]  (.D(tempResult[12]), .CK(n_0), .Q(result[12]), .QN());
   DFF_X1 \result_reg[11]  (.D(tempResult[11]), .CK(n_0), .Q(result[11]), .QN());
   DFF_X1 \result_reg[10]  (.D(tempResult[10]), .CK(n_0), .Q(result[10]), .QN());
   DFF_X1 \result_reg[9]  (.D(tempResult[9]), .CK(n_0), .Q(result[9]), .QN());
   DFF_X1 \result_reg[8]  (.D(tempResult[8]), .CK(n_0), .Q(result[8]), .QN());
   DFF_X1 \result_reg[7]  (.D(tempResult[7]), .CK(n_0), .Q(result[7]), .QN());
   DFF_X1 \result_reg[6]  (.D(tempResult[6]), .CK(n_0), .Q(result[6]), .QN());
   DFF_X1 \result_reg[5]  (.D(tempResult[5]), .CK(n_0), .Q(result[5]), .QN());
   DFF_X1 \result_reg[4]  (.D(tempResult[4]), .CK(n_0), .Q(result[4]), .QN());
   DFF_X1 \result_reg[3]  (.D(tempResult[3]), .CK(n_0), .Q(result[3]), .QN());
   DFF_X1 \result_reg[2]  (.D(tempResult[2]), .CK(n_0), .Q(result[2]), .QN());
   DFF_X1 \result_reg[1]  (.D(tempResult[1]), .CK(n_0), .Q(result[1]), .QN());
   DFF_X1 \result_reg[0]  (.D(tempResult[0]), .CK(n_0), .Q(result[0]), .QN());
   datapath__0_0 i_2 (.p_0({n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
      n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
      n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, uc_0, uc_1}), 
      .p_1({in1[31], in1[30], in1[29], in1[28], in1[27], in1[26], in1[25], 
      in1[24], in1[23], in1[22], in1[21], in1[20], in1[19], in1[18], in1[17], 
      in1[16], in1[15], in1[14], in1[13], in1[12], in1[11], in1[10], in1[9], 
      in1[8], in1[7], in1[6], in1[5], in1[4], in1[3], in1[2], in1[1], in1[0], 
      1'b0}));
   datapath__0_12 i_12 (.p_0({n_0_381, n_0_380, n_0_379, n_0_378, n_0_377, 
      n_0_376, n_0_375, n_0_374, n_0_373, n_0_372, n_0_371__0, n_0_370__0, 
      n_0_369__0, n_0_368__0, n_0_367__0, n_0_366__0, n_0_365__0, n_0_364__0, 
      n_0_363__0, n_0_362__0, n_0_361__0, n_0_360__0, n_0_359__0, n_0_358__0, 
      n_0_357__0, n_0_356__0, n_0_355__0, n_0_354__0, n_0_353__0, n_0_352__0, 
      n_0_351__0, n_0_350__0, n_0_349__0, n_0_348__0, n_0_347__0, n_0_346__0, 
      n_0_345__0, n_0_344__0, n_0_343__0, n_0_342__0, n_0_341__0, n_0_340__0, 
      n_0_339__0, n_0_338__0, n_0_337__0, n_0_336__0, n_0_335__0, n_0_334__0, 
      n_0_333__0, n_0_332__0, n_0_331__0, n_0_330__0, n_0_329__0, n_0_328__0, 
      n_0_327__0, n_0_326__0, n_0_325__0, n_0_324__0, n_0_323__0, n_0_322__0, 
      n_0_321__0, n_0_320__0, n_0_318__0, n_0_316__0}), .tempResult(tempResult), 
      .p_1({n_95, n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
      n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, 
      n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_32, n_31, n_30, 
      n_29, n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, 
      n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, 
      n_4, n_3, n_2, n_1}));
   HA_X1 i_0_0 (.A(shiftingAmount[2]), .B(shiftingAmount[1]), .CO(n_0_0), 
      .S(n_0_3));
   HA_X1 i_0_1 (.A(shiftingAmount[3]), .B(n_0_0), .CO(n_0_1), .S(n_0_4));
   HA_X1 i_0_2 (.A(shiftingAmount[4]), .B(n_0_1), .CO(n_0_2), .S(n_0_5));
   INV_X1 i_0_3 (.A(start), .ZN(n_0_6));
   AND2_X1 i_0_4 (.A1(n_0_6), .A2(n_1), .ZN(n_96));
   AND2_X1 i_0_5 (.A1(n_0_6), .A2(n_2), .ZN(n_97));
   AND2_X1 i_0_6 (.A1(n_0_6), .A2(n_3), .ZN(n_98));
   AND2_X1 i_0_7 (.A1(n_0_6), .A2(n_4), .ZN(n_99));
   AND2_X1 i_0_8 (.A1(n_0_6), .A2(n_5), .ZN(n_100));
   AND2_X1 i_0_9 (.A1(n_0_6), .A2(n_6), .ZN(n_101));
   AND2_X1 i_0_10 (.A1(n_0_6), .A2(n_7), .ZN(n_102));
   AND2_X1 i_0_11 (.A1(n_0_6), .A2(n_8), .ZN(n_103));
   AND2_X1 i_0_12 (.A1(n_0_6), .A2(n_9), .ZN(n_104));
   AND2_X1 i_0_13 (.A1(n_0_6), .A2(n_10), .ZN(n_105));
   AND2_X1 i_0_14 (.A1(n_0_6), .A2(n_11), .ZN(n_106));
   AND2_X1 i_0_15 (.A1(n_0_6), .A2(n_12), .ZN(n_107));
   AND2_X1 i_0_16 (.A1(n_0_6), .A2(n_13), .ZN(n_108));
   AND2_X1 i_0_17 (.A1(n_0_6), .A2(n_14), .ZN(n_109));
   AND2_X1 i_0_18 (.A1(n_0_6), .A2(n_15), .ZN(n_110));
   AND2_X1 i_0_19 (.A1(n_0_6), .A2(n_16), .ZN(n_111));
   AND2_X1 i_0_20 (.A1(n_0_6), .A2(n_17), .ZN(n_112));
   AND2_X1 i_0_21 (.A1(n_0_6), .A2(n_18), .ZN(n_113));
   AND2_X1 i_0_22 (.A1(n_0_6), .A2(n_19), .ZN(n_114));
   AND2_X1 i_0_23 (.A1(n_0_6), .A2(n_20), .ZN(n_115));
   AND2_X1 i_0_24 (.A1(n_0_6), .A2(n_21), .ZN(n_116));
   AND2_X1 i_0_25 (.A1(n_0_6), .A2(n_22), .ZN(n_117));
   AND2_X1 i_0_26 (.A1(n_0_6), .A2(n_23), .ZN(n_118));
   AND2_X1 i_0_27 (.A1(n_0_6), .A2(n_24), .ZN(n_119));
   AND2_X1 i_0_28 (.A1(n_0_6), .A2(n_25), .ZN(n_120));
   AND2_X1 i_0_29 (.A1(n_0_6), .A2(n_26), .ZN(n_121));
   AND2_X1 i_0_30 (.A1(n_0_6), .A2(n_27), .ZN(n_122));
   AND2_X1 i_0_31 (.A1(n_0_6), .A2(n_28), .ZN(n_123));
   AND2_X1 i_0_32 (.A1(n_0_6), .A2(n_29), .ZN(n_124));
   AND2_X1 i_0_33 (.A1(n_0_6), .A2(n_30), .ZN(n_125));
   AND2_X1 i_0_34 (.A1(n_0_6), .A2(n_31), .ZN(n_126));
   AND2_X1 i_0_35 (.A1(n_0_6), .A2(n_32), .ZN(n_127));
   AND2_X1 i_0_36 (.A1(n_0_6), .A2(n_64), .ZN(n_128));
   AND2_X1 i_0_37 (.A1(n_0_6), .A2(n_65), .ZN(n_129));
   AND2_X1 i_0_38 (.A1(n_0_6), .A2(n_66), .ZN(n_130));
   AND2_X1 i_0_39 (.A1(n_0_6), .A2(n_67), .ZN(n_131));
   AND2_X1 i_0_40 (.A1(n_0_6), .A2(n_68), .ZN(n_132));
   AND2_X1 i_0_41 (.A1(n_0_6), .A2(n_69), .ZN(n_133));
   AND2_X1 i_0_42 (.A1(n_0_6), .A2(n_70), .ZN(n_134));
   AND2_X1 i_0_43 (.A1(n_0_6), .A2(n_71), .ZN(n_135));
   AND2_X1 i_0_44 (.A1(n_0_6), .A2(n_72), .ZN(n_136));
   AND2_X1 i_0_45 (.A1(n_0_6), .A2(n_73), .ZN(n_137));
   AND2_X1 i_0_46 (.A1(n_0_6), .A2(n_74), .ZN(n_138));
   AND2_X1 i_0_47 (.A1(n_0_6), .A2(n_75), .ZN(n_139));
   AND2_X1 i_0_48 (.A1(n_0_6), .A2(n_76), .ZN(n_140));
   AND2_X1 i_0_49 (.A1(n_0_6), .A2(n_77), .ZN(n_141));
   AND2_X1 i_0_50 (.A1(n_0_6), .A2(n_78), .ZN(n_142));
   AND2_X1 i_0_51 (.A1(n_0_6), .A2(n_79), .ZN(n_143));
   AND2_X1 i_0_52 (.A1(n_0_6), .A2(n_80), .ZN(n_144));
   AND2_X1 i_0_53 (.A1(n_0_6), .A2(n_81), .ZN(n_148));
   AND2_X1 i_0_54 (.A1(n_0_6), .A2(n_82), .ZN(n_149));
   AND2_X1 i_0_55 (.A1(n_0_6), .A2(n_83), .ZN(n_150));
   AND2_X1 i_0_56 (.A1(n_0_6), .A2(n_84), .ZN(n_151));
   AND2_X1 i_0_57 (.A1(n_0_6), .A2(n_85), .ZN(n_152));
   AND2_X1 i_0_58 (.A1(n_0_6), .A2(n_86), .ZN(n_153));
   AND2_X1 i_0_59 (.A1(n_0_6), .A2(n_87), .ZN(n_154));
   AND2_X1 i_0_60 (.A1(n_0_6), .A2(n_88), .ZN(n_155));
   AND2_X1 i_0_61 (.A1(n_0_6), .A2(n_89), .ZN(n_156));
   AND2_X1 i_0_62 (.A1(n_0_6), .A2(n_90), .ZN(n_157));
   AND2_X1 i_0_63 (.A1(n_0_6), .A2(n_91), .ZN(n_158));
   AND2_X1 i_0_64 (.A1(n_0_6), .A2(n_92), .ZN(n_159));
   AND2_X1 i_0_65 (.A1(n_0_6), .A2(n_93), .ZN(n_160));
   AND2_X1 i_0_66 (.A1(n_0_6), .A2(n_94), .ZN(n_161));
   AND2_X1 i_0_67 (.A1(n_0_6), .A2(n_95), .ZN(n_162));
   NOR2_X1 i_0_68 (.A1(start), .A2(shiftingAmount[1]), .ZN(n_163));
   AND2_X1 i_0_69 (.A1(n_0_6), .A2(n_0_3), .ZN(n_164));
   AND2_X1 i_0_70 (.A1(n_0_6), .A2(n_0_4), .ZN(n_165));
   AND2_X1 i_0_71 (.A1(n_0_6), .A2(n_0_5), .ZN(n_166));
   INV_X1 i_0_72 (.A(n_0_2), .ZN(n_0_7));
   INV_X1 i_0_73 (.A(shiftingAmount[5]), .ZN(n_0_8));
   AOI221_X1 i_0_74 (.A(start), .B1(n_0_2), .B2(shiftingAmount[5]), .C1(n_0_7), 
      .C2(n_0_8), .ZN(n_167));
   NOR2_X1 i_0_75 (.A1(shiftingAmount[4]), .A2(shiftingAmount[3]), .ZN(n_0_9));
   NAND2_X1 i_0_76 (.A1(n_0_9), .A2(shiftingAmount[5]), .ZN(n_0_10));
   NOR2_X1 i_0_77 (.A1(shiftingAmount[2]), .A2(shiftingAmount[1]), .ZN(n_0_11));
   INV_X1 i_0_78 (.A(n_0_11), .ZN(n_0_12));
   NOR3_X1 i_0_79 (.A1(n_0_10), .A2(start), .A3(n_0_12), .ZN(n_168));
   INV_X1 i_0_80 (.A(newB[34]), .ZN(n_0_13));
   OR3_X1 i_0_81 (.A1(n_0_10), .A2(n_0_12), .A3(n_0_13), .ZN(n_0_14));
   NAND2_X1 i_0_82 (.A1(n_0_8), .A2(shiftingAmount[4]), .ZN(n_0_15));
   INV_X1 i_0_83 (.A(n_0_15), .ZN(n_0_16));
   INV_X1 i_0_84 (.A(shiftingAmount[3]), .ZN(n_0_17));
   NAND4_X1 i_0_85 (.A1(n_0_16), .A2(n_0_11), .A3(newB[17]), .A4(n_0_17), 
      .ZN(n_0_18));
   NAND3_X1 i_0_86 (.A1(n_0_9), .A2(n_0_11), .A3(newB[1]), .ZN(n_0_19));
   INV_X1 i_0_87 (.A(shiftingAmount[2]), .ZN(n_0_20));
   NAND2_X1 i_0_88 (.A1(n_0_20), .A2(shiftingAmount[1]), .ZN(n_0_21));
   INV_X1 i_0_89 (.A(n_0_21), .ZN(n_0_22));
   NAND2_X1 i_0_90 (.A1(n_0_22), .A2(shiftingAmount[4]), .ZN(n_0_23));
   OAI22_X1 i_0_91 (.A1(n_0_17), .A2(newB[27]), .B1(newB[19]), .B2(
      shiftingAmount[3]), .ZN(n_0_24));
   NOR2_X1 i_0_92 (.A1(n_0_17), .A2(shiftingAmount[4]), .ZN(n_0_25));
   AOI22_X1 i_0_93 (.A1(n_0_25), .A2(newB[11]), .B1(n_0_9), .B2(newB[3]), 
      .ZN(n_0_26));
   OAI221_X1 i_0_94 (.A(n_0_19), .B1(n_0_23), .B2(n_0_24), .C1(n_0_26), .C2(
      n_0_21), .ZN(n_0_27));
   INV_X1 i_0_95 (.A(shiftingAmount[4]), .ZN(n_0_28));
   NAND2_X1 i_0_96 (.A1(n_0_17), .A2(shiftingAmount[2]), .ZN(n_0_29));
   INV_X1 i_0_97 (.A(n_0_29), .ZN(n_0_30));
   NAND2_X1 i_0_98 (.A1(n_0_20), .A2(shiftingAmount[3]), .ZN(n_0_31));
   INV_X1 i_0_99 (.A(n_0_31), .ZN(n_0_32));
   AOI221_X1 i_0_100 (.A(n_0_28), .B1(n_0_30), .B2(newB[21]), .C1(newB[25]), 
      .C2(n_0_32), .ZN(n_0_33));
   NOR2_X1 i_0_101 (.A1(n_0_17), .A2(n_0_20), .ZN(n_0_34));
   AOI221_X1 i_0_102 (.A(shiftingAmount[4]), .B1(n_0_32), .B2(newB[9]), .C1(
      newB[13]), .C2(n_0_34), .ZN(n_0_35));
   AND3_X1 i_0_103 (.A1(newB[29]), .A2(shiftingAmount[4]), .A3(shiftingAmount[3]), 
      .ZN(n_0_36));
   AOI211_X1 i_0_104 (.A(shiftingAmount[1]), .B(n_0_36), .C1(newB[5]), .C2(n_0_9), 
      .ZN(n_0_37));
   INV_X1 i_0_105 (.A(shiftingAmount[1]), .ZN(n_0_38));
   AOI221_X1 i_0_106 (.A(n_0_38), .B1(n_0_9), .B2(newB[7]), .C1(n_0_25), 
      .C2(newB[15]), .ZN(n_0_39));
   OAI33_X1 i_0_107 (.A1(n_0_33), .A2(n_0_35), .A3(shiftingAmount[1]), .B1(
      n_0_37), .B2(n_0_39), .B3(n_0_20), .ZN(n_0_40));
   AOI22_X1 i_0_108 (.A1(n_0_34), .A2(newB[31]), .B1(n_0_30), .B2(newB[23]), 
      .ZN(n_0_41));
   NOR2_X1 i_0_109 (.A1(n_0_41), .A2(n_0_28), .ZN(n_0_42));
   AOI211_X1 i_0_110 (.A(n_0_27), .B(n_0_40), .C1(shiftingAmount[1]), .C2(n_0_42), 
      .ZN(n_0_43));
   OAI211_X1 i_0_111 (.A(n_0_14), .B(n_0_18), .C1(n_0_43), .C2(shiftingAmount[5]), 
      .ZN(n_0_44));
   AOI22_X1 i_0_112 (.A1(n_0_17), .A2(newB[18]), .B1(newB[26]), .B2(
      shiftingAmount[3]), .ZN(n_0_45));
   OAI33_X1 i_0_113 (.A1(n_0_10), .A2(n_0_13), .A3(shiftingAmount[2]), .B1(
      n_0_45), .B2(n_0_15), .B3(n_0_21), .ZN(n_0_46));
   AOI22_X1 i_0_114 (.A1(n_0_34), .A2(newB[14]), .B1(n_0_30), .B2(newB[6]), 
      .ZN(n_0_47));
   AOI22_X1 i_0_115 (.A1(n_0_34), .A2(newB[30]), .B1(n_0_30), .B2(newB[22]), 
      .ZN(n_0_48));
   AOI22_X1 i_0_116 (.A1(n_0_25), .A2(newB[10]), .B1(n_0_9), .B2(newB[2]), 
      .ZN(n_0_49));
   OAI222_X1 i_0_117 (.A1(shiftingAmount[4]), .A2(n_0_47), .B1(n_0_48), .B2(
      n_0_28), .C1(n_0_49), .C2(shiftingAmount[2]), .ZN(n_0_50));
   INV_X1 i_0_118 (.A(n_0_50), .ZN(n_0_51));
   NAND2_X1 i_0_119 (.A1(n_0_25), .A2(newB[8]), .ZN(n_0_52));
   OAI22_X1 i_0_120 (.A1(n_0_51), .A2(n_0_38), .B1(n_0_12), .B2(n_0_52), 
      .ZN(n_0_53));
   INV_X1 i_0_121 (.A(newB[24]), .ZN(n_0_54));
   INV_X1 i_0_122 (.A(newB[16]), .ZN(n_0_55));
   AOI221_X1 i_0_123 (.A(shiftingAmount[2]), .B1(n_0_54), .B2(shiftingAmount[3]), 
      .C1(n_0_55), .C2(n_0_17), .ZN(n_0_56));
   AOI221_X1 i_0_124 (.A(n_0_56), .B1(newB[20]), .B2(n_0_30), .C1(newB[28]), 
      .C2(n_0_34), .ZN(n_0_57));
   NOR2_X1 i_0_125 (.A1(shiftingAmount[3]), .A2(shiftingAmount[5]), .ZN(n_0_58));
   INV_X1 i_0_126 (.A(n_0_58), .ZN(n_0_59));
   NOR2_X1 i_0_127 (.A1(n_0_59), .A2(shiftingAmount[4]), .ZN(n_0_60));
   NAND2_X1 i_0_128 (.A1(n_0_8), .A2(shiftingAmount[3]), .ZN(n_0_61));
   NOR2_X1 i_0_129 (.A1(n_0_61), .A2(shiftingAmount[4]), .ZN(n_0_62));
   AOI22_X1 i_0_130 (.A1(newB[4]), .A2(n_0_60), .B1(n_0_62), .B2(newB[12]), 
      .ZN(n_0_63));
   OAI22_X1 i_0_131 (.A1(n_0_57), .A2(n_0_15), .B1(n_0_20), .B2(n_0_63), 
      .ZN(n_0_64));
   AOI221_X1 i_0_132 (.A(n_0_46), .B1(n_0_8), .B2(n_0_53), .C1(n_0_64), .C2(
      n_0_38), .ZN(n_0_65));
   INV_X1 i_0_133 (.A(n_0_65), .ZN(n_0_66));
   INV_X1 i_0_134 (.A(n_0_44), .ZN(n_0_67));
   OAI22_X1 i_0_135 (.A1(n_0_44), .A2(n_0_66), .B1(n_0_67), .B2(n_0_65), 
      .ZN(n_0_68));
   INV_X1 i_0_136 (.A(Input1_2_Positive[1]), .ZN(n_0_69));
   OR2_X1 i_0_137 (.A1(n_0_68), .A2(n_0_69), .ZN(n_0_70));
   NAND2_X1 i_0_138 (.A1(n_0_60), .A2(n_0_11), .ZN(n_0_71));
   NOR2_X1 i_0_139 (.A1(n_0_70), .A2(n_0_71), .ZN(n_0_316__0));
   NOR3_X1 i_0_140 (.A1(n_0_45), .A2(n_0_12), .A3(n_0_15), .ZN(n_0_72));
   NAND3_X1 i_0_141 (.A1(n_0_62), .A2(newB[12]), .A3(n_0_22), .ZN(n_0_73));
   NAND2_X1 i_0_142 (.A1(n_0_58), .A2(newB[20]), .ZN(n_0_74));
   OAI211_X1 i_0_143 (.A(n_0_14), .B(n_0_73), .C1(n_0_23), .C2(n_0_74), .ZN(
      n_0_75));
   INV_X1 i_0_144 (.A(newB[28]), .ZN(n_0_76));
   OAI22_X1 i_0_145 (.A1(n_0_31), .A2(n_0_76), .B1(n_0_29), .B2(n_0_54), 
      .ZN(n_0_77));
   INV_X1 i_0_146 (.A(newB[8]), .ZN(n_0_78));
   INV_X1 i_0_147 (.A(newB[4]), .ZN(n_0_79));
   OAI22_X1 i_0_148 (.A1(n_0_78), .A2(n_0_20), .B1(n_0_79), .B2(
      shiftingAmount[2]), .ZN(n_0_80));
   AOI22_X1 i_0_149 (.A1(n_0_55), .A2(n_0_28), .B1(n_0_13), .B2(
      shiftingAmount[4]), .ZN(n_0_81));
   AOI222_X1 i_0_150 (.A1(n_0_77), .A2(shiftingAmount[4]), .B1(n_0_80), .B2(
      n_0_9), .C1(n_0_81), .C2(n_0_34), .ZN(n_0_82));
   OAI22_X1 i_0_151 (.A1(n_0_51), .A2(shiftingAmount[1]), .B1(n_0_82), .B2(
      n_0_38), .ZN(n_0_83));
   AOI211_X1 i_0_152 (.A(n_0_72), .B(n_0_75), .C1(n_0_83), .C2(n_0_8), .ZN(
      n_0_84));
   INV_X1 i_0_153 (.A(n_0_84), .ZN(n_0_85));
   NAND3_X1 i_0_154 (.A1(n_0_67), .A2(n_0_65), .A3(n_0_85), .ZN(n_0_86));
   NAND3_X1 i_0_155 (.A1(n_0_44), .A2(n_0_66), .A3(n_0_84), .ZN(n_0_87));
   AOI21_X1 i_0_156 (.A(n_0_69), .B1(n_0_86), .B2(n_0_87), .ZN(n_0_88));
   NOR2_X1 i_0_157 (.A1(n_0_68), .A2(n_0_84), .ZN(n_0_89));
   NOR2_X1 i_0_158 (.A1(n_0_68), .A2(n_0_85), .ZN(n_0_90));
   AOI221_X1 i_0_159 (.A(n_0_88), .B1(n_0_89), .B2(Input1_1_Negative[1]), 
      .C1(Input1_1_Positive[1]), .C2(n_0_90), .ZN(n_0_91));
   NOR2_X1 i_0_160 (.A1(n_0_91), .A2(n_0_71), .ZN(n_0_318__0));
   INV_X1 i_0_161 (.A(n_0_87), .ZN(n_0_92));
   AOI22_X1 i_0_162 (.A1(n_0_90), .A2(Input1_2_Positive[3]), .B1(
      Input1_1_Positive[1]), .B2(n_0_92), .ZN(n_0_93));
   INV_X1 i_0_163 (.A(n_0_86), .ZN(n_0_94));
   AOI22_X1 i_0_164 (.A1(n_0_89), .A2(Input1_2_Negative[3]), .B1(
      Input1_1_Negative[1]), .B2(n_0_94), .ZN(n_0_95));
   NAND2_X1 i_0_165 (.A1(n_0_93), .A2(n_0_95), .ZN(n_0_96));
   INV_X1 i_0_166 (.A(n_0_96), .ZN(n_0_97));
   NAND2_X1 i_0_167 (.A1(n_0_60), .A2(n_0_22), .ZN(n_0_98));
   OAI22_X1 i_0_168 (.A1(n_0_97), .A2(n_0_71), .B1(n_0_70), .B2(n_0_98), 
      .ZN(n_0_320__0));
   AOI22_X1 i_0_169 (.A1(n_0_90), .A2(Input1_1_Positive[3]), .B1(
      Input1_2_Positive[3]), .B2(n_0_92), .ZN(n_0_99));
   AOI22_X1 i_0_170 (.A1(n_0_89), .A2(Input1_1_Negative[3]), .B1(
      Input1_2_Negative[3]), .B2(n_0_94), .ZN(n_0_100));
   NAND2_X1 i_0_171 (.A1(n_0_99), .A2(n_0_100), .ZN(n_0_101));
   INV_X1 i_0_172 (.A(n_0_101), .ZN(n_0_102));
   OAI22_X1 i_0_173 (.A1(n_0_91), .A2(n_0_98), .B1(n_0_71), .B2(n_0_102), 
      .ZN(n_0_321__0));
   AOI22_X1 i_0_174 (.A1(n_0_90), .A2(Input1_2_Positive[5]), .B1(
      Input1_1_Positive[3]), .B2(n_0_92), .ZN(n_0_103));
   AOI22_X1 i_0_175 (.A1(n_0_89), .A2(Input1_2_Negative[5]), .B1(
      Input1_1_Negative[3]), .B2(n_0_94), .ZN(n_0_104));
   NAND2_X1 i_0_176 (.A1(n_0_103), .A2(n_0_104), .ZN(n_0_105));
   INV_X1 i_0_177 (.A(n_0_60), .ZN(n_0_106));
   NOR2_X1 i_0_178 (.A1(n_0_106), .A2(shiftingAmount[2]), .ZN(n_0_107));
   INV_X1 i_0_179 (.A(n_0_70), .ZN(n_0_108));
   NOR2_X1 i_0_180 (.A1(shiftingAmount[4]), .A2(shiftingAmount[5]), .ZN(n_0_109));
   AND2_X1 i_0_181 (.A1(n_0_30), .A2(n_0_109), .ZN(n_0_110));
   AOI22_X1 i_0_182 (.A1(n_0_105), .A2(n_0_107), .B1(n_0_108), .B2(n_0_110), 
      .ZN(n_0_111));
   OAI22_X1 i_0_183 (.A1(n_0_111), .A2(shiftingAmount[1]), .B1(n_0_97), .B2(
      n_0_98), .ZN(n_0_322__0));
   INV_X1 i_0_184 (.A(n_0_91), .ZN(n_0_112));
   AOI22_X1 i_0_185 (.A1(n_0_89), .A2(Input1_1_Negative[5]), .B1(
      Input1_2_Positive[5]), .B2(n_0_92), .ZN(n_0_113));
   AOI22_X1 i_0_186 (.A1(n_0_90), .A2(Input1_1_Positive[5]), .B1(
      Input1_2_Negative[5]), .B2(n_0_94), .ZN(n_0_114));
   NAND2_X1 i_0_187 (.A1(n_0_113), .A2(n_0_114), .ZN(n_0_115));
   AOI22_X1 i_0_188 (.A1(n_0_112), .A2(n_0_110), .B1(n_0_107), .B2(n_0_115), 
      .ZN(n_0_116));
   OAI22_X1 i_0_189 (.A1(n_0_116), .A2(shiftingAmount[1]), .B1(n_0_102), 
      .B2(n_0_98), .ZN(n_0_323__0));
   AOI22_X1 i_0_190 (.A1(n_0_89), .A2(Input1_2_Negative[7]), .B1(
      Input1_1_Positive[5]), .B2(n_0_92), .ZN(n_0_117));
   AOI22_X1 i_0_191 (.A1(n_0_90), .A2(Input1_2_Positive[7]), .B1(
      Input1_1_Negative[5]), .B2(n_0_94), .ZN(n_0_118));
   NAND2_X1 i_0_192 (.A1(n_0_117), .A2(n_0_118), .ZN(n_0_119));
   INV_X1 i_0_193 (.A(n_0_119), .ZN(n_0_120));
   NOR2_X1 i_0_194 (.A1(n_0_120), .A2(n_0_106), .ZN(n_0_121));
   AOI22_X1 i_0_195 (.A1(n_0_121), .A2(n_0_20), .B1(n_0_96), .B2(n_0_110), 
      .ZN(n_0_122));
   OAI22_X1 i_0_196 (.A1(n_0_122), .A2(shiftingAmount[1]), .B1(n_0_38), .B2(
      n_0_111), .ZN(n_0_324__0));
   AOI22_X1 i_0_197 (.A1(n_0_90), .A2(Input1_1_Positive[7]), .B1(
      Input1_2_Positive[7]), .B2(n_0_92), .ZN(n_0_123));
   AOI22_X1 i_0_198 (.A1(n_0_89), .A2(Input1_1_Negative[7]), .B1(
      Input1_2_Negative[7]), .B2(n_0_94), .ZN(n_0_124));
   NAND2_X1 i_0_199 (.A1(n_0_123), .A2(n_0_124), .ZN(n_0_125));
   AOI22_X1 i_0_200 (.A1(n_0_125), .A2(n_0_107), .B1(n_0_101), .B2(n_0_110), 
      .ZN(n_0_126));
   OAI22_X1 i_0_201 (.A1(n_0_116), .A2(n_0_38), .B1(shiftingAmount[1]), .B2(
      n_0_126), .ZN(n_0_325__0));
   AOI22_X1 i_0_202 (.A1(n_0_90), .A2(Input1_2_Positive[9]), .B1(
      Input1_1_Positive[7]), .B2(n_0_92), .ZN(n_0_127));
   AOI22_X1 i_0_203 (.A1(n_0_89), .A2(Input1_2_Negative[9]), .B1(
      Input1_1_Negative[7]), .B2(n_0_94), .ZN(n_0_128));
   NAND2_X1 i_0_204 (.A1(n_0_127), .A2(n_0_128), .ZN(n_0_129));
   INV_X1 i_0_205 (.A(n_0_129), .ZN(n_0_130));
   INV_X1 i_0_206 (.A(n_0_62), .ZN(n_0_131));
   OAI22_X1 i_0_207 (.A1(n_0_130), .A2(n_0_106), .B1(n_0_131), .B2(n_0_70), 
      .ZN(n_0_132));
   AOI22_X1 i_0_208 (.A1(n_0_132), .A2(n_0_20), .B1(n_0_105), .B2(n_0_110), 
      .ZN(n_0_133));
   OAI22_X1 i_0_209 (.A1(n_0_133), .A2(shiftingAmount[1]), .B1(n_0_122), 
      .B2(n_0_38), .ZN(n_0_326__0));
   AOI22_X1 i_0_210 (.A1(n_0_90), .A2(Input1_1_Positive[9]), .B1(
      Input1_2_Positive[9]), .B2(n_0_92), .ZN(n_0_134));
   AOI22_X1 i_0_211 (.A1(n_0_89), .A2(Input1_1_Negative[9]), .B1(
      Input1_2_Negative[9]), .B2(n_0_94), .ZN(n_0_135));
   NAND2_X1 i_0_212 (.A1(n_0_134), .A2(n_0_135), .ZN(n_0_136));
   INV_X1 i_0_213 (.A(n_0_136), .ZN(n_0_137));
   OAI22_X1 i_0_214 (.A1(n_0_91), .A2(n_0_131), .B1(n_0_137), .B2(n_0_106), 
      .ZN(n_0_138));
   AOI22_X1 i_0_215 (.A1(n_0_138), .A2(n_0_20), .B1(n_0_110), .B2(n_0_115), 
      .ZN(n_0_139));
   OAI22_X1 i_0_216 (.A1(n_0_139), .A2(shiftingAmount[1]), .B1(n_0_38), .B2(
      n_0_126), .ZN(n_0_327__0));
   AOI22_X1 i_0_217 (.A1(n_0_89), .A2(Input1_2_Negative[11]), .B1(
      Input1_1_Positive[9]), .B2(n_0_92), .ZN(n_0_140));
   AOI22_X1 i_0_218 (.A1(n_0_90), .A2(Input1_2_Positive[11]), .B1(
      Input1_1_Negative[9]), .B2(n_0_94), .ZN(n_0_141));
   NAND2_X1 i_0_219 (.A1(n_0_140), .A2(n_0_141), .ZN(n_0_142));
   INV_X1 i_0_220 (.A(n_0_142), .ZN(n_0_143));
   OAI22_X1 i_0_221 (.A1(n_0_97), .A2(n_0_131), .B1(n_0_143), .B2(n_0_106), 
      .ZN(n_0_144));
   AOI22_X1 i_0_222 (.A1(n_0_144), .A2(n_0_20), .B1(n_0_121), .B2(
      shiftingAmount[2]), .ZN(n_0_145));
   OAI22_X1 i_0_223 (.A1(n_0_145), .A2(shiftingAmount[1]), .B1(n_0_133), 
      .B2(n_0_38), .ZN(n_0_328__0));
   AOI22_X1 i_0_224 (.A1(n_0_89), .A2(Input1_1_Negative[11]), .B1(n_0_92), 
      .B2(Input1_2_Positive[11]), .ZN(n_0_146));
   AOI22_X1 i_0_225 (.A1(n_0_90), .A2(Input1_1_Positive[11]), .B1(
      Input1_2_Negative[11]), .B2(n_0_94), .ZN(n_0_147));
   NAND2_X1 i_0_226 (.A1(n_0_146), .A2(n_0_147), .ZN(n_0_148));
   INV_X1 i_0_227 (.A(n_0_148), .ZN(n_0_149));
   OAI22_X1 i_0_228 (.A1(n_0_149), .A2(n_0_106), .B1(n_0_102), .B2(n_0_131), 
      .ZN(n_0_150));
   AOI22_X1 i_0_229 (.A1(n_0_150), .A2(n_0_20), .B1(n_0_125), .B2(n_0_110), 
      .ZN(n_0_151));
   OAI22_X1 i_0_230 (.A1(n_0_139), .A2(n_0_38), .B1(n_0_151), .B2(
      shiftingAmount[1]), .ZN(n_0_329__0));
   INV_X1 i_0_231 (.A(n_0_105), .ZN(n_0_152));
   AOI22_X1 i_0_232 (.A1(n_0_89), .A2(Input1_2_Negative[13]), .B1(
      Input1_1_Positive[11]), .B2(n_0_92), .ZN(n_0_153));
   AOI22_X1 i_0_233 (.A1(n_0_90), .A2(Input1_2_Positive[13]), .B1(
      Input1_1_Negative[11]), .B2(n_0_94), .ZN(n_0_154));
   NAND2_X1 i_0_234 (.A1(n_0_153), .A2(n_0_154), .ZN(n_0_155));
   INV_X1 i_0_235 (.A(n_0_155), .ZN(n_0_156));
   OAI22_X1 i_0_236 (.A1(n_0_152), .A2(n_0_131), .B1(n_0_156), .B2(n_0_106), 
      .ZN(n_0_157));
   AOI22_X1 i_0_237 (.A1(n_0_157), .A2(n_0_20), .B1(n_0_132), .B2(
      shiftingAmount[2]), .ZN(n_0_158));
   OAI22_X1 i_0_238 (.A1(n_0_158), .A2(shiftingAmount[1]), .B1(n_0_145), 
      .B2(n_0_38), .ZN(n_0_330__0));
   AOI22_X1 i_0_239 (.A1(n_0_90), .A2(Input1_1_Positive[13]), .B1(n_0_92), 
      .B2(Input1_2_Positive[13]), .ZN(n_0_159));
   AOI22_X1 i_0_240 (.A1(n_0_89), .A2(Input1_1_Negative[13]), .B1(
      Input1_2_Negative[13]), .B2(n_0_94), .ZN(n_0_160));
   NAND2_X1 i_0_241 (.A1(n_0_159), .A2(n_0_160), .ZN(n_0_161));
   INV_X1 i_0_242 (.A(n_0_161), .ZN(n_0_162));
   INV_X1 i_0_243 (.A(n_0_115), .ZN(n_0_163));
   OAI22_X1 i_0_244 (.A1(n_0_162), .A2(n_0_106), .B1(n_0_163), .B2(n_0_131), 
      .ZN(n_0_164));
   AOI22_X1 i_0_245 (.A1(n_0_138), .A2(shiftingAmount[2]), .B1(n_0_164), 
      .B2(n_0_20), .ZN(n_0_165));
   OAI22_X1 i_0_246 (.A1(n_0_165), .A2(shiftingAmount[1]), .B1(n_0_151), 
      .B2(n_0_38), .ZN(n_0_331__0));
   AOI22_X1 i_0_247 (.A1(n_0_89), .A2(Input1_2_Negative[15]), .B1(
      Input1_1_Negative[13]), .B2(n_0_94), .ZN(n_0_166));
   AOI22_X1 i_0_248 (.A1(n_0_90), .A2(Input1_2_Positive[15]), .B1(
      Input1_1_Positive[13]), .B2(n_0_92), .ZN(n_0_167));
   NAND2_X1 i_0_249 (.A1(n_0_166), .A2(n_0_167), .ZN(n_0_168));
   INV_X1 i_0_250 (.A(n_0_168), .ZN(n_0_169));
   OAI22_X1 i_0_251 (.A1(n_0_120), .A2(n_0_131), .B1(n_0_169), .B2(n_0_106), 
      .ZN(n_0_170));
   AOI22_X1 i_0_252 (.A1(n_0_144), .A2(shiftingAmount[2]), .B1(n_0_170), 
      .B2(n_0_20), .ZN(n_0_171));
   OAI22_X1 i_0_253 (.A1(n_0_171), .A2(shiftingAmount[1]), .B1(n_0_158), 
      .B2(n_0_38), .ZN(n_0_332__0));
   INV_X1 i_0_254 (.A(n_0_125), .ZN(n_0_172));
   AOI22_X1 i_0_255 (.A1(n_0_89), .A2(Input1_1_Negative[15]), .B1(
      Input1_2_Negative[15]), .B2(n_0_94), .ZN(n_0_173));
   AOI22_X1 i_0_256 (.A1(n_0_90), .A2(Input1_1_Positive[15]), .B1(
      Input1_2_Positive[15]), .B2(n_0_92), .ZN(n_0_174));
   NAND2_X1 i_0_257 (.A1(n_0_173), .A2(n_0_174), .ZN(n_0_175));
   INV_X1 i_0_258 (.A(n_0_175), .ZN(n_0_176));
   OAI22_X1 i_0_259 (.A1(n_0_172), .A2(n_0_131), .B1(n_0_176), .B2(n_0_106), 
      .ZN(n_0_177));
   AOI22_X1 i_0_260 (.A1(n_0_177), .A2(n_0_20), .B1(n_0_150), .B2(
      shiftingAmount[2]), .ZN(n_0_178));
   OAI22_X1 i_0_261 (.A1(n_0_165), .A2(n_0_38), .B1(n_0_178), .B2(
      shiftingAmount[1]), .ZN(n_0_333__0));
   AOI22_X1 i_0_262 (.A1(n_0_89), .A2(Input1_2_Negative[17]), .B1(
      Input1_1_Negative[15]), .B2(n_0_94), .ZN(n_0_179));
   AOI22_X1 i_0_263 (.A1(n_0_90), .A2(Input1_2_Positive[17]), .B1(
      Input1_1_Positive[15]), .B2(n_0_92), .ZN(n_0_180));
   NAND2_X1 i_0_264 (.A1(n_0_179), .A2(n_0_180), .ZN(n_0_181));
   AOI22_X1 i_0_265 (.A1(n_0_181), .A2(n_0_109), .B1(n_0_16), .B2(n_0_108), 
      .ZN(n_0_182));
   OAI22_X1 i_0_266 (.A1(n_0_182), .A2(shiftingAmount[3]), .B1(n_0_131), 
      .B2(n_0_130), .ZN(n_0_183));
   AOI22_X1 i_0_267 (.A1(n_0_183), .A2(n_0_20), .B1(shiftingAmount[2]), .B2(
      n_0_157), .ZN(n_0_184));
   OAI22_X1 i_0_268 (.A1(n_0_184), .A2(shiftingAmount[1]), .B1(n_0_171), 
      .B2(n_0_38), .ZN(n_0_334__0));
   AOI22_X1 i_0_269 (.A1(n_0_89), .A2(Input1_1_Negative[17]), .B1(
      Input1_2_Negative[17]), .B2(n_0_94), .ZN(n_0_185));
   AOI22_X1 i_0_270 (.A1(n_0_90), .A2(Input1_1_Positive[17]), .B1(
      Input1_2_Positive[17]), .B2(n_0_92), .ZN(n_0_186));
   NAND2_X1 i_0_271 (.A1(n_0_185), .A2(n_0_186), .ZN(n_0_187));
   OAI22_X1 i_0_272 (.A1(n_0_112), .A2(n_0_28), .B1(n_0_187), .B2(
      shiftingAmount[4]), .ZN(n_0_188));
   OAI22_X1 i_0_273 (.A1(n_0_188), .A2(n_0_59), .B1(n_0_131), .B2(n_0_137), 
      .ZN(n_0_189));
   AOI22_X1 i_0_274 (.A1(n_0_189), .A2(n_0_20), .B1(shiftingAmount[2]), .B2(
      n_0_164), .ZN(n_0_190));
   OAI22_X1 i_0_275 (.A1(n_0_190), .A2(shiftingAmount[1]), .B1(n_0_38), .B2(
      n_0_178), .ZN(n_0_335__0));
   AOI22_X1 i_0_276 (.A1(n_0_89), .A2(Input1_2_Negative[19]), .B1(
      Input1_1_Negative[17]), .B2(n_0_94), .ZN(n_0_191));
   AOI22_X1 i_0_277 (.A1(n_0_90), .A2(Input1_2_Positive[19]), .B1(
      Input1_1_Positive[17]), .B2(n_0_92), .ZN(n_0_192));
   NAND2_X1 i_0_278 (.A1(n_0_191), .A2(n_0_192), .ZN(n_0_193));
   OAI22_X1 i_0_279 (.A1(n_0_96), .A2(n_0_28), .B1(n_0_193), .B2(
      shiftingAmount[4]), .ZN(n_0_194));
   OAI22_X1 i_0_280 (.A1(n_0_194), .A2(n_0_59), .B1(n_0_131), .B2(n_0_143), 
      .ZN(n_0_195));
   AOI22_X1 i_0_281 (.A1(n_0_195), .A2(n_0_20), .B1(shiftingAmount[2]), .B2(
      n_0_170), .ZN(n_0_196));
   OAI22_X1 i_0_282 (.A1(n_0_196), .A2(shiftingAmount[1]), .B1(n_0_184), 
      .B2(n_0_38), .ZN(n_0_336__0));
   AOI22_X1 i_0_283 (.A1(n_0_89), .A2(Input1_1_Negative[19]), .B1(
      Input1_2_Positive[19]), .B2(n_0_92), .ZN(n_0_197));
   AOI22_X1 i_0_284 (.A1(n_0_90), .A2(Input1_1_Positive[19]), .B1(
      Input1_2_Negative[19]), .B2(n_0_94), .ZN(n_0_198));
   NAND2_X1 i_0_285 (.A1(n_0_197), .A2(n_0_198), .ZN(n_0_199));
   OAI22_X1 i_0_286 (.A1(n_0_101), .A2(n_0_28), .B1(n_0_199), .B2(
      shiftingAmount[4]), .ZN(n_0_200));
   OAI22_X1 i_0_287 (.A1(n_0_200), .A2(n_0_59), .B1(n_0_131), .B2(n_0_149), 
      .ZN(n_0_201));
   AOI22_X1 i_0_288 (.A1(n_0_201), .A2(n_0_20), .B1(shiftingAmount[2]), .B2(
      n_0_177), .ZN(n_0_202));
   OAI22_X1 i_0_289 (.A1(n_0_190), .A2(n_0_38), .B1(shiftingAmount[1]), .B2(
      n_0_202), .ZN(n_0_337__0));
   AOI22_X1 i_0_290 (.A1(n_0_89), .A2(Input1_2_Negative[21]), .B1(
      Input1_1_Negative[19]), .B2(n_0_94), .ZN(n_0_203));
   AOI22_X1 i_0_291 (.A1(n_0_90), .A2(Input1_2_Positive[21]), .B1(
      Input1_1_Positive[19]), .B2(n_0_92), .ZN(n_0_204));
   NAND2_X1 i_0_292 (.A1(n_0_203), .A2(n_0_204), .ZN(n_0_205));
   AOI22_X1 i_0_293 (.A1(n_0_205), .A2(n_0_109), .B1(n_0_105), .B2(n_0_16), 
      .ZN(n_0_206));
   OAI22_X1 i_0_294 (.A1(n_0_206), .A2(shiftingAmount[3]), .B1(n_0_131), 
      .B2(n_0_156), .ZN(n_0_207));
   AOI22_X1 i_0_295 (.A1(n_0_207), .A2(n_0_20), .B1(n_0_183), .B2(
      shiftingAmount[2]), .ZN(n_0_208));
   OAI22_X1 i_0_296 (.A1(n_0_208), .A2(shiftingAmount[1]), .B1(n_0_196), 
      .B2(n_0_38), .ZN(n_0_338__0));
   AOI22_X1 i_0_297 (.A1(n_0_89), .A2(Input1_1_Negative[21]), .B1(
      Input1_2_Negative[21]), .B2(n_0_94), .ZN(n_0_209));
   AOI22_X1 i_0_298 (.A1(n_0_90), .A2(Input1_1_Positive[21]), .B1(
      Input1_2_Positive[21]), .B2(n_0_92), .ZN(n_0_210));
   NAND2_X1 i_0_299 (.A1(n_0_209), .A2(n_0_210), .ZN(n_0_211));
   AOI22_X1 i_0_300 (.A1(n_0_115), .A2(n_0_16), .B1(n_0_211), .B2(n_0_109), 
      .ZN(n_0_212));
   OAI22_X1 i_0_301 (.A1(n_0_212), .A2(shiftingAmount[3]), .B1(n_0_131), 
      .B2(n_0_162), .ZN(n_0_213));
   AOI22_X1 i_0_302 (.A1(n_0_189), .A2(shiftingAmount[2]), .B1(n_0_213), 
      .B2(n_0_20), .ZN(n_0_214));
   OAI22_X1 i_0_303 (.A1(n_0_214), .A2(shiftingAmount[1]), .B1(n_0_38), .B2(
      n_0_202), .ZN(n_0_339__0));
   AOI22_X1 i_0_304 (.A1(n_0_89), .A2(Input1_2_Negative[23]), .B1(
      Input1_1_Positive[21]), .B2(n_0_92), .ZN(n_0_215));
   AOI22_X1 i_0_305 (.A1(n_0_90), .A2(Input1_2_Positive[23]), .B1(
      Input1_1_Negative[21]), .B2(n_0_94), .ZN(n_0_216));
   NAND2_X1 i_0_306 (.A1(n_0_215), .A2(n_0_216), .ZN(n_0_217));
   OAI22_X1 i_0_307 (.A1(n_0_119), .A2(n_0_28), .B1(n_0_217), .B2(
      shiftingAmount[4]), .ZN(n_0_218));
   OAI22_X1 i_0_308 (.A1(n_0_218), .A2(n_0_59), .B1(n_0_131), .B2(n_0_169), 
      .ZN(n_0_219));
   AOI22_X1 i_0_309 (.A1(n_0_195), .A2(shiftingAmount[2]), .B1(n_0_219), 
      .B2(n_0_20), .ZN(n_0_220));
   OAI22_X1 i_0_310 (.A1(n_0_220), .A2(shiftingAmount[1]), .B1(n_0_208), 
      .B2(n_0_38), .ZN(n_0_340__0));
   AOI22_X1 i_0_311 (.A1(n_0_89), .A2(Input1_1_Negative[23]), .B1(
      Input1_2_Positive[23]), .B2(n_0_92), .ZN(n_0_221));
   AOI22_X1 i_0_312 (.A1(n_0_90), .A2(Input1_1_Positive[23]), .B1(
      Input1_2_Negative[23]), .B2(n_0_94), .ZN(n_0_222));
   NAND2_X1 i_0_313 (.A1(n_0_221), .A2(n_0_222), .ZN(n_0_223));
   OAI22_X1 i_0_314 (.A1(n_0_125), .A2(n_0_28), .B1(n_0_223), .B2(
      shiftingAmount[4]), .ZN(n_0_224));
   OAI22_X1 i_0_315 (.A1(n_0_224), .A2(n_0_59), .B1(n_0_131), .B2(n_0_176), 
      .ZN(n_0_225));
   AOI22_X1 i_0_316 (.A1(n_0_201), .A2(shiftingAmount[2]), .B1(n_0_225), 
      .B2(n_0_20), .ZN(n_0_226));
   OAI22_X1 i_0_317 (.A1(n_0_214), .A2(n_0_38), .B1(n_0_226), .B2(
      shiftingAmount[1]), .ZN(n_0_341__0));
   AOI22_X1 i_0_318 (.A1(n_0_90), .A2(Input1_2_Positive[25]), .B1(n_0_92), 
      .B2(Input1_1_Positive[23]), .ZN(n_0_227));
   AOI22_X1 i_0_319 (.A1(n_0_89), .A2(Input1_2_Negative[25]), .B1(
      Input1_1_Negative[23]), .B2(n_0_94), .ZN(n_0_228));
   NAND2_X1 i_0_320 (.A1(n_0_227), .A2(n_0_228), .ZN(n_0_229));
   AOI22_X1 i_0_321 (.A1(n_0_229), .A2(n_0_109), .B1(n_0_129), .B2(n_0_16), 
      .ZN(n_0_230));
   OAI22_X1 i_0_322 (.A1(n_0_230), .A2(shiftingAmount[3]), .B1(n_0_182), 
      .B2(n_0_17), .ZN(n_0_231));
   AOI22_X1 i_0_323 (.A1(n_0_231), .A2(n_0_20), .B1(n_0_207), .B2(
      shiftingAmount[2]), .ZN(n_0_232));
   OAI22_X1 i_0_324 (.A1(n_0_232), .A2(shiftingAmount[1]), .B1(n_0_220), 
      .B2(n_0_38), .ZN(n_0_342__0));
   AOI22_X1 i_0_325 (.A1(n_0_90), .A2(Input1_1_Positive[25]), .B1(n_0_92), 
      .B2(Input1_2_Positive[25]), .ZN(n_0_233));
   AOI22_X1 i_0_326 (.A1(n_0_89), .A2(Input1_1_Negative[25]), .B1(
      Input1_2_Negative[25]), .B2(n_0_94), .ZN(n_0_234));
   NAND2_X1 i_0_327 (.A1(n_0_233), .A2(n_0_234), .ZN(n_0_235));
   AOI22_X1 i_0_328 (.A1(n_0_235), .A2(n_0_109), .B1(n_0_136), .B2(n_0_16), 
      .ZN(n_0_236));
   OAI22_X1 i_0_329 (.A1(n_0_188), .A2(n_0_61), .B1(shiftingAmount[3]), .B2(
      n_0_236), .ZN(n_0_237));
   AOI22_X1 i_0_330 (.A1(n_0_237), .A2(n_0_20), .B1(n_0_213), .B2(
      shiftingAmount[2]), .ZN(n_0_238));
   OAI22_X1 i_0_331 (.A1(n_0_238), .A2(shiftingAmount[1]), .B1(n_0_226), 
      .B2(n_0_38), .ZN(n_0_343__0));
   AOI22_X1 i_0_332 (.A1(n_0_89), .A2(Input1_2_Negative[27]), .B1(
      Input1_1_Negative[25]), .B2(n_0_94), .ZN(n_0_239));
   AOI22_X1 i_0_333 (.A1(n_0_90), .A2(Input1_2_Positive[27]), .B1(
      Input1_1_Positive[25]), .B2(n_0_92), .ZN(n_0_240));
   NAND2_X1 i_0_334 (.A1(n_0_239), .A2(n_0_240), .ZN(n_0_241));
   AOI22_X1 i_0_335 (.A1(n_0_142), .A2(n_0_16), .B1(n_0_241), .B2(n_0_109), 
      .ZN(n_0_242));
   OAI22_X1 i_0_336 (.A1(n_0_242), .A2(shiftingAmount[3]), .B1(n_0_194), 
      .B2(n_0_61), .ZN(n_0_243));
   AOI22_X1 i_0_337 (.A1(n_0_243), .A2(n_0_20), .B1(n_0_219), .B2(
      shiftingAmount[2]), .ZN(n_0_244));
   OAI22_X1 i_0_338 (.A1(n_0_244), .A2(shiftingAmount[1]), .B1(n_0_232), 
      .B2(n_0_38), .ZN(n_0_344__0));
   AOI22_X1 i_0_339 (.A1(n_0_89), .A2(Input1_1_Negative[27]), .B1(
      Input1_2_Negative[27]), .B2(n_0_94), .ZN(n_0_245));
   AOI22_X1 i_0_340 (.A1(n_0_90), .A2(Input1_1_Positive[27]), .B1(
      Input1_2_Positive[27]), .B2(n_0_92), .ZN(n_0_246));
   NAND2_X1 i_0_341 (.A1(n_0_245), .A2(n_0_246), .ZN(n_0_247));
   AOI22_X1 i_0_342 (.A1(n_0_148), .A2(n_0_16), .B1(n_0_247), .B2(n_0_109), 
      .ZN(n_0_248));
   OAI22_X1 i_0_343 (.A1(n_0_248), .A2(shiftingAmount[3]), .B1(n_0_200), 
      .B2(n_0_61), .ZN(n_0_249));
   AOI22_X1 i_0_344 (.A1(n_0_249), .A2(n_0_20), .B1(n_0_225), .B2(
      shiftingAmount[2]), .ZN(n_0_250));
   OAI22_X1 i_0_345 (.A1(n_0_238), .A2(n_0_38), .B1(n_0_250), .B2(
      shiftingAmount[1]), .ZN(n_0_345__0));
   AOI22_X1 i_0_346 (.A1(n_0_90), .A2(Input1_2_Positive[29]), .B1(n_0_94), 
      .B2(Input1_1_Negative[27]), .ZN(n_0_251));
   AOI22_X1 i_0_347 (.A1(n_0_89), .A2(Input1_2_Negative[29]), .B1(
      Input1_1_Positive[27]), .B2(n_0_92), .ZN(n_0_252));
   NAND2_X1 i_0_348 (.A1(n_0_251), .A2(n_0_252), .ZN(n_0_253));
   AOI22_X1 i_0_349 (.A1(n_0_253), .A2(n_0_109), .B1(n_0_155), .B2(n_0_16), 
      .ZN(n_0_254));
   OAI22_X1 i_0_350 (.A1(n_0_254), .A2(shiftingAmount[3]), .B1(n_0_206), 
      .B2(n_0_17), .ZN(n_0_255));
   AOI22_X1 i_0_351 (.A1(n_0_255), .A2(n_0_20), .B1(n_0_231), .B2(
      shiftingAmount[2]), .ZN(n_0_256));
   OAI22_X1 i_0_352 (.A1(n_0_256), .A2(shiftingAmount[1]), .B1(n_0_244), 
      .B2(n_0_38), .ZN(n_0_346__0));
   AOI22_X1 i_0_353 (.A1(n_0_90), .A2(Input1_1_Positive[29]), .B1(
      Input1_2_Positive[29]), .B2(n_0_92), .ZN(n_0_257));
   AOI22_X1 i_0_354 (.A1(n_0_89), .A2(Input1_1_Negative[29]), .B1(
      Input1_2_Negative[29]), .B2(n_0_94), .ZN(n_0_258));
   NAND2_X1 i_0_355 (.A1(n_0_257), .A2(n_0_258), .ZN(n_0_259));
   AOI22_X1 i_0_356 (.A1(n_0_161), .A2(n_0_16), .B1(n_0_259), .B2(n_0_109), 
      .ZN(n_0_260));
   OAI22_X1 i_0_357 (.A1(n_0_260), .A2(shiftingAmount[3]), .B1(n_0_212), 
      .B2(n_0_17), .ZN(n_0_261));
   AOI22_X1 i_0_358 (.A1(n_0_237), .A2(shiftingAmount[2]), .B1(n_0_261), 
      .B2(n_0_20), .ZN(n_0_262));
   OAI22_X1 i_0_359 (.A1(n_0_262), .A2(shiftingAmount[1]), .B1(n_0_250), 
      .B2(n_0_38), .ZN(n_0_347__0));
   AOI22_X1 i_0_360 (.A1(n_0_89), .A2(Input1_2_Negative[31]), .B1(
      Input1_1_Negative[29]), .B2(n_0_94), .ZN(n_0_263));
   AOI22_X1 i_0_361 (.A1(n_0_90), .A2(Input1_2_Positive[31]), .B1(
      Input1_1_Positive[29]), .B2(n_0_92), .ZN(n_0_264));
   NAND2_X1 i_0_362 (.A1(n_0_263), .A2(n_0_264), .ZN(n_0_265));
   AOI22_X1 i_0_363 (.A1(n_0_265), .A2(n_0_109), .B1(n_0_168), .B2(n_0_16), 
      .ZN(n_0_266));
   OAI22_X1 i_0_364 (.A1(n_0_266), .A2(shiftingAmount[3]), .B1(n_0_218), 
      .B2(n_0_61), .ZN(n_0_267));
   AOI22_X1 i_0_365 (.A1(n_0_243), .A2(shiftingAmount[2]), .B1(n_0_267), 
      .B2(n_0_20), .ZN(n_0_268));
   OAI22_X1 i_0_366 (.A1(n_0_268), .A2(shiftingAmount[1]), .B1(n_0_256), 
      .B2(n_0_38), .ZN(n_0_348__0));
   AOI22_X1 i_0_367 (.A1(n_0_89), .A2(Input1_1_Negative[63]), .B1(n_0_90), 
      .B2(Input1_1_Positive[63]), .ZN(n_0_269));
   AOI22_X1 i_0_368 (.A1(n_0_92), .A2(Input1_2_Positive[31]), .B1(n_0_94), 
      .B2(Input1_2_Negative[31]), .ZN(n_0_270));
   NAND2_X1 i_0_369 (.A1(n_0_269), .A2(n_0_270), .ZN(n_0_271));
   AOI22_X1 i_0_370 (.A1(n_0_271), .A2(n_0_109), .B1(n_0_175), .B2(n_0_16), 
      .ZN(n_0_272));
   OAI22_X1 i_0_371 (.A1(n_0_272), .A2(shiftingAmount[3]), .B1(n_0_224), 
      .B2(n_0_61), .ZN(n_0_273));
   AOI22_X1 i_0_372 (.A1(n_0_249), .A2(shiftingAmount[2]), .B1(n_0_273), 
      .B2(n_0_20), .ZN(n_0_274));
   OAI22_X1 i_0_373 (.A1(n_0_262), .A2(n_0_38), .B1(n_0_274), .B2(
      shiftingAmount[1]), .ZN(n_0_349__0));
   AOI22_X1 i_0_374 (.A1(n_0_92), .A2(Input1_1_Positive[63]), .B1(n_0_94), 
      .B2(Input1_1_Negative[63]), .ZN(n_0_275));
   NAND2_X1 i_0_375 (.A1(n_0_269), .A2(n_0_275), .ZN(n_0_276));
   NAND2_X1 i_0_376 (.A1(n_0_276), .A2(n_0_109), .ZN(n_0_277));
   INV_X1 i_0_377 (.A(n_0_277), .ZN(n_0_278));
   AOI221_X1 i_0_378 (.A(n_0_278), .B1(shiftingAmount[5]), .B2(n_0_108), 
      .C1(n_0_16), .C2(n_0_181), .ZN(n_0_279));
   OAI22_X1 i_0_379 (.A1(n_0_279), .A2(shiftingAmount[3]), .B1(n_0_17), .B2(
      n_0_230), .ZN(n_0_280));
   AOI22_X1 i_0_380 (.A1(n_0_280), .A2(n_0_20), .B1(shiftingAmount[2]), .B2(
      n_0_255), .ZN(n_0_281));
   OAI22_X1 i_0_381 (.A1(n_0_281), .A2(shiftingAmount[1]), .B1(n_0_38), .B2(
      n_0_268), .ZN(n_0_350__0));
   AOI221_X1 i_0_382 (.A(n_0_278), .B1(n_0_16), .B2(n_0_187), .C1(n_0_112), 
      .C2(shiftingAmount[5]), .ZN(n_0_282));
   OAI22_X1 i_0_383 (.A1(n_0_282), .A2(shiftingAmount[3]), .B1(n_0_17), .B2(
      n_0_236), .ZN(n_0_283));
   AOI22_X1 i_0_384 (.A1(n_0_283), .A2(n_0_20), .B1(shiftingAmount[2]), .B2(
      n_0_261), .ZN(n_0_284));
   OAI22_X1 i_0_385 (.A1(n_0_284), .A2(shiftingAmount[1]), .B1(n_0_38), .B2(
      n_0_274), .ZN(n_0_351__0));
   OAI21_X1 i_0_386 (.A(n_0_277), .B1(n_0_8), .B2(n_0_97), .ZN(n_0_285));
   AOI21_X1 i_0_387 (.A(n_0_285), .B1(n_0_16), .B2(n_0_193), .ZN(n_0_286));
   OAI22_X1 i_0_388 (.A1(n_0_286), .A2(shiftingAmount[3]), .B1(n_0_17), .B2(
      n_0_242), .ZN(n_0_287));
   AOI22_X1 i_0_389 (.A1(n_0_287), .A2(n_0_20), .B1(shiftingAmount[2]), .B2(
      n_0_267), .ZN(n_0_288));
   OAI22_X1 i_0_390 (.A1(n_0_281), .A2(n_0_38), .B1(n_0_288), .B2(
      shiftingAmount[1]), .ZN(n_0_352__0));
   OAI21_X1 i_0_391 (.A(n_0_277), .B1(n_0_8), .B2(n_0_102), .ZN(n_0_289));
   AOI21_X1 i_0_392 (.A(n_0_289), .B1(n_0_16), .B2(n_0_199), .ZN(n_0_290));
   OAI22_X1 i_0_393 (.A1(n_0_290), .A2(shiftingAmount[3]), .B1(n_0_17), .B2(
      n_0_248), .ZN(n_0_291));
   AOI22_X1 i_0_394 (.A1(n_0_291), .A2(n_0_20), .B1(shiftingAmount[2]), .B2(
      n_0_273), .ZN(n_0_292));
   OAI22_X1 i_0_395 (.A1(n_0_284), .A2(n_0_38), .B1(shiftingAmount[1]), .B2(
      n_0_292), .ZN(n_0_353__0));
   AOI221_X1 i_0_396 (.A(n_0_278), .B1(n_0_16), .B2(n_0_205), .C1(
      shiftingAmount[5]), .C2(n_0_105), .ZN(n_0_293));
   OAI22_X1 i_0_397 (.A1(n_0_293), .A2(shiftingAmount[3]), .B1(n_0_17), .B2(
      n_0_254), .ZN(n_0_294));
   AOI22_X1 i_0_398 (.A1(n_0_280), .A2(shiftingAmount[2]), .B1(n_0_294), 
      .B2(n_0_20), .ZN(n_0_295));
   OAI22_X1 i_0_399 (.A1(n_0_295), .A2(shiftingAmount[1]), .B1(n_0_38), .B2(
      n_0_288), .ZN(n_0_354__0));
   AOI221_X1 i_0_400 (.A(n_0_278), .B1(n_0_16), .B2(n_0_211), .C1(
      shiftingAmount[5]), .C2(n_0_115), .ZN(n_0_296));
   OAI22_X1 i_0_401 (.A1(n_0_296), .A2(shiftingAmount[3]), .B1(n_0_17), .B2(
      n_0_260), .ZN(n_0_297));
   AOI22_X1 i_0_402 (.A1(n_0_283), .A2(shiftingAmount[2]), .B1(n_0_297), 
      .B2(n_0_20), .ZN(n_0_298));
   OAI22_X1 i_0_403 (.A1(n_0_298), .A2(shiftingAmount[1]), .B1(n_0_38), .B2(
      n_0_292), .ZN(n_0_355__0));
   OAI21_X1 i_0_404 (.A(n_0_277), .B1(n_0_8), .B2(n_0_120), .ZN(n_0_299));
   AOI21_X1 i_0_405 (.A(n_0_299), .B1(n_0_16), .B2(n_0_217), .ZN(n_0_300));
   OAI22_X1 i_0_406 (.A1(n_0_300), .A2(shiftingAmount[3]), .B1(n_0_17), .B2(
      n_0_266), .ZN(n_0_301));
   AOI22_X1 i_0_407 (.A1(n_0_287), .A2(shiftingAmount[2]), .B1(n_0_301), 
      .B2(n_0_20), .ZN(n_0_302));
   OAI22_X1 i_0_408 (.A1(n_0_295), .A2(n_0_38), .B1(n_0_302), .B2(
      shiftingAmount[1]), .ZN(n_0_356__0));
   OAI21_X1 i_0_409 (.A(n_0_277), .B1(n_0_8), .B2(n_0_172), .ZN(n_0_303));
   AOI21_X1 i_0_410 (.A(n_0_303), .B1(n_0_16), .B2(n_0_223), .ZN(n_0_304));
   OAI22_X1 i_0_411 (.A1(n_0_304), .A2(shiftingAmount[3]), .B1(n_0_17), .B2(
      n_0_272), .ZN(n_0_305));
   AOI22_X1 i_0_412 (.A1(n_0_291), .A2(shiftingAmount[2]), .B1(n_0_305), 
      .B2(n_0_20), .ZN(n_0_306));
   OAI22_X1 i_0_413 (.A1(n_0_298), .A2(n_0_38), .B1(n_0_306), .B2(
      shiftingAmount[1]), .ZN(n_0_357__0));
   AOI221_X1 i_0_414 (.A(n_0_278), .B1(shiftingAmount[5]), .B2(n_0_129), 
      .C1(n_0_16), .C2(n_0_229), .ZN(n_0_307));
   AOI22_X1 i_0_415 (.A1(n_0_279), .A2(shiftingAmount[3]), .B1(n_0_307), 
      .B2(n_0_17), .ZN(n_0_308));
   AOI22_X1 i_0_416 (.A1(n_0_308), .A2(n_0_20), .B1(n_0_294), .B2(
      shiftingAmount[2]), .ZN(n_0_309));
   OAI22_X1 i_0_417 (.A1(n_0_309), .A2(shiftingAmount[1]), .B1(n_0_38), .B2(
      n_0_302), .ZN(n_0_358__0));
   AOI221_X1 i_0_418 (.A(n_0_278), .B1(shiftingAmount[5]), .B2(n_0_136), 
      .C1(n_0_16), .C2(n_0_235), .ZN(n_0_310));
   AOI22_X1 i_0_419 (.A1(n_0_282), .A2(shiftingAmount[3]), .B1(n_0_310), 
      .B2(n_0_17), .ZN(n_0_311));
   AOI22_X1 i_0_420 (.A1(n_0_311), .A2(n_0_20), .B1(n_0_297), .B2(
      shiftingAmount[2]), .ZN(n_0_312));
   OAI22_X1 i_0_421 (.A1(n_0_312), .A2(shiftingAmount[1]), .B1(n_0_38), .B2(
      n_0_306), .ZN(n_0_359__0));
   AOI221_X1 i_0_422 (.A(n_0_278), .B1(n_0_16), .B2(n_0_241), .C1(
      shiftingAmount[5]), .C2(n_0_142), .ZN(n_0_313));
   OAI22_X1 i_0_423 (.A1(n_0_313), .A2(shiftingAmount[3]), .B1(n_0_286), 
      .B2(n_0_17), .ZN(n_0_314));
   AOI22_X1 i_0_424 (.A1(n_0_314), .A2(n_0_20), .B1(shiftingAmount[2]), .B2(
      n_0_301), .ZN(n_0_315));
   OAI22_X1 i_0_425 (.A1(n_0_309), .A2(n_0_38), .B1(n_0_315), .B2(
      shiftingAmount[1]), .ZN(n_0_360__0));
   AOI221_X1 i_0_426 (.A(n_0_278), .B1(n_0_16), .B2(n_0_247), .C1(
      shiftingAmount[5]), .C2(n_0_148), .ZN(n_0_316__1));
   OAI22_X1 i_0_427 (.A1(n_0_316__1), .A2(shiftingAmount[3]), .B1(n_0_290), 
      .B2(n_0_17), .ZN(n_0_317));
   AOI22_X1 i_0_428 (.A1(n_0_317), .A2(n_0_20), .B1(shiftingAmount[2]), .B2(
      n_0_305), .ZN(n_0_318__1));
   OAI22_X1 i_0_429 (.A1(n_0_312), .A2(n_0_38), .B1(n_0_318__1), .B2(
      shiftingAmount[1]), .ZN(n_0_361__0));
   AOI221_X1 i_0_430 (.A(n_0_278), .B1(shiftingAmount[5]), .B2(n_0_155), 
      .C1(n_0_16), .C2(n_0_253), .ZN(n_0_319));
   OAI22_X1 i_0_431 (.A1(n_0_293), .A2(n_0_17), .B1(n_0_319), .B2(
      shiftingAmount[3]), .ZN(n_0_320__1));
   AOI22_X1 i_0_432 (.A1(n_0_308), .A2(shiftingAmount[2]), .B1(n_0_320__1), 
      .B2(n_0_20), .ZN(n_0_321__1));
   OAI22_X1 i_0_433 (.A1(n_0_321__1), .A2(shiftingAmount[1]), .B1(n_0_38), 
      .B2(n_0_315), .ZN(n_0_362__0));
   AOI221_X1 i_0_434 (.A(n_0_278), .B1(n_0_16), .B2(n_0_259), .C1(
      shiftingAmount[5]), .C2(n_0_161), .ZN(n_0_322__1));
   AOI22_X1 i_0_435 (.A1(n_0_296), .A2(shiftingAmount[3]), .B1(n_0_322__1), 
      .B2(n_0_17), .ZN(n_0_323__1));
   AOI22_X1 i_0_436 (.A1(n_0_311), .A2(shiftingAmount[2]), .B1(n_0_323__1), 
      .B2(n_0_20), .ZN(n_0_324__1));
   OAI22_X1 i_0_437 (.A1(n_0_324__1), .A2(shiftingAmount[1]), .B1(n_0_38), 
      .B2(n_0_318__1), .ZN(n_0_363__0));
   AOI221_X1 i_0_438 (.A(n_0_278), .B1(n_0_16), .B2(n_0_265), .C1(
      shiftingAmount[5]), .C2(n_0_168), .ZN(n_0_325__1));
   OAI22_X1 i_0_439 (.A1(n_0_325__1), .A2(shiftingAmount[3]), .B1(n_0_300), 
      .B2(n_0_17), .ZN(n_0_326__1));
   AOI22_X1 i_0_440 (.A1(n_0_314), .A2(shiftingAmount[2]), .B1(n_0_326__1), 
      .B2(n_0_20), .ZN(n_0_327__1));
   OAI22_X1 i_0_441 (.A1(n_0_321__1), .A2(n_0_38), .B1(n_0_327__1), .B2(
      shiftingAmount[1]), .ZN(n_0_364__0));
   AOI221_X1 i_0_442 (.A(n_0_278), .B1(shiftingAmount[5]), .B2(n_0_175), 
      .C1(n_0_16), .C2(n_0_271), .ZN(n_0_328__1));
   OAI22_X1 i_0_443 (.A1(n_0_328__1), .A2(shiftingAmount[3]), .B1(n_0_304), 
      .B2(n_0_17), .ZN(n_0_329__1));
   AOI22_X1 i_0_444 (.A1(n_0_317), .A2(shiftingAmount[2]), .B1(n_0_329__1), 
      .B2(n_0_20), .ZN(n_0_330__1));
   OAI22_X1 i_0_445 (.A1(n_0_324__1), .A2(n_0_38), .B1(n_0_330__1), .B2(
      shiftingAmount[1]), .ZN(n_0_365__0));
   NAND2_X1 i_0_446 (.A1(n_0_276), .A2(n_0_8), .ZN(n_0_331__1));
   NAND2_X1 i_0_447 (.A1(n_0_331__1), .A2(n_0_17), .ZN(n_0_332__1));
   AOI21_X1 i_0_448 (.A(n_0_332__1), .B1(shiftingAmount[5]), .B2(n_0_181), 
      .ZN(n_0_333__1));
   AOI21_X1 i_0_449 (.A(n_0_333__1), .B1(n_0_307), .B2(shiftingAmount[3]), 
      .ZN(n_0_334__1));
   AOI22_X1 i_0_450 (.A1(n_0_320__1), .A2(shiftingAmount[2]), .B1(n_0_334__1), 
      .B2(n_0_20), .ZN(n_0_335__1));
   OAI22_X1 i_0_451 (.A1(n_0_335__1), .A2(shiftingAmount[1]), .B1(n_0_327__1), 
      .B2(n_0_38), .ZN(n_0_366__0));
   AOI21_X1 i_0_452 (.A(n_0_332__1), .B1(shiftingAmount[5]), .B2(n_0_187), 
      .ZN(n_0_336__1));
   AOI21_X1 i_0_453 (.A(n_0_336__1), .B1(n_0_310), .B2(shiftingAmount[3]), 
      .ZN(n_0_337__1));
   AOI22_X1 i_0_454 (.A1(n_0_323__1), .A2(shiftingAmount[2]), .B1(n_0_337__1), 
      .B2(n_0_20), .ZN(n_0_338__1));
   OAI22_X1 i_0_455 (.A1(n_0_338__1), .A2(shiftingAmount[1]), .B1(n_0_330__1), 
      .B2(n_0_38), .ZN(n_0_367__0));
   AOI21_X1 i_0_456 (.A(n_0_332__1), .B1(shiftingAmount[5]), .B2(n_0_193), 
      .ZN(n_0_339__1));
   AOI21_X1 i_0_457 (.A(n_0_339__1), .B1(n_0_313), .B2(shiftingAmount[3]), 
      .ZN(n_0_340__1));
   AOI22_X1 i_0_458 (.A1(n_0_326__1), .A2(shiftingAmount[2]), .B1(n_0_340__1), 
      .B2(n_0_20), .ZN(n_0_341__1));
   OAI22_X1 i_0_459 (.A1(n_0_335__1), .A2(n_0_38), .B1(n_0_341__1), .B2(
      shiftingAmount[1]), .ZN(n_0_368__0));
   AOI21_X1 i_0_460 (.A(n_0_332__1), .B1(shiftingAmount[5]), .B2(n_0_199), 
      .ZN(n_0_342__1));
   AOI21_X1 i_0_461 (.A(n_0_342__1), .B1(n_0_316__1), .B2(shiftingAmount[3]), 
      .ZN(n_0_343__1));
   AOI22_X1 i_0_462 (.A1(n_0_329__1), .A2(shiftingAmount[2]), .B1(n_0_343__1), 
      .B2(n_0_20), .ZN(n_0_344__1));
   OAI22_X1 i_0_463 (.A1(n_0_338__1), .A2(n_0_38), .B1(n_0_344__1), .B2(
      shiftingAmount[1]), .ZN(n_0_369__0));
   AOI21_X1 i_0_464 (.A(n_0_332__1), .B1(shiftingAmount[5]), .B2(n_0_205), 
      .ZN(n_0_345__1));
   AOI21_X1 i_0_465 (.A(n_0_345__1), .B1(n_0_319), .B2(shiftingAmount[3]), 
      .ZN(n_0_346__1));
   AOI22_X1 i_0_466 (.A1(n_0_334__1), .A2(shiftingAmount[2]), .B1(n_0_346__1), 
      .B2(n_0_20), .ZN(n_0_347__1));
   OAI22_X1 i_0_467 (.A1(n_0_347__1), .A2(shiftingAmount[1]), .B1(n_0_341__1), 
      .B2(n_0_38), .ZN(n_0_370__0));
   AOI21_X1 i_0_468 (.A(n_0_332__1), .B1(shiftingAmount[5]), .B2(n_0_211), 
      .ZN(n_0_348__1));
   AOI21_X1 i_0_469 (.A(n_0_348__1), .B1(n_0_322__1), .B2(shiftingAmount[3]), 
      .ZN(n_0_349__1));
   AOI22_X1 i_0_470 (.A1(n_0_337__1), .A2(shiftingAmount[2]), .B1(n_0_349__1), 
      .B2(n_0_20), .ZN(n_0_350__1));
   OAI22_X1 i_0_471 (.A1(n_0_350__1), .A2(shiftingAmount[1]), .B1(n_0_344__1), 
      .B2(n_0_38), .ZN(n_0_371__0));
   AOI21_X1 i_0_472 (.A(n_0_332__1), .B1(shiftingAmount[5]), .B2(n_0_217), 
      .ZN(n_0_351__1));
   AOI21_X1 i_0_473 (.A(n_0_351__1), .B1(n_0_325__1), .B2(shiftingAmount[3]), 
      .ZN(n_0_352__1));
   AOI22_X1 i_0_474 (.A1(n_0_340__1), .A2(shiftingAmount[2]), .B1(n_0_352__1), 
      .B2(n_0_20), .ZN(n_0_353__1));
   OAI22_X1 i_0_475 (.A1(n_0_347__1), .A2(n_0_38), .B1(n_0_353__1), .B2(
      shiftingAmount[1]), .ZN(n_0_372));
   AOI21_X1 i_0_476 (.A(n_0_332__1), .B1(shiftingAmount[5]), .B2(n_0_223), 
      .ZN(n_0_354__1));
   AOI21_X1 i_0_477 (.A(n_0_354__1), .B1(n_0_328__1), .B2(shiftingAmount[3]), 
      .ZN(n_0_355__1));
   AOI22_X1 i_0_478 (.A1(n_0_355__1), .A2(n_0_20), .B1(n_0_343__1), .B2(
      shiftingAmount[2]), .ZN(n_0_356__1));
   OAI22_X1 i_0_479 (.A1(n_0_350__1), .A2(n_0_38), .B1(n_0_356__1), .B2(
      shiftingAmount[1]), .ZN(n_0_373));
   INV_X1 i_0_480 (.A(n_0_229), .ZN(n_0_357__1));
   OAI21_X1 i_0_481 (.A(n_0_331__1), .B1(n_0_8), .B2(n_0_357__1), .ZN(n_0_358__1));
   AOI22_X1 i_0_482 (.A1(n_0_346__1), .A2(shiftingAmount[2]), .B1(n_0_20), 
      .B2(n_0_358__1), .ZN(n_0_359__1));
   OAI22_X1 i_0_483 (.A1(n_0_353__1), .A2(n_0_38), .B1(n_0_359__1), .B2(
      shiftingAmount[1]), .ZN(n_0_374));
   INV_X1 i_0_484 (.A(n_0_235), .ZN(n_0_360__1));
   OAI21_X1 i_0_485 (.A(n_0_331__1), .B1(n_0_8), .B2(n_0_360__1), .ZN(n_0_361__1));
   AOI22_X1 i_0_486 (.A1(n_0_349__1), .A2(shiftingAmount[2]), .B1(n_0_20), 
      .B2(n_0_361__1), .ZN(n_0_362__1));
   OAI22_X1 i_0_487 (.A1(n_0_356__1), .A2(n_0_38), .B1(n_0_362__1), .B2(
      shiftingAmount[1]), .ZN(n_0_375));
   INV_X1 i_0_488 (.A(n_0_241), .ZN(n_0_363__1));
   OAI21_X1 i_0_489 (.A(n_0_331__1), .B1(n_0_8), .B2(n_0_363__1), .ZN(n_0_364__1));
   AOI22_X1 i_0_490 (.A1(n_0_352__1), .A2(shiftingAmount[2]), .B1(n_0_364__1), 
      .B2(n_0_20), .ZN(n_0_365__1));
   OAI22_X1 i_0_491 (.A1(n_0_359__1), .A2(n_0_38), .B1(n_0_365__1), .B2(
      shiftingAmount[1]), .ZN(n_0_376));
   INV_X1 i_0_492 (.A(n_0_247), .ZN(n_0_366__1));
   OAI21_X1 i_0_493 (.A(n_0_331__1), .B1(n_0_8), .B2(n_0_366__1), .ZN(n_0_367__1));
   AOI22_X1 i_0_494 (.A1(n_0_355__1), .A2(shiftingAmount[2]), .B1(n_0_367__1), 
      .B2(n_0_20), .ZN(n_0_368__1));
   OAI22_X1 i_0_495 (.A1(n_0_362__1), .A2(n_0_38), .B1(n_0_368__1), .B2(
      shiftingAmount[1]), .ZN(n_0_377));
   INV_X1 i_0_496 (.A(n_0_259), .ZN(n_0_369__1));
   OAI21_X1 i_0_497 (.A(n_0_331__1), .B1(n_0_8), .B2(n_0_369__1), .ZN(n_0_381));
   NOR2_X1 i_0_498 (.A1(n_0_381), .A2(shiftingAmount[1]), .ZN(n_0_370__1));
   AOI21_X1 i_0_499 (.A(n_0_370__1), .B1(n_0_365__1), .B2(shiftingAmount[1]), 
      .ZN(n_0_378));
   AOI21_X1 i_0_500 (.A(n_0_370__1), .B1(n_0_368__1), .B2(shiftingAmount[1]), 
      .ZN(n_0_379));
   INV_X1 i_0_501 (.A(n_0_253), .ZN(n_0_371__1));
   OAI21_X1 i_0_502 (.A(n_0_331__1), .B1(n_0_8), .B2(n_0_371__1), .ZN(n_0_380));
   DFF_X1 \tempResult_reg[63]  (.D(n_162), .CK(n_145), .Q(tempResult[63]), .QN());
   DFF_X1 \tempResult_reg[62]  (.D(n_161), .CK(n_145), .Q(tempResult[62]), .QN());
   DFF_X1 \tempResult_reg[61]  (.D(n_160), .CK(n_145), .Q(tempResult[61]), .QN());
   DFF_X1 \tempResult_reg[60]  (.D(n_159), .CK(n_145), .Q(tempResult[60]), .QN());
   DFF_X1 \tempResult_reg[59]  (.D(n_158), .CK(n_145), .Q(tempResult[59]), .QN());
   DFF_X1 \tempResult_reg[58]  (.D(n_157), .CK(n_145), .Q(tempResult[58]), .QN());
   DFF_X1 \tempResult_reg[57]  (.D(n_156), .CK(n_145), .Q(tempResult[57]), .QN());
   DFF_X1 \tempResult_reg[56]  (.D(n_155), .CK(n_145), .Q(tempResult[56]), .QN());
   DFF_X1 \tempResult_reg[55]  (.D(n_154), .CK(n_145), .Q(tempResult[55]), .QN());
   DFF_X1 \tempResult_reg[54]  (.D(n_153), .CK(n_145), .Q(tempResult[54]), .QN());
   DFF_X1 \tempResult_reg[53]  (.D(n_152), .CK(n_145), .Q(tempResult[53]), .QN());
   DFF_X1 \tempResult_reg[52]  (.D(n_151), .CK(n_145), .Q(tempResult[52]), .QN());
   DFF_X1 \tempResult_reg[51]  (.D(n_150), .CK(n_145), .Q(tempResult[51]), .QN());
   DFF_X1 \tempResult_reg[50]  (.D(n_149), .CK(n_145), .Q(tempResult[50]), .QN());
   DFF_X1 \tempResult_reg[49]  (.D(n_148), .CK(n_145), .Q(tempResult[49]), .QN());
   DFF_X1 \tempResult_reg[48]  (.D(n_144), .CK(n_145), .Q(tempResult[48]), .QN());
   DFF_X1 \tempResult_reg[47]  (.D(n_143), .CK(n_145), .Q(tempResult[47]), .QN());
   DFF_X1 \tempResult_reg[46]  (.D(n_142), .CK(n_145), .Q(tempResult[46]), .QN());
   DFF_X1 \tempResult_reg[45]  (.D(n_141), .CK(n_145), .Q(tempResult[45]), .QN());
   DFF_X1 \tempResult_reg[44]  (.D(n_140), .CK(n_145), .Q(tempResult[44]), .QN());
   DFF_X1 \tempResult_reg[43]  (.D(n_139), .CK(n_145), .Q(tempResult[43]), .QN());
   DFF_X1 \tempResult_reg[42]  (.D(n_138), .CK(n_145), .Q(tempResult[42]), .QN());
   DFF_X1 \tempResult_reg[41]  (.D(n_137), .CK(n_145), .Q(tempResult[41]), .QN());
   DFF_X1 \tempResult_reg[40]  (.D(n_136), .CK(n_145), .Q(tempResult[40]), .QN());
   DFF_X1 \tempResult_reg[39]  (.D(n_135), .CK(n_145), .Q(tempResult[39]), .QN());
   DFF_X1 \tempResult_reg[38]  (.D(n_134), .CK(n_145), .Q(tempResult[38]), .QN());
   DFF_X1 \tempResult_reg[37]  (.D(n_133), .CK(n_145), .Q(tempResult[37]), .QN());
   DFF_X1 \tempResult_reg[36]  (.D(n_132), .CK(n_145), .Q(tempResult[36]), .QN());
   DFF_X1 \tempResult_reg[35]  (.D(n_131), .CK(n_145), .Q(tempResult[35]), .QN());
   DFF_X1 \tempResult_reg[34]  (.D(n_130), .CK(n_145), .Q(tempResult[34]), .QN());
   DFF_X1 \tempResult_reg[33]  (.D(n_129), .CK(n_145), .Q(tempResult[33]), .QN());
   DFF_X1 \tempResult_reg[32]  (.D(n_128), .CK(n_145), .Q(tempResult[32]), .QN());
   DFF_X1 \tempResult_reg[31]  (.D(n_127), .CK(n_145), .Q(tempResult[31]), .QN());
   DFF_X1 \tempResult_reg[30]  (.D(n_126), .CK(n_145), .Q(tempResult[30]), .QN());
   DFF_X1 \tempResult_reg[29]  (.D(n_125), .CK(n_145), .Q(tempResult[29]), .QN());
   DFF_X1 \tempResult_reg[28]  (.D(n_124), .CK(n_145), .Q(tempResult[28]), .QN());
   DFF_X1 \tempResult_reg[27]  (.D(n_123), .CK(n_145), .Q(tempResult[27]), .QN());
   DFF_X1 \tempResult_reg[26]  (.D(n_122), .CK(n_145), .Q(tempResult[26]), .QN());
   DFF_X1 \tempResult_reg[25]  (.D(n_121), .CK(n_145), .Q(tempResult[25]), .QN());
   DFF_X1 \tempResult_reg[24]  (.D(n_120), .CK(n_145), .Q(tempResult[24]), .QN());
   DFF_X1 \tempResult_reg[23]  (.D(n_119), .CK(n_145), .Q(tempResult[23]), .QN());
   DFF_X1 \tempResult_reg[22]  (.D(n_118), .CK(n_145), .Q(tempResult[22]), .QN());
   DFF_X1 \tempResult_reg[21]  (.D(n_117), .CK(n_145), .Q(tempResult[21]), .QN());
   DFF_X1 \tempResult_reg[20]  (.D(n_116), .CK(n_145), .Q(tempResult[20]), .QN());
   DFF_X1 \tempResult_reg[19]  (.D(n_115), .CK(n_145), .Q(tempResult[19]), .QN());
   DFF_X1 \tempResult_reg[18]  (.D(n_114), .CK(n_145), .Q(tempResult[18]), .QN());
   DFF_X1 \tempResult_reg[17]  (.D(n_113), .CK(n_145), .Q(tempResult[17]), .QN());
   DFF_X1 \tempResult_reg[16]  (.D(n_112), .CK(n_145), .Q(tempResult[16]), .QN());
   DFF_X1 \tempResult_reg[15]  (.D(n_111), .CK(n_145), .Q(tempResult[15]), .QN());
   DFF_X1 \tempResult_reg[14]  (.D(n_110), .CK(n_145), .Q(tempResult[14]), .QN());
   DFF_X1 \tempResult_reg[13]  (.D(n_109), .CK(n_145), .Q(tempResult[13]), .QN());
   DFF_X1 \tempResult_reg[12]  (.D(n_108), .CK(n_145), .Q(tempResult[12]), .QN());
   DFF_X1 \tempResult_reg[11]  (.D(n_107), .CK(n_145), .Q(tempResult[11]), .QN());
   DFF_X1 \tempResult_reg[10]  (.D(n_106), .CK(n_145), .Q(tempResult[10]), .QN());
   DFF_X1 \tempResult_reg[9]  (.D(n_105), .CK(n_145), .Q(tempResult[9]), .QN());
   DFF_X1 \tempResult_reg[8]  (.D(n_104), .CK(n_145), .Q(tempResult[8]), .QN());
   DFF_X1 \tempResult_reg[7]  (.D(n_103), .CK(n_145), .Q(tempResult[7]), .QN());
   DFF_X1 \tempResult_reg[6]  (.D(n_102), .CK(n_145), .Q(tempResult[6]), .QN());
   DFF_X1 \tempResult_reg[5]  (.D(n_101), .CK(n_145), .Q(tempResult[5]), .QN());
   DFF_X1 \tempResult_reg[4]  (.D(n_100), .CK(n_145), .Q(tempResult[4]), .QN());
   DFF_X1 \tempResult_reg[3]  (.D(n_99), .CK(n_145), .Q(tempResult[3]), .QN());
   DFF_X1 \tempResult_reg[2]  (.D(n_98), .CK(n_145), .Q(tempResult[2]), .QN());
   DFF_X1 \tempResult_reg[1]  (.D(n_97), .CK(n_145), .Q(tempResult[1]), .QN());
   DFF_X1 \tempResult_reg[0]  (.D(n_96), .CK(n_145), .Q(tempResult[0]), .QN());
   DFF_X1 \shiftingAmount_reg[5]  (.D(n_167), .CK(n_145), .Q(shiftingAmount[5]), 
      .QN());
   DFF_X1 \shiftingAmount_reg[4]  (.D(n_166), .CK(n_145), .Q(shiftingAmount[4]), 
      .QN());
   DFF_X1 \shiftingAmount_reg[3]  (.D(n_165), .CK(n_145), .Q(shiftingAmount[3]), 
      .QN());
   DFF_X1 \shiftingAmount_reg[2]  (.D(n_164), .CK(n_145), .Q(shiftingAmount[2]), 
      .QN());
   DFF_X1 \shiftingAmount_reg[1]  (.D(n_163), .CK(n_145), .Q(shiftingAmount[1]), 
      .QN());
   DFF_X1 \newB_reg[34]  (.D(in2[31]), .CK(n_146), .Q(newB[34]), .QN());
   DFF_X1 \newB_reg[31]  (.D(in2[30]), .CK(n_146), .Q(newB[31]), .QN());
   DFF_X1 \newB_reg[30]  (.D(in2[29]), .CK(n_146), .Q(newB[30]), .QN());
   DFF_X1 \newB_reg[29]  (.D(in2[28]), .CK(n_146), .Q(newB[29]), .QN());
   DFF_X1 \newB_reg[28]  (.D(in2[27]), .CK(n_146), .Q(newB[28]), .QN());
   DFF_X1 \newB_reg[27]  (.D(in2[26]), .CK(n_146), .Q(newB[27]), .QN());
   DFF_X1 \newB_reg[26]  (.D(in2[25]), .CK(n_146), .Q(newB[26]), .QN());
   DFF_X1 \newB_reg[25]  (.D(in2[24]), .CK(n_146), .Q(newB[25]), .QN());
   DFF_X1 \newB_reg[24]  (.D(in2[23]), .CK(n_146), .Q(newB[24]), .QN());
   DFF_X1 \newB_reg[23]  (.D(in2[22]), .CK(n_146), .Q(newB[23]), .QN());
   DFF_X1 \newB_reg[22]  (.D(in2[21]), .CK(n_146), .Q(newB[22]), .QN());
   DFF_X1 \newB_reg[21]  (.D(in2[20]), .CK(n_146), .Q(newB[21]), .QN());
   DFF_X1 \newB_reg[20]  (.D(in2[19]), .CK(n_146), .Q(newB[20]), .QN());
   DFF_X1 \newB_reg[19]  (.D(in2[18]), .CK(n_146), .Q(newB[19]), .QN());
   DFF_X1 \newB_reg[18]  (.D(in2[17]), .CK(n_146), .Q(newB[18]), .QN());
   DFF_X1 \newB_reg[17]  (.D(in2[16]), .CK(n_146), .Q(newB[17]), .QN());
   DFF_X1 \newB_reg[16]  (.D(in2[15]), .CK(n_146), .Q(newB[16]), .QN());
   DFF_X1 \newB_reg[15]  (.D(in2[14]), .CK(n_146), .Q(newB[15]), .QN());
   DFF_X1 \newB_reg[14]  (.D(in2[13]), .CK(n_146), .Q(newB[14]), .QN());
   DFF_X1 \newB_reg[13]  (.D(in2[12]), .CK(n_146), .Q(newB[13]), .QN());
   DFF_X1 \newB_reg[12]  (.D(in2[11]), .CK(n_146), .Q(newB[12]), .QN());
   DFF_X1 \newB_reg[11]  (.D(in2[10]), .CK(n_146), .Q(newB[11]), .QN());
   DFF_X1 \newB_reg[10]  (.D(in2[9]), .CK(n_146), .Q(newB[10]), .QN());
   DFF_X1 \newB_reg[9]  (.D(in2[8]), .CK(n_146), .Q(newB[9]), .QN());
   DFF_X1 \newB_reg[8]  (.D(in2[7]), .CK(n_146), .Q(newB[8]), .QN());
   DFF_X1 \newB_reg[7]  (.D(in2[6]), .CK(n_146), .Q(newB[7]), .QN());
   DFF_X1 \newB_reg[6]  (.D(in2[5]), .CK(n_146), .Q(newB[6]), .QN());
   DFF_X1 \newB_reg[5]  (.D(in2[4]), .CK(n_146), .Q(newB[5]), .QN());
   DFF_X1 \newB_reg[4]  (.D(in2[3]), .CK(n_146), .Q(newB[4]), .QN());
   DFF_X1 \newB_reg[3]  (.D(in2[2]), .CK(n_146), .Q(newB[3]), .QN());
   DFF_X1 \newB_reg[2]  (.D(in2[1]), .CK(n_146), .Q(newB[2]), .QN());
   DFF_X1 \newB_reg[1]  (.D(in2[0]), .CK(n_146), .Q(newB[1]), .QN());
   CLKGATETST_X1 clk_gate_tempResult_reg (.CK(clk), .E(n_147), .SE(1'b0), 
      .GCK(n_145));
   CLKGATETST_X1 clk_gate_Input1_1_Positive_reg (.CK(clk), .E(start), .SE(1'b0), 
      .GCK(n_146));
   DFF_X1 \Input1_1_Negative_reg[63]  (.D(n_63), .CK(n_146), .Q(
      Input1_1_Negative[63]), .QN());
   DFF_X1 \Input1_1_Negative_reg[15]  (.D(n_47), .CK(n_146), .Q(
      Input1_1_Negative[15]), .QN());
   DFF_X1 \Input1_1_Positive_reg[15]  (.D(in1[15]), .CK(n_146), .Q(
      Input1_1_Positive[15]), .QN());
   DFF_X1 \Input1_2_Negative_reg[17]  (.D(n_48), .CK(n_146), .Q(
      Input1_2_Negative[17]), .QN());
   DFF_X1 \Input1_2_Positive_reg[17]  (.D(in1[16]), .CK(n_146), .Q(
      Input1_2_Positive[17]), .QN());
   DFF_X1 \Input1_1_Negative_reg[7]  (.D(n_39), .CK(n_146), .Q(
      Input1_1_Negative[7]), .QN());
   DFF_X1 \Input1_1_Positive_reg[7]  (.D(in1[7]), .CK(n_146), .Q(
      Input1_1_Positive[7]), .QN());
   DFF_X1 \Input1_2_Negative_reg[9]  (.D(n_40), .CK(n_146), .Q(
      Input1_2_Negative[9]), .QN());
   DFF_X1 \Input1_2_Positive_reg[9]  (.D(in1[8]), .CK(n_146), .Q(
      Input1_2_Positive[9]), .QN());
   DFF_X1 \Input1_1_Negative_reg[23]  (.D(n_55), .CK(n_146), .Q(
      Input1_1_Negative[23]), .QN());
   DFF_X1 \Input1_1_Positive_reg[23]  (.D(in1[23]), .CK(n_146), .Q(
      Input1_1_Positive[23]), .QN());
   DFF_X1 \Input1_2_Negative_reg[25]  (.D(n_56), .CK(n_146), .Q(
      Input1_2_Negative[25]), .QN());
   DFF_X1 \Input1_2_Positive_reg[25]  (.D(in1[24]), .CK(n_146), .Q(
      Input1_2_Positive[25]), .QN());
   DFF_X1 \Input1_1_Negative_reg[3]  (.D(n_35), .CK(n_146), .Q(
      Input1_1_Negative[3]), .QN());
   DFF_X1 \Input1_1_Positive_reg[3]  (.D(in1[3]), .CK(n_146), .Q(
      Input1_1_Positive[3]), .QN());
   DFF_X1 \Input1_2_Negative_reg[5]  (.D(n_36), .CK(n_146), .Q(
      Input1_2_Negative[5]), .QN());
   DFF_X1 \Input1_2_Positive_reg[5]  (.D(in1[4]), .CK(n_146), .Q(
      Input1_2_Positive[5]), .QN());
   DFF_X1 \Input1_1_Negative_reg[19]  (.D(n_51), .CK(n_146), .Q(
      Input1_1_Negative[19]), .QN());
   DFF_X1 \Input1_1_Positive_reg[19]  (.D(in1[19]), .CK(n_146), .Q(
      Input1_1_Positive[19]), .QN());
   DFF_X1 \Input1_2_Negative_reg[21]  (.D(n_52), .CK(n_146), .Q(
      Input1_2_Negative[21]), .QN());
   DFF_X1 \Input1_2_Positive_reg[21]  (.D(in1[20]), .CK(n_146), .Q(
      Input1_2_Positive[21]), .QN());
   DFF_X1 \Input1_1_Negative_reg[11]  (.D(n_43), .CK(n_146), .Q(
      Input1_1_Negative[11]), .QN());
   DFF_X1 \Input1_1_Positive_reg[11]  (.D(in1[11]), .CK(n_146), .Q(
      Input1_1_Positive[11]), .QN());
   DFF_X1 \Input1_2_Negative_reg[13]  (.D(n_44), .CK(n_146), .Q(
      Input1_2_Negative[13]), .QN());
   DFF_X1 \Input1_2_Positive_reg[13]  (.D(in1[12]), .CK(n_146), .Q(
      Input1_2_Positive[13]), .QN());
   DFF_X1 \Input1_1_Negative_reg[27]  (.D(n_59), .CK(n_146), .Q(
      Input1_1_Negative[27]), .QN());
   DFF_X1 \Input1_1_Positive_reg[27]  (.D(in1[27]), .CK(n_146), .Q(
      Input1_1_Positive[27]), .QN());
   DFF_X1 \Input1_2_Negative_reg[29]  (.D(n_60), .CK(n_146), .Q(
      Input1_2_Negative[29]), .QN());
   DFF_X1 \Input1_2_Positive_reg[29]  (.D(in1[28]), .CK(n_146), .Q(
      Input1_2_Positive[29]), .QN());
   DFF_X1 \Input1_1_Negative_reg[1]  (.D(n_33), .CK(n_146), .Q(
      Input1_1_Negative[1]), .QN());
   DFF_X1 \Input1_1_Positive_reg[1]  (.D(in1[1]), .CK(n_146), .Q(
      Input1_1_Positive[1]), .QN());
   DFF_X1 \Input1_2_Negative_reg[3]  (.D(n_34), .CK(n_146), .Q(
      Input1_2_Negative[3]), .QN());
   DFF_X1 \Input1_2_Positive_reg[3]  (.D(in1[2]), .CK(n_146), .Q(
      Input1_2_Positive[3]), .QN());
   DFF_X1 \Input1_1_Negative_reg[17]  (.D(n_49), .CK(n_146), .Q(
      Input1_1_Negative[17]), .QN());
   DFF_X1 \Input1_1_Positive_reg[17]  (.D(in1[17]), .CK(n_146), .Q(
      Input1_1_Positive[17]), .QN());
   DFF_X1 \Input1_2_Negative_reg[19]  (.D(n_50), .CK(n_146), .Q(
      Input1_2_Negative[19]), .QN());
   DFF_X1 \Input1_2_Positive_reg[19]  (.D(in1[18]), .CK(n_146), .Q(
      Input1_2_Positive[19]), .QN());
   DFF_X1 \Input1_1_Negative_reg[9]  (.D(n_41), .CK(n_146), .Q(
      Input1_1_Negative[9]), .QN());
   DFF_X1 \Input1_1_Positive_reg[9]  (.D(in1[9]), .CK(n_146), .Q(
      Input1_1_Positive[9]), .QN());
   DFF_X1 \Input1_2_Negative_reg[11]  (.D(n_42), .CK(n_146), .Q(
      Input1_2_Negative[11]), .QN());
   DFF_X1 \Input1_2_Positive_reg[11]  (.D(in1[10]), .CK(n_146), .Q(
      Input1_2_Positive[11]), .QN());
   DFF_X1 \Input1_1_Negative_reg[25]  (.D(n_57), .CK(n_146), .Q(
      Input1_1_Negative[25]), .QN());
   DFF_X1 \Input1_1_Positive_reg[25]  (.D(in1[25]), .CK(n_146), .Q(
      Input1_1_Positive[25]), .QN());
   DFF_X1 \Input1_2_Negative_reg[27]  (.D(n_58), .CK(n_146), .Q(
      Input1_2_Negative[27]), .QN());
   DFF_X1 \Input1_2_Positive_reg[27]  (.D(in1[26]), .CK(n_146), .Q(
      Input1_2_Positive[27]), .QN());
   DFF_X1 \Input1_1_Negative_reg[5]  (.D(n_37), .CK(n_146), .Q(
      Input1_1_Negative[5]), .QN());
   DFF_X1 \Input1_1_Positive_reg[5]  (.D(in1[5]), .CK(n_146), .Q(
      Input1_1_Positive[5]), .QN());
   DFF_X1 \Input1_2_Negative_reg[7]  (.D(n_38), .CK(n_146), .Q(
      Input1_2_Negative[7]), .QN());
   DFF_X1 \Input1_2_Positive_reg[7]  (.D(in1[6]), .CK(n_146), .Q(
      Input1_2_Positive[7]), .QN());
   DFF_X1 \Input1_1_Negative_reg[21]  (.D(n_53), .CK(n_146), .Q(
      Input1_1_Negative[21]), .QN());
   DFF_X1 \Input1_1_Positive_reg[21]  (.D(in1[21]), .CK(n_146), .Q(
      Input1_1_Positive[21]), .QN());
   DFF_X1 \Input1_2_Negative_reg[23]  (.D(n_54), .CK(n_146), .Q(
      Input1_2_Negative[23]), .QN());
   DFF_X1 \Input1_2_Positive_reg[23]  (.D(in1[22]), .CK(n_146), .Q(
      Input1_2_Positive[23]), .QN());
   DFF_X1 \Input1_1_Negative_reg[13]  (.D(n_45), .CK(n_146), .Q(
      Input1_1_Negative[13]), .QN());
   DFF_X1 \Input1_1_Positive_reg[13]  (.D(in1[13]), .CK(n_146), .Q(
      Input1_1_Positive[13]), .QN());
   DFF_X1 \Input1_2_Negative_reg[15]  (.D(n_46), .CK(n_146), .Q(
      Input1_2_Negative[15]), .QN());
   DFF_X1 \Input1_2_Positive_reg[15]  (.D(in1[14]), .CK(n_146), .Q(
      Input1_2_Positive[15]), .QN());
   DFF_X1 \Input1_1_Negative_reg[29]  (.D(n_61), .CK(n_146), .Q(
      Input1_1_Negative[29]), .QN());
   DFF_X1 \Input1_1_Positive_reg[29]  (.D(in1[29]), .CK(n_146), .Q(
      Input1_1_Positive[29]), .QN());
   DFF_X1 \Input1_2_Negative_reg[31]  (.D(n_62), .CK(n_146), .Q(
      Input1_2_Negative[31]), .QN());
   DFF_X1 \Input1_2_Positive_reg[31]  (.D(in1[30]), .CK(n_146), .Q(
      Input1_2_Positive[31]), .QN());
   DFF_X1 \Input1_2_Positive_reg[1]  (.D(in1[0]), .CK(n_146), .Q(
      Input1_2_Positive[1]), .QN());
   DFF_X1 \Input1_1_Positive_reg[63]  (.D(in1[31]), .CK(n_146), .Q(
      Input1_1_Positive[63]), .QN());
   INV_X1 i_14 (.A(n_168), .ZN(n_147));
endmodule

module Radix4(clk, inputA, inputB, outResult, start);
   input clk;
   input [31:0]inputA;
   input [31:0]inputB;
   output [63:0]outResult;
   input start;

   wire [63:0]result;
   wire [31:0]B;
   wire [31:0]A;

   Noaman_4_Booth mult (.start(start), .clk(clk), .in1(A), .in2(B), .result(
      result));
   DFF_X1 \outResult_reg[63]  (.D(result[63]), .CK(clk), .Q(outResult[63]), 
      .QN());
   DFF_X1 \outResult_reg[62]  (.D(result[62]), .CK(clk), .Q(outResult[62]), 
      .QN());
   DFF_X1 \outResult_reg[61]  (.D(result[61]), .CK(clk), .Q(outResult[61]), 
      .QN());
   DFF_X1 \outResult_reg[60]  (.D(result[60]), .CK(clk), .Q(outResult[60]), 
      .QN());
   DFF_X1 \outResult_reg[59]  (.D(result[59]), .CK(clk), .Q(outResult[59]), 
      .QN());
   DFF_X1 \outResult_reg[58]  (.D(result[58]), .CK(clk), .Q(outResult[58]), 
      .QN());
   DFF_X1 \outResult_reg[57]  (.D(result[57]), .CK(clk), .Q(outResult[57]), 
      .QN());
   DFF_X1 \outResult_reg[56]  (.D(result[56]), .CK(clk), .Q(outResult[56]), 
      .QN());
   DFF_X1 \outResult_reg[55]  (.D(result[55]), .CK(clk), .Q(outResult[55]), 
      .QN());
   DFF_X1 \outResult_reg[54]  (.D(result[54]), .CK(clk), .Q(outResult[54]), 
      .QN());
   DFF_X1 \outResult_reg[53]  (.D(result[53]), .CK(clk), .Q(outResult[53]), 
      .QN());
   DFF_X1 \outResult_reg[52]  (.D(result[52]), .CK(clk), .Q(outResult[52]), 
      .QN());
   DFF_X1 \outResult_reg[51]  (.D(result[51]), .CK(clk), .Q(outResult[51]), 
      .QN());
   DFF_X1 \outResult_reg[50]  (.D(result[50]), .CK(clk), .Q(outResult[50]), 
      .QN());
   DFF_X1 \outResult_reg[49]  (.D(result[49]), .CK(clk), .Q(outResult[49]), 
      .QN());
   DFF_X1 \outResult_reg[48]  (.D(result[48]), .CK(clk), .Q(outResult[48]), 
      .QN());
   DFF_X1 \outResult_reg[47]  (.D(result[47]), .CK(clk), .Q(outResult[47]), 
      .QN());
   DFF_X1 \outResult_reg[46]  (.D(result[46]), .CK(clk), .Q(outResult[46]), 
      .QN());
   DFF_X1 \outResult_reg[45]  (.D(result[45]), .CK(clk), .Q(outResult[45]), 
      .QN());
   DFF_X1 \outResult_reg[44]  (.D(result[44]), .CK(clk), .Q(outResult[44]), 
      .QN());
   DFF_X1 \outResult_reg[43]  (.D(result[43]), .CK(clk), .Q(outResult[43]), 
      .QN());
   DFF_X1 \outResult_reg[42]  (.D(result[42]), .CK(clk), .Q(outResult[42]), 
      .QN());
   DFF_X1 \outResult_reg[41]  (.D(result[41]), .CK(clk), .Q(outResult[41]), 
      .QN());
   DFF_X1 \outResult_reg[40]  (.D(result[40]), .CK(clk), .Q(outResult[40]), 
      .QN());
   DFF_X1 \outResult_reg[39]  (.D(result[39]), .CK(clk), .Q(outResult[39]), 
      .QN());
   DFF_X1 \outResult_reg[38]  (.D(result[38]), .CK(clk), .Q(outResult[38]), 
      .QN());
   DFF_X1 \outResult_reg[37]  (.D(result[37]), .CK(clk), .Q(outResult[37]), 
      .QN());
   DFF_X1 \outResult_reg[36]  (.D(result[36]), .CK(clk), .Q(outResult[36]), 
      .QN());
   DFF_X1 \outResult_reg[35]  (.D(result[35]), .CK(clk), .Q(outResult[35]), 
      .QN());
   DFF_X1 \outResult_reg[34]  (.D(result[34]), .CK(clk), .Q(outResult[34]), 
      .QN());
   DFF_X1 \outResult_reg[33]  (.D(result[33]), .CK(clk), .Q(outResult[33]), 
      .QN());
   DFF_X1 \outResult_reg[32]  (.D(result[32]), .CK(clk), .Q(outResult[32]), 
      .QN());
   DFF_X1 \outResult_reg[31]  (.D(result[31]), .CK(clk), .Q(outResult[31]), 
      .QN());
   DFF_X1 \outResult_reg[30]  (.D(result[30]), .CK(clk), .Q(outResult[30]), 
      .QN());
   DFF_X1 \outResult_reg[29]  (.D(result[29]), .CK(clk), .Q(outResult[29]), 
      .QN());
   DFF_X1 \outResult_reg[28]  (.D(result[28]), .CK(clk), .Q(outResult[28]), 
      .QN());
   DFF_X1 \outResult_reg[27]  (.D(result[27]), .CK(clk), .Q(outResult[27]), 
      .QN());
   DFF_X1 \outResult_reg[26]  (.D(result[26]), .CK(clk), .Q(outResult[26]), 
      .QN());
   DFF_X1 \outResult_reg[25]  (.D(result[25]), .CK(clk), .Q(outResult[25]), 
      .QN());
   DFF_X1 \outResult_reg[24]  (.D(result[24]), .CK(clk), .Q(outResult[24]), 
      .QN());
   DFF_X1 \outResult_reg[23]  (.D(result[23]), .CK(clk), .Q(outResult[23]), 
      .QN());
   DFF_X1 \outResult_reg[22]  (.D(result[22]), .CK(clk), .Q(outResult[22]), 
      .QN());
   DFF_X1 \outResult_reg[21]  (.D(result[21]), .CK(clk), .Q(outResult[21]), 
      .QN());
   DFF_X1 \outResult_reg[20]  (.D(result[20]), .CK(clk), .Q(outResult[20]), 
      .QN());
   DFF_X1 \outResult_reg[19]  (.D(result[19]), .CK(clk), .Q(outResult[19]), 
      .QN());
   DFF_X1 \outResult_reg[18]  (.D(result[18]), .CK(clk), .Q(outResult[18]), 
      .QN());
   DFF_X1 \outResult_reg[17]  (.D(result[17]), .CK(clk), .Q(outResult[17]), 
      .QN());
   DFF_X1 \outResult_reg[16]  (.D(result[16]), .CK(clk), .Q(outResult[16]), 
      .QN());
   DFF_X1 \outResult_reg[15]  (.D(result[15]), .CK(clk), .Q(outResult[15]), 
      .QN());
   DFF_X1 \outResult_reg[14]  (.D(result[14]), .CK(clk), .Q(outResult[14]), 
      .QN());
   DFF_X1 \outResult_reg[13]  (.D(result[13]), .CK(clk), .Q(outResult[13]), 
      .QN());
   DFF_X1 \outResult_reg[12]  (.D(result[12]), .CK(clk), .Q(outResult[12]), 
      .QN());
   DFF_X1 \outResult_reg[11]  (.D(result[11]), .CK(clk), .Q(outResult[11]), 
      .QN());
   DFF_X1 \outResult_reg[10]  (.D(result[10]), .CK(clk), .Q(outResult[10]), 
      .QN());
   DFF_X1 \outResult_reg[9]  (.D(result[9]), .CK(clk), .Q(outResult[9]), .QN());
   DFF_X1 \outResult_reg[8]  (.D(result[8]), .CK(clk), .Q(outResult[8]), .QN());
   DFF_X1 \outResult_reg[7]  (.D(result[7]), .CK(clk), .Q(outResult[7]), .QN());
   DFF_X1 \outResult_reg[6]  (.D(result[6]), .CK(clk), .Q(outResult[6]), .QN());
   DFF_X1 \outResult_reg[5]  (.D(result[5]), .CK(clk), .Q(outResult[5]), .QN());
   DFF_X1 \outResult_reg[4]  (.D(result[4]), .CK(clk), .Q(outResult[4]), .QN());
   DFF_X1 \outResult_reg[3]  (.D(result[3]), .CK(clk), .Q(outResult[3]), .QN());
   DFF_X1 \outResult_reg[2]  (.D(result[2]), .CK(clk), .Q(outResult[2]), .QN());
   DFF_X1 \outResult_reg[1]  (.D(result[1]), .CK(clk), .Q(outResult[1]), .QN());
   DFF_X1 \outResult_reg[0]  (.D(result[0]), .CK(clk), .Q(outResult[0]), .QN());
   DFF_X1 \B_reg[31]  (.D(inputB[31]), .CK(clk), .Q(B[31]), .QN());
   DFF_X1 \B_reg[30]  (.D(inputB[30]), .CK(clk), .Q(B[30]), .QN());
   DFF_X1 \B_reg[29]  (.D(inputB[29]), .CK(clk), .Q(B[29]), .QN());
   DFF_X1 \B_reg[28]  (.D(inputB[28]), .CK(clk), .Q(B[28]), .QN());
   DFF_X1 \B_reg[27]  (.D(inputB[27]), .CK(clk), .Q(B[27]), .QN());
   DFF_X1 \B_reg[26]  (.D(inputB[26]), .CK(clk), .Q(B[26]), .QN());
   DFF_X1 \B_reg[25]  (.D(inputB[25]), .CK(clk), .Q(B[25]), .QN());
   DFF_X1 \B_reg[24]  (.D(inputB[24]), .CK(clk), .Q(B[24]), .QN());
   DFF_X1 \B_reg[23]  (.D(inputB[23]), .CK(clk), .Q(B[23]), .QN());
   DFF_X1 \B_reg[22]  (.D(inputB[22]), .CK(clk), .Q(B[22]), .QN());
   DFF_X1 \B_reg[21]  (.D(inputB[21]), .CK(clk), .Q(B[21]), .QN());
   DFF_X1 \B_reg[20]  (.D(inputB[20]), .CK(clk), .Q(B[20]), .QN());
   DFF_X1 \B_reg[19]  (.D(inputB[19]), .CK(clk), .Q(B[19]), .QN());
   DFF_X1 \B_reg[18]  (.D(inputB[18]), .CK(clk), .Q(B[18]), .QN());
   DFF_X1 \B_reg[17]  (.D(inputB[17]), .CK(clk), .Q(B[17]), .QN());
   DFF_X1 \B_reg[16]  (.D(inputB[16]), .CK(clk), .Q(B[16]), .QN());
   DFF_X1 \B_reg[15]  (.D(inputB[15]), .CK(clk), .Q(B[15]), .QN());
   DFF_X1 \B_reg[14]  (.D(inputB[14]), .CK(clk), .Q(B[14]), .QN());
   DFF_X1 \B_reg[13]  (.D(inputB[13]), .CK(clk), .Q(B[13]), .QN());
   DFF_X1 \B_reg[12]  (.D(inputB[12]), .CK(clk), .Q(B[12]), .QN());
   DFF_X1 \B_reg[11]  (.D(inputB[11]), .CK(clk), .Q(B[11]), .QN());
   DFF_X1 \B_reg[10]  (.D(inputB[10]), .CK(clk), .Q(B[10]), .QN());
   DFF_X1 \B_reg[9]  (.D(inputB[9]), .CK(clk), .Q(B[9]), .QN());
   DFF_X1 \B_reg[8]  (.D(inputB[8]), .CK(clk), .Q(B[8]), .QN());
   DFF_X1 \B_reg[7]  (.D(inputB[7]), .CK(clk), .Q(B[7]), .QN());
   DFF_X1 \B_reg[6]  (.D(inputB[6]), .CK(clk), .Q(B[6]), .QN());
   DFF_X1 \B_reg[5]  (.D(inputB[5]), .CK(clk), .Q(B[5]), .QN());
   DFF_X1 \B_reg[4]  (.D(inputB[4]), .CK(clk), .Q(B[4]), .QN());
   DFF_X1 \B_reg[3]  (.D(inputB[3]), .CK(clk), .Q(B[3]), .QN());
   DFF_X1 \B_reg[2]  (.D(inputB[2]), .CK(clk), .Q(B[2]), .QN());
   DFF_X1 \B_reg[1]  (.D(inputB[1]), .CK(clk), .Q(B[1]), .QN());
   DFF_X1 \B_reg[0]  (.D(inputB[0]), .CK(clk), .Q(B[0]), .QN());
   DFF_X1 \A_reg[31]  (.D(inputA[31]), .CK(clk), .Q(A[31]), .QN());
   DFF_X1 \A_reg[30]  (.D(inputA[30]), .CK(clk), .Q(A[30]), .QN());
   DFF_X1 \A_reg[29]  (.D(inputA[29]), .CK(clk), .Q(A[29]), .QN());
   DFF_X1 \A_reg[28]  (.D(inputA[28]), .CK(clk), .Q(A[28]), .QN());
   DFF_X1 \A_reg[27]  (.D(inputA[27]), .CK(clk), .Q(A[27]), .QN());
   DFF_X1 \A_reg[26]  (.D(inputA[26]), .CK(clk), .Q(A[26]), .QN());
   DFF_X1 \A_reg[25]  (.D(inputA[25]), .CK(clk), .Q(A[25]), .QN());
   DFF_X1 \A_reg[24]  (.D(inputA[24]), .CK(clk), .Q(A[24]), .QN());
   DFF_X1 \A_reg[23]  (.D(inputA[23]), .CK(clk), .Q(A[23]), .QN());
   DFF_X1 \A_reg[22]  (.D(inputA[22]), .CK(clk), .Q(A[22]), .QN());
   DFF_X1 \A_reg[21]  (.D(inputA[21]), .CK(clk), .Q(A[21]), .QN());
   DFF_X1 \A_reg[20]  (.D(inputA[20]), .CK(clk), .Q(A[20]), .QN());
   DFF_X1 \A_reg[19]  (.D(inputA[19]), .CK(clk), .Q(A[19]), .QN());
   DFF_X1 \A_reg[18]  (.D(inputA[18]), .CK(clk), .Q(A[18]), .QN());
   DFF_X1 \A_reg[17]  (.D(inputA[17]), .CK(clk), .Q(A[17]), .QN());
   DFF_X1 \A_reg[16]  (.D(inputA[16]), .CK(clk), .Q(A[16]), .QN());
   DFF_X1 \A_reg[15]  (.D(inputA[15]), .CK(clk), .Q(A[15]), .QN());
   DFF_X1 \A_reg[14]  (.D(inputA[14]), .CK(clk), .Q(A[14]), .QN());
   DFF_X1 \A_reg[13]  (.D(inputA[13]), .CK(clk), .Q(A[13]), .QN());
   DFF_X1 \A_reg[12]  (.D(inputA[12]), .CK(clk), .Q(A[12]), .QN());
   DFF_X1 \A_reg[11]  (.D(inputA[11]), .CK(clk), .Q(A[11]), .QN());
   DFF_X1 \A_reg[10]  (.D(inputA[10]), .CK(clk), .Q(A[10]), .QN());
   DFF_X1 \A_reg[9]  (.D(inputA[9]), .CK(clk), .Q(A[9]), .QN());
   DFF_X1 \A_reg[8]  (.D(inputA[8]), .CK(clk), .Q(A[8]), .QN());
   DFF_X1 \A_reg[7]  (.D(inputA[7]), .CK(clk), .Q(A[7]), .QN());
   DFF_X1 \A_reg[6]  (.D(inputA[6]), .CK(clk), .Q(A[6]), .QN());
   DFF_X1 \A_reg[5]  (.D(inputA[5]), .CK(clk), .Q(A[5]), .QN());
   DFF_X1 \A_reg[4]  (.D(inputA[4]), .CK(clk), .Q(A[4]), .QN());
   DFF_X1 \A_reg[3]  (.D(inputA[3]), .CK(clk), .Q(A[3]), .QN());
   DFF_X1 \A_reg[2]  (.D(inputA[2]), .CK(clk), .Q(A[2]), .QN());
   DFF_X1 \A_reg[1]  (.D(inputA[1]), .CK(clk), .Q(A[1]), .QN());
   DFF_X1 \A_reg[0]  (.D(inputA[0]), .CK(clk), .Q(A[0]), .QN());
endmodule
