/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Dec 27 14:02:28 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 748255416 */

module datapath(p_0, a);
   output [31:0]p_0;
   input [31:0]a;

   AOI21_X1 i_0 (.A(n_62), .B1(a[1]), .B2(a[0]), .ZN(p_0[1]));
   AOI21_X1 i_1 (.A(n_60), .B1(a[2]), .B2(n_61), .ZN(p_0[2]));
   AOI21_X1 i_2 (.A(n_58), .B1(a[3]), .B2(n_59), .ZN(p_0[3]));
   AOI21_X1 i_3 (.A(n_5), .B1(a[4]), .B2(n_57), .ZN(p_0[4]));
   AOI21_X1 i_5 (.A(n_1), .B1(a[6]), .B2(n_2), .ZN(p_0[6]));
   AOI21_X1 i_6 (.A(n_55), .B1(a[7]), .B2(n_0), .ZN(p_0[7]));
   INV_X1 i_7 (.A(n_1), .ZN(n_0));
   NOR2_X1 i_8 (.A1(n_57), .A2(n_56), .ZN(n_1));
   INV_X1 i_9 (.A(n_3), .ZN(n_2));
   AOI21_X1 i_13 (.A(n_11), .B1(a[8]), .B2(n_54), .ZN(p_0[8]));
   AOI21_X1 i_15 (.A(n_7), .B1(a[10]), .B2(n_8), .ZN(p_0[10]));
   AOI21_X1 i_16 (.A(n_52), .B1(a[11]), .B2(n_6), .ZN(p_0[11]));
   INV_X1 i_17 (.A(n_7), .ZN(n_6));
   NOR2_X1 i_18 (.A1(n_54), .A2(n_53), .ZN(n_7));
   INV_X1 i_19 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_23 (.A(n_17), .B1(a[12]), .B2(n_51), .ZN(p_0[12]));
   AOI21_X1 i_25 (.A(n_13), .B1(a[14]), .B2(n_14), .ZN(p_0[14]));
   AOI21_X1 i_26 (.A(n_49), .B1(a[15]), .B2(n_12), .ZN(p_0[15]));
   INV_X1 i_27 (.A(n_13), .ZN(n_12));
   NOR2_X1 i_28 (.A1(n_51), .A2(n_50), .ZN(n_13));
   INV_X1 i_29 (.A(n_15), .ZN(n_14));
   AOI21_X1 i_33 (.A(n_23), .B1(a[16]), .B2(n_48), .ZN(p_0[16]));
   AOI21_X1 i_34 (.A(n_21), .B1(a[17]), .B2(n_22), .ZN(p_0[17]));
   AOI21_X1 i_35 (.A(n_19), .B1(a[18]), .B2(n_20), .ZN(p_0[18]));
   AOI21_X1 i_36 (.A(n_45), .B1(a[19]), .B2(n_18), .ZN(p_0[19]));
   INV_X1 i_37 (.A(n_19), .ZN(n_18));
   NOR2_X1 i_38 (.A1(n_48), .A2(n_46), .ZN(n_19));
   INV_X1 i_39 (.A(n_21), .ZN(n_20));
   NOR2_X1 i_40 (.A1(a[17]), .A2(n_22), .ZN(n_21));
   INV_X1 i_41 (.A(n_23), .ZN(n_22));
   NOR2_X1 i_42 (.A1(a[16]), .A2(n_48), .ZN(n_23));
   AOI21_X1 i_43 (.A(n_25), .B1(a[20]), .B2(n_44), .ZN(p_0[20]));
   NOR2_X1 i_46 (.A1(a[20]), .A2(n_44), .ZN(n_25));
   AOI21_X1 i_64 (.A(n_37), .B1(a[30]), .B2(n_35), .ZN(p_0[30]));
   INV_X1 i_65 (.A(n_36), .ZN(n_35));
   XNOR2_X1 i_67 (.A(a[31]), .B(n_37), .ZN(p_0[31]));
   NOR4_X1 i_68 (.A1(a[29]), .A2(a[28]), .A3(a[30]), .A4(n_38), .ZN(n_37));
   INV_X1 i_4 (.A(n_4), .ZN(n_36));
   OR2_X1 i_10 (.A1(n_74), .A2(a[29]), .ZN(n_4));
   INV_X1 i_11 (.A(n_39), .ZN(n_15));
   INV_X1 i_12 (.A(n_29), .ZN(n_9));
   INV_X1 i_14 (.A(n_10), .ZN(n_3));
   NAND2_X1 i_20 (.A1(n_5), .A2(n_26), .ZN(n_10));
   INV_X1 i_21 (.A(n_16), .ZN(n_5));
   XNOR2_X1 i_22 (.A(n_16), .B(n_26), .ZN(p_0[5]));
   NAND2_X1 i_24 (.A1(n_58), .A2(n_24), .ZN(n_16));
   INV_X1 i_30 (.A(a[4]), .ZN(n_24));
   INV_X1 i_31 (.A(a[5]), .ZN(n_26));
   INV_X1 i_32 (.A(n_27), .ZN(p_0[9]));
   NAND2_X1 i_44 (.A1(n_29), .A2(n_28), .ZN(n_27));
   NAND2_X1 i_45 (.A1(n_30), .A2(a[9]), .ZN(n_28));
   NAND2_X1 i_47 (.A1(n_11), .A2(n_32), .ZN(n_29));
   INV_X1 i_48 (.A(n_30), .ZN(n_11));
   NAND2_X1 i_49 (.A1(n_55), .A2(n_31), .ZN(n_30));
   INV_X1 i_50 (.A(a[8]), .ZN(n_31));
   INV_X1 i_51 (.A(a[9]), .ZN(n_32));
   INV_X1 i_52 (.A(n_33), .ZN(p_0[13]));
   NAND2_X1 i_53 (.A1(n_39), .A2(n_34), .ZN(n_33));
   NAND2_X1 i_54 (.A1(n_40), .A2(a[13]), .ZN(n_34));
   NAND2_X1 i_55 (.A1(n_17), .A2(n_42), .ZN(n_39));
   INV_X1 i_56 (.A(n_40), .ZN(n_17));
   NAND2_X1 i_57 (.A1(n_52), .A2(n_41), .ZN(n_40));
   INV_X1 i_58 (.A(a[12]), .ZN(n_41));
   INV_X1 i_59 (.A(a[13]), .ZN(n_42));
   AOI21_X1 i_60 (.A(n_43), .B1(n_47), .B2(a[21]), .ZN(p_0[21]));
   INV_X1 i_61 (.A(n_63), .ZN(n_43));
   INV_X1 i_62 (.A(n_25), .ZN(n_47));
   AOI21_X1 i_63 (.A(n_84), .B1(n_63), .B2(a[22]), .ZN(p_0[22]));
   NAND3_X1 i_66 (.A1(n_45), .A2(n_65), .A3(n_64), .ZN(n_63));
   INV_X1 i_69 (.A(a[20]), .ZN(n_64));
   INV_X1 i_70 (.A(a[21]), .ZN(n_65));
   INV_X1 i_71 (.A(n_66), .ZN(p_0[23]));
   NAND2_X1 i_72 (.A1(n_83), .A2(n_67), .ZN(n_66));
   NAND2_X1 i_73 (.A1(n_85), .A2(a[23]), .ZN(n_67));
   INV_X1 i_74 (.A(n_68), .ZN(p_0[24]));
   XNOR2_X1 i_75 (.A(n_83), .B(a[24]), .ZN(n_68));
   AND2_X1 i_76 (.A1(n_69), .A2(n_70), .ZN(p_0[25]));
   OAI21_X1 i_77 (.A(a[25]), .B1(n_83), .B2(a[24]), .ZN(n_69));
   AOI22_X1 i_78 (.A1(n_70), .A2(a[26]), .B1(n_82), .B2(n_72), .ZN(p_0[26]));
   NAND3_X1 i_79 (.A1(n_82), .A2(n_80), .A3(n_79), .ZN(n_70));
   AOI21_X1 i_80 (.A(n_75), .B1(n_71), .B2(a[27]), .ZN(p_0[27]));
   NAND2_X1 i_81 (.A1(n_82), .A2(n_72), .ZN(n_71));
   INV_X1 i_82 (.A(n_78), .ZN(n_72));
   XNOR2_X1 i_83 (.A(n_38), .B(n_101), .ZN(p_0[28]));
   INV_X1 i_84 (.A(n_73), .ZN(p_0[29]));
   XNOR2_X1 i_85 (.A(n_74), .B(a[29]), .ZN(n_73));
   NAND2_X1 i_86 (.A1(n_75), .A2(n_101), .ZN(n_74));
   INV_X1 i_87 (.A(n_38), .ZN(n_75));
   NAND2_X1 i_88 (.A1(n_82), .A2(n_76), .ZN(n_38));
   INV_X1 i_89 (.A(n_77), .ZN(n_76));
   OR2_X1 i_90 (.A1(n_78), .A2(a[27]), .ZN(n_77));
   NAND3_X1 i_91 (.A1(n_81), .A2(n_80), .A3(n_79), .ZN(n_78));
   INV_X1 i_92 (.A(a[24]), .ZN(n_79));
   INV_X1 i_93 (.A(a[25]), .ZN(n_80));
   INV_X1 i_94 (.A(a[26]), .ZN(n_81));
   INV_X1 i_95 (.A(n_83), .ZN(n_82));
   NAND2_X1 i_96 (.A1(n_84), .A2(n_100), .ZN(n_83));
   INV_X1 i_97 (.A(n_85), .ZN(n_84));
   NAND2_X1 i_98 (.A1(n_45), .A2(n_86), .ZN(n_85));
   INV_X1 i_99 (.A(n_87), .ZN(n_86));
   OR3_X1 i_100 (.A1(a[22]), .A2(a[21]), .A3(a[20]), .ZN(n_87));
   INV_X1 i_101 (.A(n_44), .ZN(n_45));
   NAND2_X1 i_102 (.A1(n_49), .A2(n_88), .ZN(n_44));
   INV_X1 i_103 (.A(n_89), .ZN(n_88));
   OR2_X1 i_104 (.A1(n_46), .A2(a[19]), .ZN(n_89));
   OR3_X1 i_105 (.A1(a[18]), .A2(a[17]), .A3(a[16]), .ZN(n_46));
   INV_X1 i_106 (.A(n_48), .ZN(n_49));
   NAND2_X1 i_107 (.A1(n_52), .A2(n_90), .ZN(n_48));
   INV_X1 i_108 (.A(n_91), .ZN(n_90));
   OR2_X1 i_109 (.A1(n_50), .A2(a[15]), .ZN(n_91));
   OR3_X1 i_110 (.A1(a[14]), .A2(a[13]), .A3(a[12]), .ZN(n_50));
   INV_X1 i_111 (.A(n_51), .ZN(n_52));
   NAND2_X1 i_112 (.A1(n_55), .A2(n_92), .ZN(n_51));
   INV_X1 i_113 (.A(n_93), .ZN(n_92));
   OR2_X1 i_114 (.A1(n_53), .A2(a[11]), .ZN(n_93));
   OR3_X1 i_115 (.A1(a[10]), .A2(a[9]), .A3(a[8]), .ZN(n_53));
   INV_X1 i_116 (.A(n_54), .ZN(n_55));
   NAND2_X1 i_117 (.A1(n_94), .A2(n_58), .ZN(n_54));
   INV_X1 i_118 (.A(n_95), .ZN(n_94));
   OR2_X1 i_119 (.A1(n_56), .A2(a[7]), .ZN(n_95));
   OR3_X1 i_120 (.A1(a[6]), .A2(a[5]), .A3(a[4]), .ZN(n_56));
   INV_X1 i_121 (.A(n_57), .ZN(n_58));
   NAND2_X1 i_122 (.A1(n_60), .A2(n_99), .ZN(n_57));
   INV_X1 i_123 (.A(n_59), .ZN(n_60));
   NAND2_X1 i_124 (.A1(n_62), .A2(n_98), .ZN(n_59));
   INV_X1 i_125 (.A(n_61), .ZN(n_62));
   NAND2_X1 i_126 (.A1(n_97), .A2(n_96), .ZN(n_61));
   INV_X1 i_127 (.A(a[0]), .ZN(n_96));
   INV_X1 i_128 (.A(a[1]), .ZN(n_97));
   INV_X1 i_129 (.A(a[2]), .ZN(n_98));
   INV_X1 i_130 (.A(a[3]), .ZN(n_99));
   INV_X1 i_131 (.A(a[23]), .ZN(n_100));
   INV_X1 i_132 (.A(a[28]), .ZN(n_101));
endmodule

module datapath__0_65(A, p_0, multiplicand);
   input [31:0]A;
   output [31:0]p_0;
   input [31:0]multiplicand;

   OAI21_X1 i_0 (.A(n_102), .B1(n_123), .B2(multiplicand[0]), .ZN(p_0[0]));
   XNOR2_X1 i_1 (.A(n_101), .B(n_0), .ZN(p_0[1]));
   NOR2_X1 i_2 (.A1(n_111), .A2(n_104), .ZN(n_0));
   XOR2_X1 i_3 (.A(n_3), .B(n_1), .Z(p_0[2]));
   NOR2_X1 i_4 (.A1(n_109), .A2(n_100), .ZN(n_1));
   XOR2_X1 i_5 (.A(n_4), .B(n_2), .Z(p_0[3]));
   OAI21_X1 i_6 (.A(n_110), .B1(n_100), .B2(n_3), .ZN(n_2));
   OAI22_X1 i_7 (.A1(n_124), .A2(multiplicand[1]), .B1(n_111), .B2(n_101), 
      .ZN(n_3));
   OAI21_X1 i_8 (.A(n_108), .B1(n_126), .B2(multiplicand[3]), .ZN(n_4));
   XNOR2_X1 i_9 (.A(n_97), .B(n_5), .ZN(p_0[4]));
   NOR2_X1 i_10 (.A1(n_112), .A2(n_96), .ZN(n_5));
   XNOR2_X1 i_11 (.A(n_11), .B(n_6), .ZN(p_0[5]));
   OAI21_X1 i_12 (.A(n_115), .B1(n_128), .B2(multiplicand[5]), .ZN(n_6));
   XNOR2_X1 i_13 (.A(n_9), .B(n_7), .ZN(p_0[6]));
   OAI21_X1 i_14 (.A(n_116), .B1(n_129), .B2(multiplicand[6]), .ZN(n_7));
   XOR2_X1 i_15 (.A(n_12), .B(n_8), .Z(p_0[7]));
   OAI21_X1 i_16 (.A(n_116), .B1(n_93), .B2(n_9), .ZN(n_8));
   INV_X1 i_17 (.A(n_10), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_115), .B1(n_95), .B2(n_11), .ZN(n_10));
   OAI22_X1 i_19 (.A1(n_112), .A2(n_97), .B1(n_127), .B2(multiplicand[4]), 
      .ZN(n_11));
   OAI21_X1 i_20 (.A(n_114), .B1(n_130), .B2(multiplicand[7]), .ZN(n_12));
   XNOR2_X1 i_21 (.A(n_28), .B(n_13), .ZN(p_0[8]));
   NOR2_X1 i_22 (.A1(n_118), .A2(n_229), .ZN(n_13));
   XOR2_X1 i_23 (.A(n_18), .B(n_14), .Z(p_0[9]));
   NOR2_X1 i_24 (.A1(n_161), .A2(n_227), .ZN(n_14));
   XNOR2_X1 i_25 (.A(n_17), .B(n_15), .ZN(p_0[10]));
   NOR2_X1 i_26 (.A1(n_224), .A2(n_218), .ZN(n_15));
   XNOR2_X1 i_27 (.A(n_19), .B(n_16), .ZN(p_0[11]));
   OAI21_X1 i_28 (.A(n_160), .B1(n_224), .B2(n_17), .ZN(n_16));
   OAI21_X1 i_29 (.A(n_223), .B1(n_227), .B2(n_18), .ZN(n_17));
   OAI22_X1 i_30 (.A1(n_131), .A2(multiplicand[8]), .B1(n_118), .B2(n_28), 
      .ZN(n_18));
   OAI21_X1 i_31 (.A(n_222), .B1(n_230), .B2(multiplicand[11]), .ZN(n_19));
   XNOR2_X1 i_32 (.A(n_27), .B(n_20), .ZN(p_0[12]));
   OAI21_X1 i_33 (.A(n_213), .B1(n_132), .B2(multiplicand[12]), .ZN(n_20));
   XNOR2_X1 i_34 (.A(n_26), .B(n_21), .ZN(p_0[13]));
   NOR2_X1 i_35 (.A1(n_159), .A2(n_202), .ZN(n_21));
   XNOR2_X1 i_36 (.A(n_24), .B(n_22), .ZN(p_0[14]));
   NOR2_X1 i_37 (.A1(n_158), .A2(n_200), .ZN(n_22));
   XNOR2_X1 i_38 (.A(n_29), .B(n_23), .ZN(p_0[15]));
   OAI21_X1 i_39 (.A(n_157), .B1(n_158), .B2(n_24), .ZN(n_23));
   OAI21_X1 i_40 (.A(n_209), .B1(n_202), .B2(n_25), .ZN(n_24));
   INV_X1 i_41 (.A(n_26), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_213), .B1(n_203), .B2(n_27), .ZN(n_26));
   OAI21_X1 i_43 (.A(n_215), .B1(n_117), .B2(n_28), .ZN(n_27));
   NOR2_X1 i_44 (.A1(n_234), .A2(n_233), .ZN(n_28));
   OAI21_X1 i_45 (.A(n_207), .B1(n_208), .B2(multiplicand[15]), .ZN(n_29));
   XNOR2_X1 i_46 (.A(n_156), .B(n_30), .ZN(p_0[16]));
   NOR2_X1 i_47 (.A1(n_155), .A2(n_88), .ZN(n_30));
   INV_X1 i_48 (.A(n_31), .ZN(p_0[17]));
   AOI21_X1 i_49 (.A(n_35), .B1(n_37), .B2(n_36), .ZN(n_31));
   XNOR2_X1 i_50 (.A(n_33), .B(n_32), .ZN(p_0[18]));
   OAI21_X1 i_51 (.A(n_91), .B1(n_87), .B2(n_37), .ZN(n_32));
   NOR2_X1 i_52 (.A1(n_89), .A2(n_85), .ZN(n_33));
   XOR2_X1 i_53 (.A(n_38), .B(n_34), .Z(p_0[19]));
   OAI21_X1 i_54 (.A(n_84), .B1(n_154), .B2(n_35), .ZN(n_34));
   NOR2_X1 i_55 (.A1(n_37), .A2(n_36), .ZN(n_35));
   OR2_X1 i_56 (.A1(n_90), .A2(n_87), .ZN(n_36));
   OAI22_X1 i_57 (.A1(n_133), .A2(multiplicand[16]), .B1(n_156), .B2(n_155), 
      .ZN(n_37));
   NOR2_X1 i_58 (.A1(n_240), .A2(n_153), .ZN(n_38));
   XOR2_X1 i_59 (.A(n_152), .B(n_39), .Z(p_0[20]));
   OAI22_X1 i_60 (.A1(A[20]), .A2(n_120), .B1(n_137), .B2(multiplicand[20]), 
      .ZN(n_39));
   INV_X1 i_61 (.A(n_40), .ZN(p_0[21]));
   AOI21_X1 i_62 (.A(n_44), .B1(n_46), .B2(n_45), .ZN(n_40));
   XNOR2_X1 i_63 (.A(n_42), .B(n_41), .ZN(p_0[22]));
   OAI21_X1 i_64 (.A(n_83), .B1(n_80), .B2(n_46), .ZN(n_41));
   NOR2_X1 i_65 (.A1(n_81), .A2(n_78), .ZN(n_42));
   XOR2_X1 i_66 (.A(n_47), .B(n_43), .Z(p_0[23]));
   OAI21_X1 i_67 (.A(n_77), .B1(n_185), .B2(n_44), .ZN(n_43));
   NOR2_X1 i_68 (.A1(n_46), .A2(n_45), .ZN(n_44));
   OR2_X1 i_69 (.A1(n_82), .A2(n_80), .ZN(n_45));
   OAI22_X1 i_70 (.A1(n_137), .A2(multiplicand[20]), .B1(n_152), .B2(n_151), 
      .ZN(n_46));
   NOR2_X1 i_71 (.A1(n_150), .A2(n_149), .ZN(n_47));
   XOR2_X1 i_72 (.A(n_148), .B(n_48), .Z(p_0[24]));
   OAI22_X1 i_73 (.A1(A[24]), .A2(n_121), .B1(n_141), .B2(multiplicand[24]), 
      .ZN(n_48));
   INV_X1 i_74 (.A(n_49), .ZN(p_0[25]));
   AOI21_X1 i_75 (.A(n_53), .B1(n_55), .B2(n_54), .ZN(n_49));
   XNOR2_X1 i_76 (.A(n_51), .B(n_50), .ZN(p_0[26]));
   OAI21_X1 i_77 (.A(n_76), .B1(n_73), .B2(n_55), .ZN(n_50));
   NOR2_X1 i_78 (.A1(n_74), .A2(n_71), .ZN(n_51));
   XOR2_X1 i_79 (.A(n_56), .B(n_52), .Z(p_0[27]));
   OAI21_X1 i_80 (.A(n_70), .B1(n_172), .B2(n_53), .ZN(n_52));
   NOR2_X1 i_81 (.A1(n_55), .A2(n_54), .ZN(n_53));
   OR2_X1 i_82 (.A1(n_75), .A2(n_73), .ZN(n_54));
   OAI22_X1 i_83 (.A1(n_141), .A2(multiplicand[24]), .B1(n_148), .B2(n_179), 
      .ZN(n_55));
   NOR2_X1 i_84 (.A1(n_147), .A2(n_146), .ZN(n_56));
   XOR2_X1 i_85 (.A(n_68), .B(n_63), .Z(p_0[29]));
   XNOR2_X1 i_86 (.A(n_58), .B(n_57), .ZN(p_0[30]));
   OAI22_X1 i_87 (.A1(n_145), .A2(multiplicand[29]), .B1(n_68), .B2(n_64), 
      .ZN(n_57));
   OAI21_X1 i_88 (.A(n_67), .B1(A[31]), .B2(n_122), .ZN(n_58));
   XOR2_X1 i_89 (.A(n_60), .B(n_59), .Z(p_0[31]));
   XOR2_X1 i_90 (.A(A[31]), .B(multiplicand[31]), .Z(n_59));
   OAI221_X1 i_91 (.A(n_61), .B1(A[31]), .B2(n_122), .C1(n_66), .C2(n_65), 
      .ZN(n_60));
   NAND3_X1 i_92 (.A1(n_67), .A2(n_62), .A3(n_68), .ZN(n_61));
   INV_X1 i_93 (.A(n_63), .ZN(n_62));
   OAI21_X1 i_94 (.A(n_65), .B1(n_145), .B2(multiplicand[29]), .ZN(n_63));
   INV_X1 i_95 (.A(n_65), .ZN(n_64));
   NAND2_X1 i_96 (.A1(n_145), .A2(multiplicand[29]), .ZN(n_65));
   INV_X1 i_97 (.A(n_67), .ZN(n_66));
   NAND2_X1 i_98 (.A1(A[31]), .A2(n_122), .ZN(n_67));
   OAI21_X1 i_99 (.A(n_69), .B1(A[28]), .B2(n_164), .ZN(n_68));
   NAND2_X1 i_100 (.A1(multiplicand[28]), .A2(n_163), .ZN(n_69));
   INV_X1 i_101 (.A(n_71), .ZN(n_70));
   NOR2_X1 i_102 (.A1(n_143), .A2(multiplicand[26]), .ZN(n_71));
   AOI21_X1 i_103 (.A(n_73), .B1(A[24]), .B2(n_121), .ZN(n_72));
   NOR2_X1 i_104 (.A1(n_142), .A2(multiplicand[25]), .ZN(n_73));
   AND2_X1 i_105 (.A1(n_143), .A2(multiplicand[26]), .ZN(n_74));
   INV_X1 i_106 (.A(n_76), .ZN(n_75));
   NAND2_X1 i_107 (.A1(n_142), .A2(multiplicand[25]), .ZN(n_76));
   INV_X1 i_108 (.A(n_78), .ZN(n_77));
   NOR2_X1 i_109 (.A1(n_139), .A2(multiplicand[22]), .ZN(n_78));
   AOI21_X1 i_110 (.A(n_80), .B1(A[20]), .B2(n_120), .ZN(n_79));
   NOR2_X1 i_111 (.A1(n_138), .A2(multiplicand[21]), .ZN(n_80));
   AND2_X1 i_112 (.A1(n_139), .A2(multiplicand[22]), .ZN(n_81));
   INV_X1 i_113 (.A(n_83), .ZN(n_82));
   NAND2_X1 i_114 (.A1(n_138), .A2(multiplicand[21]), .ZN(n_83));
   INV_X1 i_115 (.A(n_85), .ZN(n_84));
   NOR2_X1 i_116 (.A1(n_135), .A2(multiplicand[18]), .ZN(n_85));
   NOR2_X1 i_117 (.A1(n_88), .A2(n_87), .ZN(n_86));
   NOR2_X1 i_118 (.A1(n_134), .A2(multiplicand[17]), .ZN(n_87));
   NOR2_X1 i_119 (.A1(n_133), .A2(multiplicand[16]), .ZN(n_88));
   AND2_X1 i_120 (.A1(n_135), .A2(multiplicand[18]), .ZN(n_89));
   INV_X1 i_121 (.A(n_91), .ZN(n_90));
   NAND2_X1 i_122 (.A1(n_134), .A2(multiplicand[17]), .ZN(n_91));
   NAND2_X1 i_123 (.A1(n_114), .A2(n_93), .ZN(n_92));
   NOR2_X1 i_124 (.A1(n_129), .A2(multiplicand[6]), .ZN(n_93));
   NOR2_X1 i_125 (.A1(n_96), .A2(n_95), .ZN(n_94));
   NOR2_X1 i_126 (.A1(n_128), .A2(multiplicand[5]), .ZN(n_95));
   NOR2_X1 i_127 (.A1(n_127), .A2(multiplicand[4]), .ZN(n_96));
   AOI21_X1 i_128 (.A(n_98), .B1(n_106), .B2(n_102), .ZN(n_97));
   OAI221_X1 i_129 (.A(n_103), .B1(n_107), .B2(n_99), .C1(n_126), .C2(
      multiplicand[3]), .ZN(n_98));
   INV_X1 i_130 (.A(n_100), .ZN(n_99));
   NOR2_X1 i_131 (.A1(n_125), .A2(multiplicand[2]), .ZN(n_100));
   INV_X1 i_132 (.A(n_102), .ZN(n_101));
   NAND2_X1 i_133 (.A1(n_123), .A2(multiplicand[0]), .ZN(n_102));
   OAI21_X1 i_134 (.A(n_106), .B1(n_105), .B2(n_104), .ZN(n_103));
   NOR2_X1 i_135 (.A1(n_124), .A2(multiplicand[1]), .ZN(n_104));
   NOR2_X1 i_136 (.A1(n_123), .A2(multiplicand[0]), .ZN(n_105));
   NOR3_X1 i_137 (.A1(n_111), .A2(n_107), .A3(n_109), .ZN(n_106));
   INV_X1 i_138 (.A(n_108), .ZN(n_107));
   NAND2_X1 i_139 (.A1(n_126), .A2(multiplicand[3]), .ZN(n_108));
   INV_X1 i_140 (.A(n_110), .ZN(n_109));
   NAND2_X1 i_141 (.A1(n_125), .A2(multiplicand[2]), .ZN(n_110));
   AND2_X1 i_142 (.A1(n_124), .A2(multiplicand[1]), .ZN(n_111));
   AND2_X1 i_143 (.A1(n_127), .A2(multiplicand[4]), .ZN(n_112));
   NAND3_X1 i_144 (.A1(n_116), .A2(n_114), .A3(n_115), .ZN(n_113));
   NAND2_X1 i_145 (.A1(n_130), .A2(multiplicand[7]), .ZN(n_114));
   NAND2_X1 i_146 (.A1(n_128), .A2(multiplicand[5]), .ZN(n_115));
   NAND2_X1 i_147 (.A1(n_129), .A2(multiplicand[6]), .ZN(n_116));
   NAND2_X1 i_148 (.A1(n_220), .A2(n_119), .ZN(n_117));
   INV_X1 i_149 (.A(n_119), .ZN(n_118));
   NAND2_X1 i_150 (.A1(n_131), .A2(multiplicand[8]), .ZN(n_119));
   INV_X1 i_151 (.A(multiplicand[20]), .ZN(n_120));
   INV_X1 i_152 (.A(multiplicand[24]), .ZN(n_121));
   INV_X1 i_153 (.A(multiplicand[30]), .ZN(n_122));
   INV_X1 i_154 (.A(A[0]), .ZN(n_123));
   INV_X1 i_155 (.A(A[1]), .ZN(n_124));
   INV_X1 i_156 (.A(A[2]), .ZN(n_125));
   INV_X1 i_157 (.A(A[3]), .ZN(n_126));
   INV_X1 i_158 (.A(A[4]), .ZN(n_127));
   INV_X1 i_159 (.A(A[5]), .ZN(n_128));
   INV_X1 i_160 (.A(A[6]), .ZN(n_129));
   INV_X1 i_161 (.A(A[7]), .ZN(n_130));
   INV_X1 i_162 (.A(A[8]), .ZN(n_131));
   INV_X1 i_163 (.A(A[12]), .ZN(n_132));
   INV_X1 i_164 (.A(A[16]), .ZN(n_133));
   INV_X1 i_165 (.A(A[17]), .ZN(n_134));
   INV_X1 i_166 (.A(A[18]), .ZN(n_135));
   INV_X1 i_167 (.A(A[19]), .ZN(n_136));
   INV_X1 i_168 (.A(A[20]), .ZN(n_137));
   INV_X1 i_169 (.A(A[21]), .ZN(n_138));
   INV_X1 i_170 (.A(A[22]), .ZN(n_139));
   INV_X1 i_171 (.A(A[23]), .ZN(n_140));
   INV_X1 i_172 (.A(A[24]), .ZN(n_141));
   INV_X1 i_173 (.A(A[25]), .ZN(n_142));
   INV_X1 i_174 (.A(A[26]), .ZN(n_143));
   INV_X1 i_175 (.A(A[27]), .ZN(n_144));
   INV_X1 i_176 (.A(A[29]), .ZN(n_145));
   NOR2_X1 i_177 (.A1(multiplicand[27]), .A2(n_144), .ZN(n_146));
   INV_X1 i_178 (.A(n_176), .ZN(n_147));
   INV_X1 i_179 (.A(n_180), .ZN(n_148));
   NOR2_X1 i_180 (.A1(multiplicand[23]), .A2(n_140), .ZN(n_149));
   INV_X1 i_181 (.A(n_190), .ZN(n_150));
   NOR2_X1 i_182 (.A1(n_120), .A2(A[20]), .ZN(n_151));
   NOR2_X1 i_183 (.A1(n_235), .A2(n_191), .ZN(n_152));
   NOR2_X1 i_184 (.A1(multiplicand[19]), .A2(n_136), .ZN(n_153));
   NAND2_X1 i_185 (.A1(n_238), .A2(n_239), .ZN(n_154));
   INV_X1 i_186 (.A(n_195), .ZN(n_155));
   INV_X1 i_187 (.A(n_196), .ZN(n_156));
   INV_X1 i_188 (.A(n_200), .ZN(n_157));
   INV_X1 i_189 (.A(n_211), .ZN(n_158));
   INV_X1 i_190 (.A(n_209), .ZN(n_159));
   INV_X1 i_191 (.A(n_218), .ZN(n_160));
   INV_X1 i_192 (.A(n_223), .ZN(n_161));
   NAND2_X1 i_193 (.A1(n_165), .A2(n_162), .ZN(p_0[28]));
   NAND3_X1 i_194 (.A1(n_163), .A2(multiplicand[28]), .A3(n_167), .ZN(n_162));
   NAND2_X1 i_195 (.A1(n_164), .A2(A[28]), .ZN(n_163));
   NAND2_X1 i_196 (.A1(n_173), .A2(n_169), .ZN(n_164));
   OAI21_X1 i_197 (.A(n_243), .B1(n_166), .B2(n_168), .ZN(n_165));
   INV_X1 i_198 (.A(n_167), .ZN(n_166));
   NAND3_X1 i_199 (.A1(n_173), .A2(n_242), .A3(n_169), .ZN(n_167));
   AOI21_X1 i_200 (.A(n_242), .B1(n_173), .B2(n_169), .ZN(n_168));
   OAI21_X1 i_201 (.A(n_176), .B1(n_171), .B2(n_170), .ZN(n_169));
   OAI21_X1 i_202 (.A(n_70), .B1(multiplicand[27]), .B2(n_144), .ZN(n_170));
   NOR2_X1 i_203 (.A1(n_172), .A2(n_72), .ZN(n_171));
   NAND2_X1 i_204 (.A1(n_177), .A2(n_178), .ZN(n_172));
   NAND2_X1 i_205 (.A1(n_180), .A2(n_174), .ZN(n_173));
   NOR2_X1 i_206 (.A1(n_175), .A2(n_179), .ZN(n_174));
   NAND3_X1 i_207 (.A1(n_177), .A2(n_178), .A3(n_176), .ZN(n_175));
   NAND2_X1 i_208 (.A1(multiplicand[27]), .A2(n_144), .ZN(n_176));
   INV_X1 i_209 (.A(n_75), .ZN(n_177));
   INV_X1 i_210 (.A(n_74), .ZN(n_178));
   NOR2_X1 i_211 (.A1(n_121), .A2(A[24]), .ZN(n_179));
   NAND2_X1 i_212 (.A1(n_186), .A2(n_181), .ZN(n_180));
   OAI21_X1 i_213 (.A(n_190), .B1(n_183), .B2(n_182), .ZN(n_181));
   OAI21_X1 i_214 (.A(n_77), .B1(multiplicand[23]), .B2(n_140), .ZN(n_182));
   INV_X1 i_215 (.A(n_184), .ZN(n_183));
   OR2_X1 i_216 (.A1(n_185), .A2(n_79), .ZN(n_184));
   INV_X1 i_217 (.A(n_189), .ZN(n_185));
   OAI21_X1 i_218 (.A(n_187), .B1(n_235), .B2(n_191), .ZN(n_186));
   INV_X1 i_219 (.A(n_188), .ZN(n_187));
   OAI211_X1 i_220 (.A(n_190), .B(n_189), .C1(A[20]), .C2(n_120), .ZN(n_188));
   NOR2_X1 i_221 (.A1(n_82), .A2(n_81), .ZN(n_189));
   NAND2_X1 i_222 (.A1(multiplicand[23]), .A2(n_140), .ZN(n_190));
   OAI21_X1 i_223 (.A(n_192), .B1(multiplicand[19]), .B2(n_136), .ZN(n_191));
   NAND3_X1 i_224 (.A1(n_238), .A2(n_193), .A3(n_239), .ZN(n_192));
   INV_X1 i_225 (.A(n_194), .ZN(n_193));
   NAND3_X1 i_226 (.A1(n_196), .A2(n_241), .A3(n_195), .ZN(n_194));
   NAND2_X1 i_227 (.A1(multiplicand[16]), .A2(n_133), .ZN(n_195));
   NAND2_X1 i_228 (.A1(n_204), .A2(n_197), .ZN(n_196));
   INV_X1 i_229 (.A(n_198), .ZN(n_197));
   OAI211_X1 i_230 (.A(n_201), .B(n_199), .C1(n_208), .C2(multiplicand[15]), 
      .ZN(n_198));
   NAND2_X1 i_231 (.A1(n_200), .A2(n_207), .ZN(n_199));
   NOR2_X1 i_232 (.A1(multiplicand[14]), .A2(n_212), .ZN(n_200));
   OAI211_X1 i_233 (.A(n_211), .B(n_205), .C1(n_203), .C2(n_202), .ZN(n_201));
   NOR2_X1 i_234 (.A1(multiplicand[13]), .A2(n_210), .ZN(n_202));
   NOR2_X1 i_235 (.A1(multiplicand[12]), .A2(n_132), .ZN(n_203));
   NAND4_X1 i_236 (.A1(n_214), .A2(n_213), .A3(n_211), .A4(n_205), .ZN(n_204));
   INV_X1 i_237 (.A(n_206), .ZN(n_205));
   NAND2_X1 i_238 (.A1(n_209), .A2(n_207), .ZN(n_206));
   NAND2_X1 i_239 (.A1(multiplicand[15]), .A2(n_208), .ZN(n_207));
   INV_X1 i_240 (.A(A[15]), .ZN(n_208));
   NAND2_X1 i_241 (.A1(multiplicand[13]), .A2(n_210), .ZN(n_209));
   INV_X1 i_242 (.A(A[13]), .ZN(n_210));
   NAND2_X1 i_243 (.A1(multiplicand[14]), .A2(n_212), .ZN(n_211));
   INV_X1 i_244 (.A(A[14]), .ZN(n_212));
   NAND2_X1 i_245 (.A1(multiplicand[12]), .A2(n_132), .ZN(n_213));
   OAI21_X1 i_246 (.A(n_215), .B1(n_117), .B2(n_231), .ZN(n_214));
   INV_X1 i_247 (.A(n_216), .ZN(n_215));
   OAI211_X1 i_248 (.A(n_219), .B(n_217), .C1(n_230), .C2(multiplicand[11]), 
      .ZN(n_216));
   NAND2_X1 i_249 (.A1(n_218), .A2(n_222), .ZN(n_217));
   NOR2_X1 i_250 (.A1(multiplicand[10]), .A2(n_226), .ZN(n_218));
   OAI21_X1 i_251 (.A(n_220), .B1(n_229), .B2(n_227), .ZN(n_219));
   NOR2_X1 i_252 (.A1(n_224), .A2(n_221), .ZN(n_220));
   NAND2_X1 i_253 (.A1(n_223), .A2(n_222), .ZN(n_221));
   NAND2_X1 i_254 (.A1(multiplicand[11]), .A2(n_230), .ZN(n_222));
   NAND2_X1 i_255 (.A1(multiplicand[9]), .A2(n_228), .ZN(n_223));
   INV_X1 i_256 (.A(n_225), .ZN(n_224));
   NAND2_X1 i_257 (.A1(multiplicand[10]), .A2(n_226), .ZN(n_225));
   INV_X1 i_258 (.A(A[10]), .ZN(n_226));
   NOR2_X1 i_259 (.A1(multiplicand[9]), .A2(n_228), .ZN(n_227));
   INV_X1 i_260 (.A(A[9]), .ZN(n_228));
   NOR2_X1 i_261 (.A1(multiplicand[8]), .A2(n_131), .ZN(n_229));
   INV_X1 i_262 (.A(A[11]), .ZN(n_230));
   INV_X1 i_263 (.A(n_232), .ZN(n_231));
   OR2_X1 i_264 (.A1(n_233), .A2(n_234), .ZN(n_232));
   OAI221_X1 i_265 (.A(n_92), .B1(multiplicand[7]), .B2(n_130), .C1(n_113), 
      .C2(n_94), .ZN(n_233));
   NOR3_X1 i_266 (.A1(n_97), .A2(n_112), .A3(n_113), .ZN(n_234));
   AOI21_X1 i_267 (.A(n_240), .B1(n_236), .B2(n_84), .ZN(n_235));
   NAND3_X1 i_268 (.A1(n_237), .A2(n_239), .A3(n_238), .ZN(n_236));
   INV_X1 i_269 (.A(n_86), .ZN(n_237));
   INV_X1 i_270 (.A(n_90), .ZN(n_238));
   INV_X1 i_271 (.A(n_89), .ZN(n_239));
   INV_X1 i_272 (.A(n_241), .ZN(n_240));
   NAND2_X1 i_273 (.A1(multiplicand[19]), .A2(n_136), .ZN(n_241));
   INV_X1 i_274 (.A(A[28]), .ZN(n_242));
   INV_X1 i_275 (.A(multiplicand[28]), .ZN(n_243));
endmodule

module datapath__0_66(multiplicand, A, p_0);
   input [31:0]multiplicand;
   input [31:0]A;
   output [31:0]p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0[0]));
   OAI21_X1 i_1 (.A(n_154), .B1(multiplicand[0]), .B2(A[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_154), .B(n_1), .Z(p_0[1]));
   OAI21_X1 i_3 (.A(n_153), .B1(multiplicand[1]), .B2(A[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_152), .B(n_2), .ZN(p_0[2]));
   OAI21_X1 i_5 (.A(n_157), .B1(multiplicand[2]), .B2(A[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_151), .B(n_3), .Z(p_0[3]));
   OAI21_X1 i_7 (.A(n_158), .B1(n_164), .B2(n_161), .ZN(n_3));
   XOR2_X1 i_8 (.A(n_149), .B(n_10), .Z(p_0[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_0[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_0[6]));
   NOR2_X1 i_11 (.A1(n_146), .A2(n_137), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_0[7]));
   OAI22_X1 i_13 (.A1(multiplicand[6]), .A2(A[6]), .B1(n_137), .B2(n_7), 
      .ZN(n_5));
   AOI21_X1 i_14 (.A(n_147), .B1(multiplicand[5]), .B2(A[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_147), .B1(n_141), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_144), .B1(n_149), .B2(n_142), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_142), .B1(multiplicand[4]), .B2(A[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_148), .A2(n_139), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_135), .B(n_18), .ZN(p_0[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_0[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_0[10]));
   NOR2_X1 i_23 (.A1(n_132), .A2(n_123), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_0[11]));
   OAI22_X1 i_25 (.A1(multiplicand[10]), .A2(A[10]), .B1(n_123), .B2(n_15), 
      .ZN(n_13));
   AOI21_X1 i_26 (.A(n_133), .B1(multiplicand[9]), .B2(A[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_133), .B1(n_127), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_130), .B1(n_135), .B2(n_128), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_130), .B1(multiplicand[8]), .B2(A[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_134), .A2(n_125), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_121), .B(n_26), .Z(p_0[12]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(p_0[13]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(p_0[14]));
   NOR2_X1 i_35 (.A1(n_118), .A2(n_109), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(p_0[15]));
   OAI22_X1 i_37 (.A1(multiplicand[14]), .A2(A[14]), .B1(n_109), .B2(n_23), 
      .ZN(n_21));
   AOI21_X1 i_38 (.A(n_119), .B1(multiplicand[13]), .B2(A[13]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_119), .B1(n_113), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_116), .B1(n_121), .B2(n_114), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_114), .B1(multiplicand[12]), .B2(A[12]), .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_120), .A2(n_111), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_107), .B(n_34), .Z(p_0[16]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(p_0[17]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(p_0[18]));
   NOR2_X1 i_47 (.A1(n_104), .A2(n_95), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(p_0[19]));
   OAI22_X1 i_49 (.A1(multiplicand[18]), .A2(A[18]), .B1(n_95), .B2(n_31), 
      .ZN(n_29));
   AOI21_X1 i_50 (.A(n_105), .B1(multiplicand[17]), .B2(A[17]), .ZN(n_30));
   AOI21_X1 i_51 (.A(n_105), .B1(n_99), .B2(n_32), .ZN(n_31));
   INV_X1 i_52 (.A(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_102), .B1(n_107), .B2(n_100), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_100), .B1(multiplicand[16]), .B2(A[16]), .ZN(n_34));
   NOR2_X1 i_55 (.A1(n_106), .A2(n_97), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_93), .B(n_42), .Z(p_0[20]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(p_0[21]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(p_0[22]));
   NOR2_X1 i_59 (.A1(n_82), .A2(n_72), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(p_0[23]));
   OAI21_X1 i_61 (.A(n_81), .B1(n_72), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_84), .A2(n_74), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_83), .B1(n_74), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_79), .B1(n_93), .B2(n_76), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_76), .B1(multiplicand[20]), .B2(A[20]), .ZN(n_42));
   AOI21_X1 i_67 (.A(n_86), .B1(multiplicand[23]), .B2(A[23]), .ZN(n_43));
   XOR2_X1 i_68 (.A(n_51), .B(n_50), .Z(p_0[24]));
   OAI21_X1 i_78 (.A(n_69), .B1(multiplicand[24]), .B2(A[24]), .ZN(n_50));
   XNOR2_X1 i_82 (.A(n_64), .B(n_63), .ZN(p_0[28]));
   XOR2_X1 i_83 (.A(n_62), .B(n_58), .Z(p_0[29]));
   XNOR2_X1 i_84 (.A(n_55), .B(n_54), .ZN(p_0[30]));
   OAI21_X1 i_85 (.A(n_160), .B1(n_166), .B2(n_163), .ZN(n_54));
   NOR2_X1 i_86 (.A1(n_61), .A2(n_60), .ZN(n_55));
   XOR2_X1 i_87 (.A(n_57), .B(n_56), .Z(p_0[31]));
   XNOR2_X1 i_88 (.A(multiplicand[31]), .B(multiplicand[30]), .ZN(n_56));
   OAI21_X1 i_89 (.A(n_160), .B1(n_61), .B2(n_59), .ZN(n_57));
   AOI21_X1 i_90 (.A(n_60), .B1(multiplicand[29]), .B2(A[29]), .ZN(n_58));
   OAI22_X1 i_91 (.A1(n_166), .A2(n_163), .B1(multiplicand[29]), .B2(A[29]), 
      .ZN(n_59));
   NOR2_X1 i_92 (.A1(multiplicand[29]), .A2(A[29]), .ZN(n_60));
   AOI21_X1 i_93 (.A(n_62), .B1(multiplicand[29]), .B2(A[29]), .ZN(n_61));
   AOI21_X1 i_94 (.A(n_159), .B1(n_64), .B2(n_63), .ZN(n_62));
   AOI21_X1 i_95 (.A(n_159), .B1(multiplicand[28]), .B2(A[28]), .ZN(n_63));
   NOR4_X1 i_96 (.A1(n_67), .A2(n_65), .A3(n_70), .A4(n_77), .ZN(n_64));
   OAI22_X1 i_97 (.A1(n_165), .A2(n_162), .B1(n_92), .B2(n_66), .ZN(n_65));
   AOI21_X1 i_99 (.A(n_89), .B1(n_69), .B2(n_68), .ZN(n_67));
   NAND2_X1 i_100 (.A1(multiplicand[25]), .A2(A[25]), .ZN(n_68));
   NOR2_X1 i_102 (.A1(n_87), .A2(n_71), .ZN(n_70));
   INV_X1 i_106 (.A(n_75), .ZN(n_74));
   NOR3_X1 i_109 (.A1(n_87), .A2(n_78), .A3(n_93), .ZN(n_77));
   NOR2_X1 i_111 (.A1(multiplicand[20]), .A2(A[20]), .ZN(n_79));
   NOR2_X1 i_116 (.A1(multiplicand[21]), .A2(A[21]), .ZN(n_84));
   OR2_X1 i_119 (.A1(n_89), .A2(n_88), .ZN(n_87));
   OR2_X1 i_121 (.A1(n_92), .A2(n_90), .ZN(n_89));
   NOR2_X1 i_124 (.A1(multiplicand[27]), .A2(A[27]), .ZN(n_92));
   NOR2_X1 i_126 (.A1(n_106), .A2(n_96), .ZN(n_94));
   INV_X1 i_127 (.A(n_96), .ZN(n_95));
   NAND2_X1 i_128 (.A1(multiplicand[18]), .A2(A[18]), .ZN(n_96));
   AND2_X1 i_129 (.A1(multiplicand[19]), .A2(A[19]), .ZN(n_97));
   AOI21_X1 i_130 (.A(n_103), .B1(n_100), .B2(n_99), .ZN(n_98));
   NAND2_X1 i_131 (.A1(multiplicand[17]), .A2(A[17]), .ZN(n_99));
   NAND2_X1 i_132 (.A1(multiplicand[16]), .A2(A[16]), .ZN(n_100));
   NOR3_X1 i_133 (.A1(n_103), .A2(n_102), .A3(n_107), .ZN(n_101));
   NOR2_X1 i_134 (.A1(multiplicand[16]), .A2(A[16]), .ZN(n_102));
   OR3_X1 i_135 (.A1(n_106), .A2(n_104), .A3(n_105), .ZN(n_103));
   NOR2_X1 i_136 (.A1(multiplicand[18]), .A2(A[18]), .ZN(n_104));
   NOR2_X1 i_137 (.A1(multiplicand[17]), .A2(A[17]), .ZN(n_105));
   NOR2_X1 i_138 (.A1(multiplicand[19]), .A2(A[19]), .ZN(n_106));
   NOR4_X1 i_139 (.A1(n_111), .A2(n_108), .A3(n_112), .A4(n_115), .ZN(n_107));
   NOR2_X1 i_140 (.A1(n_120), .A2(n_110), .ZN(n_108));
   INV_X1 i_141 (.A(n_110), .ZN(n_109));
   NAND2_X1 i_142 (.A1(multiplicand[14]), .A2(A[14]), .ZN(n_110));
   AND2_X1 i_143 (.A1(multiplicand[15]), .A2(A[15]), .ZN(n_111));
   AOI21_X1 i_144 (.A(n_117), .B1(n_114), .B2(n_113), .ZN(n_112));
   NAND2_X1 i_145 (.A1(multiplicand[13]), .A2(A[13]), .ZN(n_113));
   NAND2_X1 i_146 (.A1(multiplicand[12]), .A2(A[12]), .ZN(n_114));
   NOR3_X1 i_147 (.A1(n_117), .A2(n_116), .A3(n_121), .ZN(n_115));
   NOR2_X1 i_148 (.A1(multiplicand[12]), .A2(A[12]), .ZN(n_116));
   OR3_X1 i_149 (.A1(n_120), .A2(n_118), .A3(n_119), .ZN(n_117));
   NOR2_X1 i_150 (.A1(multiplicand[14]), .A2(A[14]), .ZN(n_118));
   NOR2_X1 i_151 (.A1(multiplicand[13]), .A2(A[13]), .ZN(n_119));
   NOR2_X1 i_152 (.A1(multiplicand[15]), .A2(A[15]), .ZN(n_120));
   NOR4_X1 i_153 (.A1(n_125), .A2(n_122), .A3(n_126), .A4(n_129), .ZN(n_121));
   NOR2_X1 i_154 (.A1(n_134), .A2(n_124), .ZN(n_122));
   INV_X1 i_155 (.A(n_124), .ZN(n_123));
   NAND2_X1 i_156 (.A1(multiplicand[10]), .A2(A[10]), .ZN(n_124));
   AND2_X1 i_157 (.A1(multiplicand[11]), .A2(A[11]), .ZN(n_125));
   AOI21_X1 i_158 (.A(n_131), .B1(n_128), .B2(n_127), .ZN(n_126));
   NAND2_X1 i_159 (.A1(multiplicand[9]), .A2(A[9]), .ZN(n_127));
   NAND2_X1 i_160 (.A1(multiplicand[8]), .A2(A[8]), .ZN(n_128));
   NOR3_X1 i_161 (.A1(n_131), .A2(n_130), .A3(n_135), .ZN(n_129));
   NOR2_X1 i_162 (.A1(multiplicand[8]), .A2(A[8]), .ZN(n_130));
   OR3_X1 i_163 (.A1(n_134), .A2(n_132), .A3(n_133), .ZN(n_131));
   NOR2_X1 i_164 (.A1(multiplicand[10]), .A2(A[10]), .ZN(n_132));
   NOR2_X1 i_165 (.A1(multiplicand[9]), .A2(A[9]), .ZN(n_133));
   NOR2_X1 i_166 (.A1(multiplicand[11]), .A2(A[11]), .ZN(n_134));
   NOR4_X1 i_167 (.A1(n_139), .A2(n_136), .A3(n_140), .A4(n_143), .ZN(n_135));
   NOR2_X1 i_168 (.A1(n_148), .A2(n_138), .ZN(n_136));
   INV_X1 i_169 (.A(n_138), .ZN(n_137));
   NAND2_X1 i_170 (.A1(multiplicand[6]), .A2(A[6]), .ZN(n_138));
   AND2_X1 i_171 (.A1(multiplicand[7]), .A2(A[7]), .ZN(n_139));
   AOI21_X1 i_172 (.A(n_145), .B1(n_142), .B2(n_141), .ZN(n_140));
   NAND2_X1 i_173 (.A1(multiplicand[5]), .A2(A[5]), .ZN(n_141));
   NAND2_X1 i_174 (.A1(multiplicand[4]), .A2(A[4]), .ZN(n_142));
   NOR3_X1 i_175 (.A1(n_145), .A2(n_144), .A3(n_149), .ZN(n_143));
   NOR2_X1 i_176 (.A1(multiplicand[4]), .A2(A[4]), .ZN(n_144));
   OR3_X1 i_177 (.A1(n_148), .A2(n_146), .A3(n_147), .ZN(n_145));
   NOR2_X1 i_178 (.A1(multiplicand[6]), .A2(A[6]), .ZN(n_146));
   NOR2_X1 i_179 (.A1(multiplicand[5]), .A2(A[5]), .ZN(n_147));
   NOR2_X1 i_180 (.A1(multiplicand[7]), .A2(A[7]), .ZN(n_148));
   NAND2_X1 i_181 (.A1(n_158), .A2(n_150), .ZN(n_149));
   OAI21_X1 i_182 (.A(n_151), .B1(n_164), .B2(n_161), .ZN(n_150));
   OAI22_X1 i_183 (.A1(multiplicand[2]), .A2(A[2]), .B1(n_156), .B2(n_152), 
      .ZN(n_151));
   AOI21_X1 i_184 (.A(n_155), .B1(n_154), .B2(n_153), .ZN(n_152));
   NAND2_X1 i_185 (.A1(multiplicand[1]), .A2(A[1]), .ZN(n_153));
   NAND2_X1 i_186 (.A1(multiplicand[0]), .A2(A[0]), .ZN(n_154));
   NOR2_X1 i_187 (.A1(multiplicand[1]), .A2(A[1]), .ZN(n_155));
   INV_X1 i_188 (.A(n_157), .ZN(n_156));
   NAND2_X1 i_189 (.A1(multiplicand[2]), .A2(A[2]), .ZN(n_157));
   NAND2_X1 i_190 (.A1(n_164), .A2(n_161), .ZN(n_158));
   NOR2_X1 i_191 (.A1(multiplicand[28]), .A2(A[28]), .ZN(n_159));
   NAND2_X1 i_192 (.A1(n_166), .A2(n_163), .ZN(n_160));
   INV_X1 i_193 (.A(A[3]), .ZN(n_161));
   INV_X1 i_194 (.A(A[27]), .ZN(n_162));
   INV_X1 i_195 (.A(A[31]), .ZN(n_163));
   INV_X1 i_196 (.A(multiplicand[3]), .ZN(n_164));
   INV_X1 i_197 (.A(multiplicand[27]), .ZN(n_165));
   INV_X1 i_198 (.A(multiplicand[30]), .ZN(n_166));
   INV_X1 i_69 (.A(n_179), .ZN(n_88));
   INV_X1 i_70 (.A(n_184), .ZN(n_90));
   INV_X1 i_71 (.A(n_169), .ZN(n_51));
   INV_X1 i_72 (.A(n_171), .ZN(n_72));
   XNOR2_X1 i_73 (.A(n_44), .B(n_45), .ZN(p_0[25]));
   NAND2_X1 i_74 (.A1(n_53), .A2(n_183), .ZN(n_44));
   INV_X1 i_75 (.A(n_168), .ZN(n_45));
   OR2_X1 i_76 (.A1(n_46), .A2(n_48), .ZN(p_0[26]));
   INV_X1 i_77 (.A(n_47), .ZN(n_46));
   NAND3_X1 i_79 (.A1(n_167), .A2(n_53), .A3(n_49), .ZN(n_47));
   AOI21_X1 i_80 (.A(n_49), .B1(n_167), .B2(n_53), .ZN(n_48));
   NAND2_X1 i_81 (.A1(n_52), .A2(n_66), .ZN(n_49));
   INV_X1 i_98 (.A(n_185), .ZN(n_52));
   NAND2_X1 i_101 (.A1(n_187), .A2(n_186), .ZN(n_53));
   NAND2_X1 i_103 (.A1(n_73), .A2(n_85), .ZN(p_0[27]));
   NAND2_X1 i_104 (.A1(n_80), .A2(n_189), .ZN(n_73));
   NAND2_X1 i_105 (.A1(n_91), .A2(n_66), .ZN(n_80));
   NAND3_X1 i_107 (.A1(n_91), .A2(n_188), .A3(n_66), .ZN(n_85));
   NAND2_X1 i_108 (.A1(n_184), .A2(n_167), .ZN(n_91));
   NAND2_X1 i_110 (.A1(n_183), .A2(n_168), .ZN(n_167));
   AOI21_X1 i_112 (.A(n_182), .B1(n_169), .B2(n_179), .ZN(n_168));
   NAND2_X1 i_113 (.A1(n_71), .A2(n_175), .ZN(n_169));
   INV_X1 i_114 (.A(n_170), .ZN(n_71));
   OAI211_X1 i_115 (.A(n_173), .B(n_172), .C1(n_86), .C2(n_171), .ZN(n_170));
   NAND2_X1 i_117 (.A1(multiplicand[22]), .A2(A[22]), .ZN(n_171));
   NAND2_X1 i_118 (.A1(multiplicand[23]), .A2(A[23]), .ZN(n_172));
   OAI211_X1 i_120 (.A(n_176), .B(n_174), .C1(multiplicand[23]), .C2(A[23]), 
      .ZN(n_173));
   NAND2_X1 i_122 (.A1(n_75), .A2(n_76), .ZN(n_174));
   NAND2_X1 i_123 (.A1(multiplicand[21]), .A2(A[21]), .ZN(n_75));
   NAND2_X1 i_125 (.A1(multiplicand[20]), .A2(A[20]), .ZN(n_76));
   NOR2_X1 i_199 (.A1(multiplicand[23]), .A2(A[23]), .ZN(n_86));
   OR2_X1 i_200 (.A1(n_78), .A2(n_93), .ZN(n_175));
   NOR4_X1 i_201 (.A1(n_101), .A2(n_98), .A3(n_97), .A4(n_94), .ZN(n_93));
   OAI211_X1 i_202 (.A(n_178), .B(n_176), .C1(multiplicand[23]), .C2(A[23]), 
      .ZN(n_78));
   INV_X1 i_203 (.A(n_177), .ZN(n_176));
   NAND2_X1 i_204 (.A1(n_81), .A2(n_83), .ZN(n_177));
   INV_X1 i_205 (.A(n_82), .ZN(n_81));
   NOR2_X1 i_206 (.A1(multiplicand[22]), .A2(A[22]), .ZN(n_82));
   INV_X1 i_207 (.A(n_84), .ZN(n_83));
   INV_X1 i_208 (.A(n_79), .ZN(n_178));
   NAND2_X1 i_209 (.A1(n_181), .A2(n_180), .ZN(n_179));
   INV_X1 i_210 (.A(A[24]), .ZN(n_180));
   INV_X1 i_211 (.A(multiplicand[24]), .ZN(n_181));
   INV_X1 i_212 (.A(n_69), .ZN(n_182));
   NAND2_X1 i_213 (.A1(multiplicand[24]), .A2(A[24]), .ZN(n_69));
   NAND2_X1 i_214 (.A1(multiplicand[25]), .A2(A[25]), .ZN(n_183));
   AOI21_X1 i_215 (.A(n_185), .B1(n_187), .B2(n_186), .ZN(n_184));
   NOR2_X1 i_216 (.A1(multiplicand[26]), .A2(A[26]), .ZN(n_185));
   INV_X1 i_217 (.A(A[25]), .ZN(n_186));
   INV_X1 i_218 (.A(multiplicand[25]), .ZN(n_187));
   NAND2_X1 i_219 (.A1(multiplicand[26]), .A2(A[26]), .ZN(n_66));
   INV_X1 i_220 (.A(n_189), .ZN(n_188));
   OAI22_X1 i_221 (.A1(n_165), .A2(n_162), .B1(multiplicand[27]), .B2(A[27]), 
      .ZN(n_189));
endmodule

module datapath__0_67(p_0, b);
   output [31:0]p_0;
   input [31:0]b;

   AOI21_X1 i_0 (.A(n_62), .B1(b[1]), .B2(b[0]), .ZN(p_0[1]));
   AOI21_X1 i_1 (.A(n_60), .B1(b[2]), .B2(n_61), .ZN(p_0[2]));
   AOI21_X1 i_2 (.A(n_58), .B1(b[3]), .B2(n_59), .ZN(p_0[3]));
   AOI21_X1 i_3 (.A(n_5), .B1(b[4]), .B2(n_57), .ZN(p_0[4]));
   AOI21_X1 i_5 (.A(n_1), .B1(b[6]), .B2(n_2), .ZN(p_0[6]));
   NOR2_X1 i_8 (.A1(n_57), .A2(n_56), .ZN(n_1));
   INV_X1 i_9 (.A(n_3), .ZN(n_2));
   AOI21_X1 i_15 (.A(n_7), .B1(b[10]), .B2(n_8), .ZN(p_0[10]));
   NOR2_X1 i_18 (.A1(n_54), .A2(n_53), .ZN(n_7));
   INV_X1 i_19 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_25 (.A(n_13), .B1(b[14]), .B2(n_14), .ZN(p_0[14]));
   NOR2_X1 i_28 (.A1(n_51), .A2(n_50), .ZN(n_13));
   INV_X1 i_29 (.A(n_15), .ZN(n_14));
   AOI21_X1 i_34 (.A(n_21), .B1(b[17]), .B2(n_22), .ZN(p_0[17]));
   AOI21_X1 i_35 (.A(n_19), .B1(b[18]), .B2(n_20), .ZN(p_0[18]));
   AOI21_X1 i_36 (.A(n_45), .B1(b[19]), .B2(n_18), .ZN(p_0[19]));
   INV_X1 i_37 (.A(n_19), .ZN(n_18));
   NOR2_X1 i_38 (.A1(n_48), .A2(n_46), .ZN(n_19));
   INV_X1 i_39 (.A(n_21), .ZN(n_20));
   NOR2_X1 i_40 (.A1(b[17]), .A2(n_22), .ZN(n_21));
   INV_X1 i_41 (.A(n_23), .ZN(n_22));
   AOI21_X1 i_43 (.A(n_25), .B1(b[20]), .B2(n_44), .ZN(p_0[20]));
   AOI21_X1 i_44 (.A(n_27), .B1(b[21]), .B2(n_24), .ZN(p_0[21]));
   INV_X1 i_45 (.A(n_25), .ZN(n_24));
   NOR2_X1 i_46 (.A1(b[20]), .A2(n_44), .ZN(n_25));
   AOI21_X1 i_47 (.A(n_43), .B1(b[22]), .B2(n_26), .ZN(p_0[22]));
   INV_X1 i_48 (.A(n_27), .ZN(n_26));
   NOR3_X1 i_49 (.A1(b[21]), .A2(b[20]), .A3(n_44), .ZN(n_27));
   AOI21_X1 i_50 (.A(n_41), .B1(b[23]), .B2(n_42), .ZN(p_0[23]));
   AOI21_X1 i_51 (.A(n_29), .B1(b[24]), .B2(n_40), .ZN(p_0[24]));
   INV_X1 i_52 (.A(n_28), .ZN(p_0[25]));
   OAI21_X1 i_53 (.A(n_30), .B1(n_63), .B2(n_29), .ZN(n_28));
   NOR2_X1 i_54 (.A1(b[24]), .A2(n_40), .ZN(n_29));
   AOI21_X1 i_55 (.A(n_32), .B1(b[26]), .B2(n_30), .ZN(p_0[26]));
   OR3_X1 i_56 (.A1(b[25]), .A2(b[24]), .A3(n_40), .ZN(n_30));
   AOI21_X1 i_57 (.A(n_39), .B1(b[27]), .B2(n_31), .ZN(p_0[27]));
   INV_X1 i_58 (.A(n_32), .ZN(n_31));
   NOR2_X1 i_59 (.A1(n_47), .A2(n_40), .ZN(n_32));
   AOI21_X1 i_60 (.A(n_34), .B1(b[28]), .B2(n_38), .ZN(p_0[28]));
   AOI21_X1 i_61 (.A(n_36), .B1(b[29]), .B2(n_33), .ZN(p_0[29]));
   INV_X1 i_62 (.A(n_34), .ZN(n_33));
   NOR2_X1 i_63 (.A1(b[28]), .A2(n_38), .ZN(n_34));
   AOI21_X1 i_64 (.A(n_37), .B1(b[30]), .B2(n_35), .ZN(p_0[30]));
   INV_X1 i_65 (.A(n_36), .ZN(n_35));
   NOR3_X1 i_66 (.A1(b[29]), .A2(b[28]), .A3(n_38), .ZN(n_36));
   XNOR2_X1 i_67 (.A(b[31]), .B(n_37), .ZN(p_0[31]));
   NOR4_X1 i_68 (.A1(b[29]), .A2(b[28]), .A3(b[30]), .A4(n_38), .ZN(n_37));
   INV_X1 i_69 (.A(n_39), .ZN(n_38));
   NOR3_X1 i_70 (.A1(b[27]), .A2(n_47), .A3(n_40), .ZN(n_39));
   INV_X1 i_71 (.A(n_41), .ZN(n_40));
   NOR2_X1 i_72 (.A1(b[23]), .A2(n_42), .ZN(n_41));
   INV_X1 i_73 (.A(n_43), .ZN(n_42));
   NOR4_X1 i_74 (.A1(b[22]), .A2(b[21]), .A3(b[20]), .A4(n_44), .ZN(n_43));
   INV_X1 i_75 (.A(n_45), .ZN(n_44));
   NOR3_X1 i_76 (.A1(b[19]), .A2(n_46), .A3(n_48), .ZN(n_45));
   OR3_X1 i_77 (.A1(b[18]), .A2(b[16]), .A3(b[17]), .ZN(n_46));
   OR3_X1 i_78 (.A1(b[26]), .A2(b[25]), .A3(b[24]), .ZN(n_47));
   INV_X1 i_94 (.A(b[25]), .ZN(n_63));
   INV_X1 i_4 (.A(n_0), .ZN(n_23));
   OR2_X1 i_6 (.A1(n_48), .A2(b[16]), .ZN(n_0));
   INV_X1 i_7 (.A(n_68), .ZN(n_15));
   INV_X1 i_10 (.A(n_49), .ZN(n_9));
   INV_X1 i_11 (.A(n_4), .ZN(n_3));
   NAND2_X1 i_12 (.A1(n_5), .A2(n_11), .ZN(n_4));
   INV_X1 i_13 (.A(n_6), .ZN(n_5));
   XNOR2_X1 i_14 (.A(n_6), .B(n_11), .ZN(p_0[5]));
   NAND2_X1 i_16 (.A1(n_58), .A2(n_10), .ZN(n_6));
   INV_X1 i_17 (.A(b[4]), .ZN(n_10));
   INV_X1 i_20 (.A(b[5]), .ZN(n_11));
   AOI21_X1 i_21 (.A(n_79), .B1(n_12), .B2(b[7]), .ZN(p_0[7]));
   INV_X1 i_22 (.A(n_1), .ZN(n_12));
   XNOR2_X1 i_23 (.A(n_54), .B(n_52), .ZN(p_0[8]));
   INV_X1 i_24 (.A(n_16), .ZN(p_0[9]));
   NAND2_X1 i_26 (.A1(n_17), .A2(n_49), .ZN(n_16));
   OAI21_X1 i_27 (.A(b[9]), .B1(n_54), .B2(b[8]), .ZN(n_17));
   NAND3_X1 i_30 (.A1(n_79), .A2(n_55), .A3(n_52), .ZN(n_49));
   INV_X1 i_31 (.A(b[8]), .ZN(n_52));
   INV_X1 i_32 (.A(b[9]), .ZN(n_55));
   AOI21_X1 i_33 (.A(n_76), .B1(n_64), .B2(b[11]), .ZN(p_0[11]));
   INV_X1 i_42 (.A(n_7), .ZN(n_64));
   INV_X1 i_79 (.A(n_65), .ZN(p_0[12]));
   XNOR2_X1 i_80 (.A(n_51), .B(b[12]), .ZN(n_65));
   INV_X1 i_81 (.A(n_66), .ZN(p_0[13]));
   NAND2_X1 i_82 (.A1(n_67), .A2(n_68), .ZN(n_66));
   OAI21_X1 i_83 (.A(b[13]), .B1(n_51), .B2(b[12]), .ZN(n_67));
   NAND3_X1 i_84 (.A1(n_76), .A2(n_70), .A3(n_69), .ZN(n_68));
   INV_X1 i_85 (.A(b[12]), .ZN(n_69));
   INV_X1 i_86 (.A(b[13]), .ZN(n_70));
   AOI21_X1 i_87 (.A(n_71), .B1(n_72), .B2(b[15]), .ZN(p_0[15]));
   INV_X1 i_88 (.A(n_48), .ZN(n_71));
   INV_X1 i_89 (.A(n_13), .ZN(n_72));
   INV_X1 i_90 (.A(n_73), .ZN(p_0[16]));
   XNOR2_X1 i_91 (.A(n_48), .B(b[16]), .ZN(n_73));
   NAND2_X1 i_92 (.A1(n_76), .A2(n_74), .ZN(n_48));
   INV_X1 i_93 (.A(n_75), .ZN(n_74));
   OR2_X1 i_95 (.A1(n_50), .A2(b[15]), .ZN(n_75));
   OR3_X1 i_96 (.A1(b[14]), .A2(b[13]), .A3(b[12]), .ZN(n_50));
   INV_X1 i_97 (.A(n_51), .ZN(n_76));
   NAND2_X1 i_98 (.A1(n_79), .A2(n_77), .ZN(n_51));
   INV_X1 i_99 (.A(n_78), .ZN(n_77));
   OR2_X1 i_100 (.A1(n_53), .A2(b[11]), .ZN(n_78));
   OR3_X1 i_101 (.A1(b[10]), .A2(b[9]), .A3(b[8]), .ZN(n_53));
   INV_X1 i_102 (.A(n_54), .ZN(n_79));
   NAND2_X1 i_103 (.A1(n_80), .A2(n_58), .ZN(n_54));
   INV_X1 i_104 (.A(n_81), .ZN(n_80));
   OR2_X1 i_105 (.A1(n_56), .A2(b[7]), .ZN(n_81));
   OR3_X1 i_106 (.A1(b[6]), .A2(b[5]), .A3(b[4]), .ZN(n_56));
   INV_X1 i_107 (.A(n_57), .ZN(n_58));
   NAND2_X1 i_108 (.A1(n_60), .A2(n_85), .ZN(n_57));
   INV_X1 i_109 (.A(n_59), .ZN(n_60));
   NAND2_X1 i_110 (.A1(n_62), .A2(n_84), .ZN(n_59));
   INV_X1 i_111 (.A(n_61), .ZN(n_62));
   NAND2_X1 i_112 (.A1(n_83), .A2(n_82), .ZN(n_61));
   INV_X1 i_113 (.A(b[0]), .ZN(n_82));
   INV_X1 i_114 (.A(b[1]), .ZN(n_83));
   INV_X1 i_115 (.A(b[2]), .ZN(n_84));
   INV_X1 i_116 (.A(b[3]), .ZN(n_85));
endmodule

module datapath__0_72(p_0, p_1);
   output [63:0]p_0;
   input [63:0]p_1;

   AOI21_X1 i_0 (.A(n_127), .B1(p_1[1]), .B2(p_1[0]), .ZN(p_0[1]));
   AOI21_X1 i_1 (.A(n_125), .B1(p_1[2]), .B2(n_126), .ZN(p_0[2]));
   AOI21_X1 i_2 (.A(n_123), .B1(p_1[3]), .B2(n_124), .ZN(p_0[3]));
   AOI21_X1 i_3 (.A(n_5), .B1(p_1[4]), .B2(n_122), .ZN(p_0[4]));
   AOI21_X1 i_4 (.A(n_3), .B1(p_1[5]), .B2(n_4), .ZN(p_0[5]));
   AOI21_X1 i_5 (.A(n_1), .B1(p_1[6]), .B2(n_2), .ZN(p_0[6]));
   AOI21_X1 i_6 (.A(n_120), .B1(p_1[7]), .B2(n_0), .ZN(p_0[7]));
   INV_X1 i_7 (.A(n_1), .ZN(n_0));
   NOR2_X1 i_8 (.A1(n_122), .A2(n_121), .ZN(n_1));
   INV_X1 i_9 (.A(n_3), .ZN(n_2));
   NOR2_X1 i_10 (.A1(p_1[5]), .A2(n_4), .ZN(n_3));
   INV_X1 i_11 (.A(n_5), .ZN(n_4));
   NOR2_X1 i_12 (.A1(p_1[4]), .A2(n_122), .ZN(n_5));
   AOI21_X1 i_13 (.A(n_11), .B1(p_1[8]), .B2(n_119), .ZN(p_0[8]));
   AOI21_X1 i_14 (.A(n_9), .B1(p_1[9]), .B2(n_10), .ZN(p_0[9]));
   AOI21_X1 i_15 (.A(n_7), .B1(p_1[10]), .B2(n_8), .ZN(p_0[10]));
   AOI21_X1 i_16 (.A(n_117), .B1(p_1[11]), .B2(n_6), .ZN(p_0[11]));
   INV_X1 i_17 (.A(n_7), .ZN(n_6));
   NOR2_X1 i_18 (.A1(n_119), .A2(n_118), .ZN(n_7));
   INV_X1 i_19 (.A(n_9), .ZN(n_8));
   NOR2_X1 i_20 (.A1(p_1[9]), .A2(n_10), .ZN(n_9));
   INV_X1 i_21 (.A(n_11), .ZN(n_10));
   NOR2_X1 i_22 (.A1(p_1[8]), .A2(n_119), .ZN(n_11));
   AOI21_X1 i_23 (.A(n_17), .B1(p_1[12]), .B2(n_116), .ZN(p_0[12]));
   AOI21_X1 i_24 (.A(n_15), .B1(p_1[13]), .B2(n_16), .ZN(p_0[13]));
   AOI21_X1 i_25 (.A(n_13), .B1(p_1[14]), .B2(n_14), .ZN(p_0[14]));
   AOI21_X1 i_26 (.A(n_114), .B1(p_1[15]), .B2(n_12), .ZN(p_0[15]));
   INV_X1 i_27 (.A(n_13), .ZN(n_12));
   NOR2_X1 i_28 (.A1(n_116), .A2(n_115), .ZN(n_13));
   INV_X1 i_29 (.A(n_15), .ZN(n_14));
   NOR2_X1 i_30 (.A1(p_1[13]), .A2(n_16), .ZN(n_15));
   INV_X1 i_31 (.A(n_17), .ZN(n_16));
   NOR2_X1 i_32 (.A1(p_1[12]), .A2(n_116), .ZN(n_17));
   AOI21_X1 i_33 (.A(n_112), .B1(p_1[16]), .B2(n_113), .ZN(p_0[16]));
   AOI21_X1 i_34 (.A(n_110), .B1(p_1[17]), .B2(n_111), .ZN(p_0[17]));
   AOI21_X1 i_35 (.A(n_108), .B1(p_1[18]), .B2(n_109), .ZN(p_0[18]));
   AOI21_X1 i_36 (.A(n_106), .B1(p_1[19]), .B2(n_107), .ZN(p_0[19]));
   AOI21_X1 i_37 (.A(n_104), .B1(p_1[20]), .B2(n_105), .ZN(p_0[20]));
   AOI21_X1 i_38 (.A(n_102), .B1(p_1[21]), .B2(n_103), .ZN(p_0[21]));
   AOI21_X1 i_39 (.A(n_100), .B1(p_1[22]), .B2(n_101), .ZN(p_0[22]));
   AOI21_X1 i_40 (.A(n_98), .B1(p_1[23]), .B2(n_99), .ZN(p_0[23]));
   AOI21_X1 i_41 (.A(n_96), .B1(p_1[24]), .B2(n_97), .ZN(p_0[24]));
   AOI21_X1 i_42 (.A(n_94), .B1(p_1[25]), .B2(n_95), .ZN(p_0[25]));
   AOI21_X1 i_43 (.A(n_92), .B1(p_1[26]), .B2(n_93), .ZN(p_0[26]));
   AOI21_X1 i_44 (.A(n_90), .B1(p_1[27]), .B2(n_91), .ZN(p_0[27]));
   AOI21_X1 i_45 (.A(n_88), .B1(p_1[28]), .B2(n_89), .ZN(p_0[28]));
   AOI21_X1 i_46 (.A(n_86), .B1(p_1[29]), .B2(n_87), .ZN(p_0[29]));
   AOI21_X1 i_47 (.A(n_84), .B1(p_1[30]), .B2(n_85), .ZN(p_0[30]));
   AOI21_X1 i_48 (.A(n_82), .B1(p_1[31]), .B2(n_83), .ZN(p_0[31]));
   AOI21_X1 i_49 (.A(n_23), .B1(p_1[32]), .B2(n_81), .ZN(p_0[32]));
   AOI21_X1 i_50 (.A(n_21), .B1(p_1[33]), .B2(n_22), .ZN(p_0[33]));
   AOI21_X1 i_51 (.A(n_19), .B1(p_1[34]), .B2(n_20), .ZN(p_0[34]));
   AOI21_X1 i_52 (.A(n_31), .B1(p_1[35]), .B2(n_18), .ZN(p_0[35]));
   INV_X1 i_53 (.A(n_19), .ZN(n_18));
   NOR2_X1 i_54 (.A1(p_1[34]), .A2(n_20), .ZN(n_19));
   INV_X1 i_55 (.A(n_21), .ZN(n_20));
   NOR2_X1 i_56 (.A1(p_1[33]), .A2(n_22), .ZN(n_21));
   INV_X1 i_57 (.A(n_23), .ZN(n_22));
   NOR2_X1 i_58 (.A1(p_1[32]), .A2(n_81), .ZN(n_23));
   AOI21_X1 i_59 (.A(n_29), .B1(p_1[36]), .B2(n_30), .ZN(p_0[36]));
   AOI21_X1 i_60 (.A(n_27), .B1(p_1[37]), .B2(n_28), .ZN(p_0[37]));
   AOI21_X1 i_61 (.A(n_25), .B1(p_1[38]), .B2(n_26), .ZN(p_0[38]));
   AOI21_X1 i_62 (.A(n_77), .B1(p_1[39]), .B2(n_24), .ZN(p_0[39]));
   INV_X1 i_63 (.A(n_25), .ZN(n_24));
   NOR2_X1 i_64 (.A1(p_1[38]), .A2(n_26), .ZN(n_25));
   INV_X1 i_65 (.A(n_27), .ZN(n_26));
   NOR2_X1 i_66 (.A1(p_1[37]), .A2(n_28), .ZN(n_27));
   INV_X1 i_67 (.A(n_29), .ZN(n_28));
   NOR2_X1 i_68 (.A1(p_1[36]), .A2(n_30), .ZN(n_29));
   INV_X1 i_69 (.A(n_31), .ZN(n_30));
   NOR2_X1 i_70 (.A1(n_81), .A2(n_79), .ZN(n_31));
   AOI21_X1 i_71 (.A(n_37), .B1(p_1[40]), .B2(n_76), .ZN(p_0[40]));
   AOI21_X1 i_72 (.A(n_35), .B1(p_1[41]), .B2(n_36), .ZN(p_0[41]));
   AOI21_X1 i_73 (.A(n_33), .B1(p_1[42]), .B2(n_34), .ZN(p_0[42]));
   AOI21_X1 i_74 (.A(n_75), .B1(p_1[43]), .B2(n_32), .ZN(p_0[43]));
   INV_X1 i_75 (.A(n_33), .ZN(n_32));
   NOR2_X1 i_76 (.A1(n_80), .A2(n_76), .ZN(n_33));
   INV_X1 i_77 (.A(n_35), .ZN(n_34));
   NOR2_X1 i_78 (.A1(p_1[41]), .A2(n_36), .ZN(n_35));
   INV_X1 i_79 (.A(n_37), .ZN(n_36));
   NOR2_X1 i_80 (.A1(p_1[40]), .A2(n_76), .ZN(n_37));
   AOI21_X1 i_81 (.A(n_73), .B1(p_1[44]), .B2(n_74), .ZN(p_0[44]));
   AOI21_X1 i_82 (.A(n_71), .B1(p_1[45]), .B2(n_72), .ZN(p_0[45]));
   AOI21_X1 i_83 (.A(n_69), .B1(p_1[46]), .B2(n_70), .ZN(p_0[46]));
   AOI21_X1 i_84 (.A(n_67), .B1(p_1[47]), .B2(n_68), .ZN(p_0[47]));
   AOI21_X1 i_85 (.A(n_43), .B1(p_1[48]), .B2(n_66), .ZN(p_0[48]));
   AOI21_X1 i_86 (.A(n_41), .B1(p_1[49]), .B2(n_42), .ZN(p_0[49]));
   AOI21_X1 i_87 (.A(n_39), .B1(p_1[50]), .B2(n_40), .ZN(p_0[50]));
   INV_X1 i_88 (.A(n_38), .ZN(p_0[51]));
   OAI21_X1 i_89 (.A(n_49), .B1(n_128), .B2(n_39), .ZN(n_38));
   NOR2_X1 i_90 (.A1(p_1[50]), .A2(n_40), .ZN(n_39));
   INV_X1 i_91 (.A(n_41), .ZN(n_40));
   NOR2_X1 i_92 (.A1(p_1[49]), .A2(n_42), .ZN(n_41));
   INV_X1 i_93 (.A(n_43), .ZN(n_42));
   NOR2_X1 i_94 (.A1(p_1[48]), .A2(n_66), .ZN(n_43));
   AOI21_X1 i_95 (.A(n_45), .B1(p_1[52]), .B2(n_49), .ZN(p_0[52]));
   INV_X1 i_96 (.A(n_44), .ZN(p_0[53]));
   OAI21_X1 i_97 (.A(n_46), .B1(n_129), .B2(n_45), .ZN(n_44));
   NOR2_X1 i_98 (.A1(p_1[52]), .A2(n_49), .ZN(n_45));
   AOI21_X1 i_99 (.A(n_48), .B1(p_1[54]), .B2(n_46), .ZN(p_0[54]));
   OR3_X1 i_100 (.A1(p_1[53]), .A2(p_1[52]), .A3(n_49), .ZN(n_46));
   AOI21_X1 i_101 (.A(n_62), .B1(p_1[55]), .B2(n_47), .ZN(p_0[55]));
   INV_X1 i_102 (.A(n_48), .ZN(n_47));
   NOR2_X1 i_103 (.A1(n_63), .A2(n_49), .ZN(n_48));
   OR2_X1 i_104 (.A1(n_66), .A2(n_64), .ZN(n_49));
   AOI21_X1 i_105 (.A(n_51), .B1(p_1[56]), .B2(n_61), .ZN(p_0[56]));
   INV_X1 i_106 (.A(n_50), .ZN(p_0[57]));
   OAI21_X1 i_107 (.A(n_52), .B1(n_130), .B2(n_51), .ZN(n_50));
   NOR2_X1 i_108 (.A1(p_1[56]), .A2(n_61), .ZN(n_51));
   AOI21_X1 i_109 (.A(n_54), .B1(p_1[58]), .B2(n_52), .ZN(p_0[58]));
   OR3_X1 i_110 (.A1(p_1[57]), .A2(p_1[56]), .A3(n_61), .ZN(n_52));
   AOI21_X1 i_111 (.A(n_60), .B1(p_1[59]), .B2(n_53), .ZN(p_0[59]));
   INV_X1 i_112 (.A(n_54), .ZN(n_53));
   NOR2_X1 i_113 (.A1(n_65), .A2(n_61), .ZN(n_54));
   INV_X1 i_191 (.A(p_1[51]), .ZN(n_128));
   INV_X1 i_192 (.A(p_1[53]), .ZN(n_129));
   INV_X1 i_193 (.A(p_1[57]), .ZN(n_130));
   NAND3_X1 i_114 (.A1(n_134), .A2(n_133), .A3(n_132), .ZN(n_65));
   INV_X1 i_115 (.A(n_66), .ZN(n_67));
   INV_X1 i_116 (.A(n_88), .ZN(n_87));
   INV_X1 i_117 (.A(n_91), .ZN(n_92));
   INV_X1 i_118 (.A(n_96), .ZN(n_95));
   INV_X1 i_119 (.A(n_107), .ZN(n_108));
   INV_X1 i_120 (.A(n_112), .ZN(n_111));
   NAND2_X1 i_121 (.A1(n_78), .A2(n_155), .ZN(n_115));
   INV_X1 i_122 (.A(n_113), .ZN(n_114));
   INV_X1 i_123 (.A(n_117), .ZN(n_116));
   NAND2_X1 i_124 (.A1(n_169), .A2(n_58), .ZN(n_121));
   INV_X1 i_125 (.A(n_119), .ZN(n_120));
   OR2_X1 i_126 (.A1(n_80), .A2(p_1[43]), .ZN(n_55));
   OR3_X1 i_127 (.A1(p_1[42]), .A2(p_1[41]), .A3(p_1[40]), .ZN(n_80));
   OR4_X1 i_128 (.A1(p_1[39]), .A2(n_57), .A3(p_1[38]), .A4(p_1[37]), .ZN(n_56));
   OR2_X1 i_129 (.A1(n_79), .A2(p_1[36]), .ZN(n_57));
   OR4_X1 i_130 (.A1(p_1[35]), .A2(p_1[34]), .A3(p_1[33]), .A4(p_1[32]), 
      .ZN(n_79));
   INV_X1 i_131 (.A(n_59), .ZN(n_58));
   NAND2_X1 i_132 (.A1(n_168), .A2(n_167), .ZN(n_59));
   INV_X1 i_133 (.A(n_131), .ZN(n_78));
   NAND2_X1 i_134 (.A1(n_157), .A2(n_156), .ZN(n_131));
   INV_X1 i_135 (.A(p_1[56]), .ZN(n_132));
   INV_X1 i_136 (.A(p_1[57]), .ZN(n_133));
   INV_X1 i_137 (.A(p_1[58]), .ZN(n_134));
   NAND2_X1 i_138 (.A1(n_69), .A2(n_196), .ZN(n_66));
   INV_X1 i_139 (.A(n_72), .ZN(n_73));
   NAND2_X1 i_140 (.A1(n_75), .A2(n_193), .ZN(n_72));
   INV_X1 i_141 (.A(n_81), .ZN(n_82));
   NAND2_X1 i_142 (.A1(n_84), .A2(n_192), .ZN(n_81));
   INV_X1 i_143 (.A(n_135), .ZN(n_88));
   NAND2_X1 i_144 (.A1(n_90), .A2(n_187), .ZN(n_135));
   INV_X1 i_145 (.A(n_93), .ZN(n_94));
   NAND2_X1 i_146 (.A1(n_96), .A2(n_184), .ZN(n_93));
   INV_X1 i_147 (.A(n_99), .ZN(n_100));
   NAND2_X1 i_148 (.A1(n_102), .A2(n_181), .ZN(n_99));
   INV_X1 i_149 (.A(n_105), .ZN(n_106));
   NAND2_X1 i_150 (.A1(n_151), .A2(n_178), .ZN(n_105));
   INV_X1 i_151 (.A(n_136), .ZN(n_112));
   NAND2_X1 i_152 (.A1(n_152), .A2(n_175), .ZN(n_136));
   NAND3_X1 i_153 (.A1(n_163), .A2(n_162), .A3(n_161), .ZN(n_118));
   NAND2_X1 i_154 (.A1(n_123), .A2(n_165), .ZN(n_119));
   INV_X1 i_155 (.A(n_124), .ZN(n_125));
   NAND2_X1 i_156 (.A1(n_127), .A2(n_173), .ZN(n_124));
   INV_X1 i_157 (.A(n_126), .ZN(n_127));
   NAND2_X1 i_158 (.A1(n_172), .A2(n_171), .ZN(n_126));
   INV_X1 i_159 (.A(n_137), .ZN(p_0[60]));
   XNOR2_X1 i_160 (.A(n_145), .B(p_1[60]), .ZN(n_137));
   NOR2_X1 i_161 (.A1(n_138), .A2(n_139), .ZN(p_0[61]));
   AOI21_X1 i_162 (.A(n_198), .B1(n_60), .B2(n_197), .ZN(n_138));
   INV_X1 i_163 (.A(n_142), .ZN(n_139));
   INV_X1 i_164 (.A(n_140), .ZN(p_0[62]));
   NAND2_X1 i_165 (.A1(n_141), .A2(p_0[63]), .ZN(n_140));
   NAND2_X1 i_166 (.A1(n_142), .A2(p_1[62]), .ZN(n_141));
   NAND4_X1 i_167 (.A1(n_62), .A2(n_198), .A3(n_197), .A4(n_146), .ZN(n_142));
   INV_X1 i_168 (.A(n_61), .ZN(n_62));
   NAND4_X1 i_169 (.A1(n_71), .A2(n_196), .A3(n_195), .A4(n_148), .ZN(n_61));
   INV_X1 i_170 (.A(n_70), .ZN(n_71));
   NAND4_X1 i_171 (.A1(n_77), .A2(n_194), .A3(n_193), .A4(n_191), .ZN(n_70));
   INV_X1 i_172 (.A(n_76), .ZN(n_77));
   NAND4_X1 i_173 (.A1(n_86), .A2(n_192), .A3(n_189), .A4(n_190), .ZN(n_76));
   INV_X1 i_174 (.A(n_85), .ZN(n_86));
   NAND4_X1 i_175 (.A1(n_143), .A2(n_188), .A3(n_187), .A4(n_186), .ZN(n_85));
   INV_X1 i_176 (.A(n_91), .ZN(n_143));
   NAND4_X1 i_177 (.A1(n_98), .A2(n_185), .A3(n_184), .A4(n_183), .ZN(n_91));
   INV_X1 i_178 (.A(n_97), .ZN(n_98));
   NAND4_X1 i_179 (.A1(n_104), .A2(n_182), .A3(n_181), .A4(n_180), .ZN(n_97));
   INV_X1 i_180 (.A(n_103), .ZN(n_104));
   NAND4_X1 i_181 (.A1(n_110), .A2(n_179), .A3(n_178), .A4(n_177), .ZN(n_103));
   INV_X1 i_182 (.A(n_109), .ZN(n_110));
   NAND4_X1 i_183 (.A1(n_117), .A2(n_176), .A3(n_175), .A4(n_153), .ZN(n_109));
   INV_X1 i_184 (.A(n_144), .ZN(n_117));
   NAND3_X1 i_185 (.A1(n_123), .A2(n_165), .A3(n_159), .ZN(n_144));
   NAND4_X1 i_186 (.A1(n_60), .A2(n_199), .A3(n_198), .A4(n_197), .ZN(p_0[63]));
   INV_X1 i_187 (.A(n_145), .ZN(n_60));
   NAND4_X1 i_188 (.A1(n_69), .A2(n_196), .A3(n_148), .A4(n_146), .ZN(n_145));
   INV_X1 i_189 (.A(n_147), .ZN(n_146));
   OR4_X1 i_190 (.A1(p_1[59]), .A2(p_1[58]), .A3(p_1[57]), .A4(p_1[56]), 
      .ZN(n_147));
   INV_X1 i_194 (.A(n_149), .ZN(n_148));
   OR3_X1 i_195 (.A1(n_64), .A2(n_63), .A3(p_1[55]), .ZN(n_149));
   OR3_X1 i_196 (.A1(p_1[54]), .A2(p_1[53]), .A3(p_1[52]), .ZN(n_63));
   OR4_X1 i_197 (.A1(p_1[51]), .A2(p_1[50]), .A3(p_1[49]), .A4(p_1[48]), 
      .ZN(n_64));
   INV_X1 i_198 (.A(n_68), .ZN(n_69));
   NAND4_X1 i_199 (.A1(n_75), .A2(n_195), .A3(n_194), .A4(n_193), .ZN(n_68));
   INV_X1 i_200 (.A(n_74), .ZN(n_75));
   NAND4_X1 i_201 (.A1(n_84), .A2(n_192), .A3(n_191), .A4(n_190), .ZN(n_74));
   INV_X1 i_202 (.A(n_83), .ZN(n_84));
   NAND4_X1 i_203 (.A1(n_90), .A2(n_189), .A3(n_188), .A4(n_187), .ZN(n_83));
   INV_X1 i_204 (.A(n_89), .ZN(n_90));
   NAND4_X1 i_205 (.A1(n_96), .A2(n_186), .A3(n_185), .A4(n_184), .ZN(n_89));
   INV_X1 i_206 (.A(n_150), .ZN(n_96));
   NAND4_X1 i_207 (.A1(n_102), .A2(n_183), .A3(n_182), .A4(n_181), .ZN(n_150));
   INV_X1 i_208 (.A(n_101), .ZN(n_102));
   NAND4_X1 i_209 (.A1(n_151), .A2(n_180), .A3(n_179), .A4(n_178), .ZN(n_101));
   INV_X1 i_210 (.A(n_107), .ZN(n_151));
   NAND4_X1 i_211 (.A1(n_152), .A2(n_177), .A3(n_176), .A4(n_175), .ZN(n_107));
   INV_X1 i_212 (.A(n_113), .ZN(n_152));
   NAND4_X1 i_213 (.A1(n_123), .A2(n_165), .A3(n_159), .A4(n_153), .ZN(n_113));
   INV_X1 i_214 (.A(n_154), .ZN(n_153));
   NAND4_X1 i_215 (.A1(n_158), .A2(n_157), .A3(n_156), .A4(n_155), .ZN(n_154));
   INV_X1 i_216 (.A(p_1[12]), .ZN(n_155));
   INV_X1 i_217 (.A(p_1[13]), .ZN(n_156));
   INV_X1 i_218 (.A(p_1[14]), .ZN(n_157));
   INV_X1 i_219 (.A(p_1[15]), .ZN(n_158));
   INV_X1 i_220 (.A(n_160), .ZN(n_159));
   NAND4_X1 i_221 (.A1(n_164), .A2(n_163), .A3(n_162), .A4(n_161), .ZN(n_160));
   INV_X1 i_222 (.A(p_1[8]), .ZN(n_161));
   INV_X1 i_223 (.A(p_1[9]), .ZN(n_162));
   INV_X1 i_224 (.A(p_1[10]), .ZN(n_163));
   INV_X1 i_225 (.A(p_1[11]), .ZN(n_164));
   INV_X1 i_226 (.A(n_166), .ZN(n_165));
   NAND4_X1 i_227 (.A1(n_170), .A2(n_169), .A3(n_168), .A4(n_167), .ZN(n_166));
   INV_X1 i_228 (.A(p_1[4]), .ZN(n_167));
   INV_X1 i_229 (.A(p_1[5]), .ZN(n_168));
   INV_X1 i_230 (.A(p_1[6]), .ZN(n_169));
   INV_X1 i_231 (.A(p_1[7]), .ZN(n_170));
   INV_X1 i_232 (.A(n_122), .ZN(n_123));
   NAND4_X1 i_233 (.A1(n_174), .A2(n_173), .A3(n_172), .A4(n_171), .ZN(n_122));
   INV_X1 i_234 (.A(p_1[0]), .ZN(n_171));
   INV_X1 i_235 (.A(p_1[1]), .ZN(n_172));
   INV_X1 i_236 (.A(p_1[2]), .ZN(n_173));
   INV_X1 i_237 (.A(p_1[3]), .ZN(n_174));
   INV_X1 i_238 (.A(p_1[16]), .ZN(n_175));
   INV_X1 i_239 (.A(p_1[17]), .ZN(n_176));
   INV_X1 i_240 (.A(p_1[18]), .ZN(n_177));
   INV_X1 i_241 (.A(p_1[19]), .ZN(n_178));
   INV_X1 i_242 (.A(p_1[20]), .ZN(n_179));
   INV_X1 i_243 (.A(p_1[21]), .ZN(n_180));
   INV_X1 i_244 (.A(p_1[22]), .ZN(n_181));
   INV_X1 i_245 (.A(p_1[23]), .ZN(n_182));
   INV_X1 i_246 (.A(p_1[24]), .ZN(n_183));
   INV_X1 i_247 (.A(p_1[25]), .ZN(n_184));
   INV_X1 i_248 (.A(p_1[26]), .ZN(n_185));
   INV_X1 i_249 (.A(p_1[27]), .ZN(n_186));
   INV_X1 i_250 (.A(p_1[28]), .ZN(n_187));
   INV_X1 i_251 (.A(p_1[29]), .ZN(n_188));
   INV_X1 i_252 (.A(p_1[30]), .ZN(n_189));
   INV_X1 i_253 (.A(n_56), .ZN(n_190));
   INV_X1 i_254 (.A(n_55), .ZN(n_191));
   INV_X1 i_255 (.A(p_1[31]), .ZN(n_192));
   INV_X1 i_256 (.A(p_1[44]), .ZN(n_193));
   INV_X1 i_257 (.A(p_1[45]), .ZN(n_194));
   INV_X1 i_258 (.A(p_1[46]), .ZN(n_195));
   INV_X1 i_259 (.A(p_1[47]), .ZN(n_196));
   INV_X1 i_260 (.A(p_1[60]), .ZN(n_197));
   INV_X1 i_261 (.A(p_1[61]), .ZN(n_198));
   INV_X1 i_262 (.A(p_1[62]), .ZN(n_199));
endmodule

module booth_multiplier(clk, rst, en, a, b, c);
   input clk;
   input rst;
   input en;
   input [31:0]a;
   input [31:0]b;
   output [63:0]c;

   wire n_64_0;
   wire n_64_3;
   wire n_64_4;
   wire n_64_5;
   wire n_64_6;
   wire n_64_7;
   wire n_64_8;
   wire n_64_9;
   wire n_64_10;
   wire n_64_11;
   wire n_64_12;
   wire n_64_13;
   wire n_64_14;
   wire n_64_15;
   wire n_64_16;
   wire n_64_17;
   wire n_64_18;
   wire n_64_19;
   wire n_64_20;
   wire n_64_21;
   wire n_64_22;
   wire n_64_23;
   wire n_64_24;
   wire n_64_25;
   wire n_64_26;
   wire n_64_27;
   wire n_64_28;
   wire n_64_29;
   wire n_64_30;
   wire n_64_31;
   wire n_64_32;
   wire n_64_33;
   wire n_64_34;
   wire n_64_35;
   wire n_64_36;
   wire n_64_37;
   wire n_64_38;
   wire n_64_39;
   wire n_64_40;
   wire n_64_41;
   wire n_64_42;
   wire n_64_43;
   wire n_64_44;
   wire n_64_45;
   wire n_64_46;
   wire n_64_47;
   wire n_64_48;
   wire n_64_49;
   wire n_64_50;
   wire n_64_51;
   wire n_64_52;
   wire n_64_53;
   wire n_64_54;
   wire n_64_55;
   wire n_64_56;
   wire n_64_57;
   wire n_64_58;
   wire n_64_59;
   wire n_64_60;
   wire n_64_61;
   wire n_64_62;
   wire n_64_63;
   wire n_64_64;
   wire n_64_65;
   wire n_64_66;
   wire n_64_67;
   wire n_64_68;
   wire n_64_69;
   wire n_64_70;
   wire n_64_71;
   wire n_64_72;
   wire n_64_73;
   wire n_64_74;
   wire n_64_75;
   wire n_64_76;
   wire n_64_77;
   wire n_64_78;
   wire n_64_79;
   wire n_64_80;
   wire n_64_81;
   wire n_64_82;
   wire n_64_83;
   wire n_64_84;
   wire n_64_85;
   wire n_64_86;
   wire n_64_87;
   wire n_64_88;
   wire n_64_89;
   wire n_64_90;
   wire n_64_91;
   wire n_64_92;
   wire n_64_93;
   wire n_64_94;
   wire n_64_95;
   wire n_64_96;
   wire n_64_97;
   wire n_64_98;
   wire n_64_99;
   wire n_64_100;
   wire n_64_101;
   wire n_64_102;
   wire n_64_103;
   wire n_64_104;
   wire n_64_105;
   wire n_64_106;
   wire n_64_107;
   wire n_64_108;
   wire n_64_109;
   wire n_64_110;
   wire n_64_111;
   wire n_64_112;
   wire n_64_113;
   wire n_64_114;
   wire n_64_115;
   wire n_64_116;
   wire n_64_117;
   wire n_64_118;
   wire n_64_119;
   wire n_64_120;
   wire n_64_121;
   wire n_64_122;
   wire n_64_123;
   wire n_64_124;
   wire n_64_125;
   wire n_64_126;
   wire n_64_127;
   wire n_64_128;
   wire n_64_129;
   wire n_64_130;
   wire n_64_131;
   wire n_64_132;
   wire n_64_133;
   wire n_64_134;
   wire n_64_135;
   wire n_64_136;
   wire n_64_137;
   wire n_64_138;
   wire n_64_139;
   wire n_64_140;
   wire n_64_141;
   wire n_64_142;
   wire n_64_143;
   wire n_64_144;
   wire n_64_145;
   wire n_64_146;
   wire n_64_147;
   wire n_64_148;
   wire n_64_149;
   wire n_64_150;
   wire n_64_151;
   wire n_64_152;
   wire n_64_153;
   wire n_64_154;
   wire n_64_155;
   wire n_64_156;
   wire n_64_157;
   wire n_64_158;
   wire n_64_159;
   wire n_64_160;
   wire n_64_161;
   wire n_64_162;
   wire n_64_163;
   wire n_64_164;
   wire n_64_165;
   wire n_64_166;
   wire n_64_167;
   wire n_64_168;
   wire n_64_169;
   wire n_64_170;
   wire n_64_171;
   wire n_64_172;
   wire n_64_173;
   wire n_64_174;
   wire n_64_175;
   wire n_64_176;
   wire n_64_177;
   wire n_64_178;
   wire n_64_179;
   wire n_64_180;
   wire n_64_181;
   wire n_64_182;
   wire n_64_183;
   wire n_64_184;
   wire n_64_185;
   wire n_64_186;
   wire n_64_187;
   wire n_64_188;
   wire n_64_189;
   wire n_64_190;
   wire n_64_191;
   wire n_64_192;
   wire [31:0]A;
   wire [6:0]SC;
   wire [31:0]multiplicand;
   wire [32:0]Q;
   wire out_sign;
   wire n_64_1;
   wire n_64_2;
   wire n_64_1_5;
   wire n_64_1_0;
   wire n_64_1_6;
   wire n_64_1_1;
   wire n_64_1_7;
   wire n_64_1_2;
   wire n_64_1_8;
   wire n_64_1_3;
   wire n_64_1_9;
   wire n_64_1_4;
   wire n_64_193;
   wire n_64_194;
   wire n_64_195;
   wire n_64_196;
   wire n_64_197;
   wire n_64_198;
   wire n_64_199;
   wire n_64_1_10;
   wire n_64_1_11;
   wire n_64_1_12;
   wire n_64_200;
   wire n_64_1_13;
   wire n_64_1_14;
   wire n_64_1_15;
   wire n_64_201;
   wire n_64_1_16;
   wire n_64_202;
   wire n_64_1_17;
   wire n_64_203;
   wire n_64_1_18;
   wire n_64_204;
   wire n_64_1_19;
   wire n_64_205;
   wire n_64_1_20;
   wire n_64_206;
   wire n_64_1_21;
   wire n_64_207;
   wire n_64_1_22;
   wire n_64_208;
   wire n_64_1_23;
   wire n_64_209;
   wire n_64_1_24;
   wire n_64_210;
   wire n_64_1_25;
   wire n_64_211;
   wire n_64_1_26;
   wire n_64_212;
   wire n_64_1_27;
   wire n_64_213;
   wire n_64_1_28;
   wire n_64_214;
   wire n_64_1_29;
   wire n_64_215;
   wire n_64_1_30;
   wire n_64_216;
   wire n_64_1_31;
   wire n_64_217;
   wire n_64_1_32;
   wire n_64_218;
   wire n_64_1_33;
   wire n_64_219;
   wire n_64_1_34;
   wire n_64_220;
   wire n_64_1_35;
   wire n_64_221;
   wire n_64_1_36;
   wire n_64_222;
   wire n_64_1_37;
   wire n_64_223;
   wire n_64_1_38;
   wire n_64_224;
   wire n_64_1_39;
   wire n_64_225;
   wire n_64_1_40;
   wire n_64_226;
   wire n_64_1_41;
   wire n_64_227;
   wire n_64_1_42;
   wire n_64_228;
   wire n_64_1_43;
   wire n_64_229;
   wire n_64_1_44;
   wire n_64_230;
   wire n_64_1_45;
   wire n_64_231;
   wire n_64_1_46;
   wire n_64_232;
   wire n_64_1_47;
   wire n_64_233;
   wire n_64_1_48;
   wire n_64_234;
   wire n_64_1_49;
   wire n_64_235;
   wire n_64_1_50;
   wire n_64_236;
   wire n_64_1_51;
   wire n_64_237;
   wire n_64_1_52;
   wire n_64_238;
   wire n_64_1_53;
   wire n_64_239;
   wire n_64_1_54;
   wire n_64_240;
   wire n_64_1_55;
   wire n_64_241;
   wire n_64_1_56;
   wire n_64_242;
   wire n_64_1_57;
   wire n_64_243;
   wire n_64_1_58;
   wire n_64_244;
   wire n_64_1_59;
   wire n_64_245;
   wire n_64_1_60;
   wire n_64_246;
   wire n_64_1_61;
   wire n_64_247;
   wire n_64_1_62;
   wire n_64_248;
   wire n_64_1_63;
   wire n_64_249;
   wire n_64_1_64;
   wire n_64_250;
   wire n_64_1_65;
   wire n_64_251;
   wire n_64_1_66;
   wire n_64_252;
   wire n_64_1_67;
   wire n_64_253;
   wire n_64_1_68;
   wire n_64_254;
   wire n_64_1_69;
   wire n_64_255;
   wire n_64_1_70;
   wire n_64_256;
   wire n_64_1_71;
   wire n_64_257;
   wire n_64_1_72;
   wire n_64_258;
   wire n_64_1_73;
   wire n_64_259;
   wire n_64_1_74;
   wire n_64_260;
   wire n_64_1_75;
   wire n_64_265;
   wire n_64_266;
   wire n_64_267;
   wire n_64_268;
   wire n_64_269;
   wire n_64_270;
   wire n_64_271;
   wire n_64_272;
   wire n_64_273;
   wire n_64_274;
   wire n_64_275;
   wire n_64_276;
   wire n_64_277;
   wire n_64_278;
   wire n_64_279;
   wire n_64_280;
   wire n_64_281;
   wire n_64_282;
   wire n_64_283;
   wire n_64_284;
   wire n_64_285;
   wire n_64_286;
   wire n_64_287;
   wire n_64_288;
   wire n_64_289;
   wire n_64_290;
   wire n_64_291;
   wire n_64_292;
   wire n_64_293;
   wire n_64_294;
   wire n_64_295;
   wire n_64_296;
   wire n_64_300;
   wire n_64_1_81;
   wire n_64_301;
   wire n_64_1_82;
   wire n_64_302;
   wire n_64_1_83;
   wire n_64_303;
   wire n_64_1_84;
   wire n_64_310;
   wire n_64_1_91;
   wire n_64_311;
   wire n_64_1_92;
   wire n_64_312;
   wire n_64_1_93;
   wire n_64_313;
   wire n_64_1_94;
   wire n_64_314;
   wire n_64_1_95;
   wire n_64_315;
   wire n_64_1_96;
   wire n_64_316;
   wire n_64_1_97;
   wire n_64_317;
   wire n_64_1_98;
   wire n_64_318;
   wire n_64_1_99;
   wire n_64_319;
   wire n_64_1_100;
   wire n_64_320;
   wire n_64_1_101;
   wire n_64_321;
   wire n_64_1_102;
   wire n_64_322;
   wire n_64_1_103;
   wire n_64_323;
   wire n_64_1_104;
   wire n_64_324;
   wire n_64_1_105;
   wire n_64_325;
   wire n_64_1_106;
   wire n_64_326;
   wire n_64_1_107;
   wire n_64_327;
   wire n_64_1_108;
   wire n_64_328;
   wire n_64_1_110;
   wire n_64_1_111;
   wire n_64_329;
   wire n_64_1_113;
   wire n_64_330;
   wire n_64_1_114;
   wire n_64_331;
   wire n_64_1_115;
   wire n_64_332;
   wire n_64_1_116;
   wire n_64_333;
   wire n_64_1_117;
   wire n_64_334;
   wire n_64_1_118;
   wire n_64_335;
   wire n_64_1_119;
   wire n_64_336;
   wire n_64_1_120;
   wire n_64_337;
   wire n_64_1_121;
   wire n_64_338;
   wire n_64_1_122;
   wire n_64_339;
   wire n_64_1_123;
   wire n_64_340;
   wire n_64_1_124;
   wire n_64_341;
   wire n_64_1_125;
   wire n_64_342;
   wire n_64_1_126;
   wire n_64_343;
   wire n_64_1_127;
   wire n_64_344;
   wire n_64_1_128;
   wire n_64_345;
   wire n_64_1_129;
   wire n_64_346;
   wire n_64_1_130;
   wire n_64_347;
   wire n_64_1_131;
   wire n_64_348;
   wire n_64_1_132;
   wire n_64_349;
   wire n_64_1_133;
   wire n_64_350;
   wire n_64_1_134;
   wire n_64_351;
   wire n_64_1_135;
   wire n_64_352;
   wire n_64_1_136;
   wire n_64_353;
   wire n_64_1_137;
   wire n_64_354;
   wire n_64_1_138;
   wire n_64_355;
   wire n_64_1_139;
   wire n_64_356;
   wire n_64_1_140;
   wire n_64_357;
   wire n_64_1_141;
   wire n_64_358;
   wire n_64_1_142;
   wire n_64_359;
   wire n_64_360;
   wire n_64_1_145;
   wire n_64_1_146;
   wire n_64_1_147;
   wire n_64_1_148;
   wire n_64_297;
   wire n_64_1_149;
   wire n_64_361;
   wire n_64_1_150;
   wire n_64_362;
   wire n_64_1_151;
   wire n_64_363;
   wire n_64_1_152;
   wire n_64_364;
   wire n_64_1_153;
   wire n_64_365;
   wire n_64_1_154;
   wire n_64_366;
   wire n_64_1_155;
   wire n_64_367;
   wire n_64_1_156;
   wire n_64_368;
   wire n_64_1_157;
   wire n_64_369;
   wire n_64_1_158;
   wire n_64_370;
   wire n_64_1_159;
   wire n_64_371;
   wire n_64_1_160;
   wire n_64_372;
   wire n_64_1_161;
   wire n_64_373;
   wire n_64_1_162;
   wire n_64_374;
   wire n_64_1_163;
   wire n_64_375;
   wire n_64_1_164;
   wire n_64_376;
   wire n_64_1_165;
   wire n_64_377;
   wire n_64_1_166;
   wire n_64_378;
   wire n_64_1_167;
   wire n_64_379;
   wire n_64_1_168;
   wire n_64_380;
   wire n_64_1_169;
   wire n_64_381;
   wire n_64_1_170;
   wire n_64_382;
   wire n_64_1_171;
   wire n_64_383;
   wire n_64_1_172;
   wire n_64_384;
   wire n_64_1_173;
   wire n_64_385;
   wire n_64_1_174;
   wire n_64_386;
   wire n_64_1_175;
   wire n_64_387;
   wire n_64_1_176;
   wire n_64_388;
   wire n_64_1_177;
   wire n_64_389;
   wire n_64_1_178;
   wire n_64_390;
   wire n_64_1_179;
   wire n_64_391;
   wire n_64_1_180;
   wire n_64_1_181;
   wire n_64_392;
   wire n_64_1_182;
   wire n_64_1_183;
   wire n_64_1_186;
   wire n_64_1_187;
   wire n_64_393;
   wire n_64_394;
   wire n_64_1_188;
   wire n_64_1_189;
   wire n_64_1_190;
   wire n_64_1_191;
   wire n_64_1_192;
   wire n_64_264;
   wire n_64_1_193;
   wire n_64_1_194;
   wire n_64_1_144;
   wire n_64_261;
   wire n_64_1_143;
   wire n_64_1_76;
   wire n_64_262;
   wire n_64_1_77;
   wire n_64_1_79;
   wire n_64_1_195;
   wire n_64_1_196;
   wire n_64_1_197;
   wire n_64_1_198;
   wire n_64_1_199;
   wire n_64_1_200;
   wire n_64_263;
   wire n_64_1_201;
   wire n_64_1_78;
   wire n_64_1_202;
   wire n_64_298;
   wire n_64_1_203;
   wire n_64_1_204;
   wire n_64_299;
   wire n_64_1_80;
   wire n_64_1_205;
   wire n_64_304;
   wire n_64_1_85;
   wire n_64_1_206;
   wire n_64_305;
   wire n_64_1_86;
   wire n_64_1_207;
   wire n_64_306;
   wire n_64_1_87;
   wire n_64_1_208;
   wire n_64_307;
   wire n_64_1_88;
   wire n_64_1_209;
   wire n_64_308;
   wire n_64_1_89;
   wire n_64_1_210;
   wire n_64_309;
   wire n_64_1_90;
   wire n_64_1_211;
   wire n_64_1_109;
   wire n_64_1_212;
   wire n_64_1_112;
   wire n_64_1_184;
   wire n_64_1_185;

   TBUF_X1 i_0 (.A(n_64), .EN(n_0), .Z(c[0]));
   TBUF_X1 i_1 (.A(n_63), .EN(n_0), .Z(c[1]));
   TBUF_X1 i_2 (.A(n_62), .EN(n_0), .Z(c[2]));
   TBUF_X1 i_3 (.A(n_61), .EN(n_0), .Z(c[3]));
   TBUF_X1 i_4 (.A(n_60), .EN(n_0), .Z(c[4]));
   TBUF_X1 i_5 (.A(n_59), .EN(n_0), .Z(c[5]));
   TBUF_X1 i_6 (.A(n_58), .EN(n_0), .Z(c[6]));
   TBUF_X1 i_7 (.A(n_57), .EN(n_0), .Z(c[7]));
   TBUF_X1 i_8 (.A(n_56), .EN(n_0), .Z(c[8]));
   TBUF_X1 i_9 (.A(n_55), .EN(n_0), .Z(c[9]));
   TBUF_X1 i_10 (.A(n_54), .EN(n_0), .Z(c[10]));
   TBUF_X1 i_11 (.A(n_53), .EN(n_0), .Z(c[11]));
   TBUF_X1 i_12 (.A(n_52), .EN(n_0), .Z(c[12]));
   TBUF_X1 i_13 (.A(n_51), .EN(n_0), .Z(c[13]));
   TBUF_X1 i_14 (.A(n_50), .EN(n_0), .Z(c[14]));
   TBUF_X1 i_15 (.A(n_49), .EN(n_0), .Z(c[15]));
   TBUF_X1 i_16 (.A(n_48), .EN(n_0), .Z(c[16]));
   TBUF_X1 i_17 (.A(n_47), .EN(n_0), .Z(c[17]));
   TBUF_X1 i_18 (.A(n_46), .EN(n_0), .Z(c[18]));
   TBUF_X1 i_19 (.A(n_45), .EN(n_0), .Z(c[19]));
   TBUF_X1 i_20 (.A(n_44), .EN(n_0), .Z(c[20]));
   TBUF_X1 i_21 (.A(n_43), .EN(n_0), .Z(c[21]));
   TBUF_X1 i_22 (.A(n_42), .EN(n_0), .Z(c[22]));
   TBUF_X1 i_23 (.A(n_41), .EN(n_0), .Z(c[23]));
   TBUF_X1 i_24 (.A(n_40), .EN(n_0), .Z(c[24]));
   TBUF_X1 i_25 (.A(n_39), .EN(n_0), .Z(c[25]));
   TBUF_X1 i_26 (.A(n_38), .EN(n_0), .Z(c[26]));
   TBUF_X1 i_27 (.A(n_37), .EN(n_0), .Z(c[27]));
   TBUF_X1 i_28 (.A(n_36), .EN(n_0), .Z(c[28]));
   TBUF_X1 i_29 (.A(n_35), .EN(n_0), .Z(c[29]));
   TBUF_X1 i_30 (.A(n_34), .EN(n_0), .Z(c[30]));
   TBUF_X1 i_31 (.A(n_33), .EN(n_0), .Z(c[31]));
   TBUF_X1 i_32 (.A(n_32), .EN(n_0), .Z(c[32]));
   TBUF_X1 i_33 (.A(n_31), .EN(n_0), .Z(c[33]));
   TBUF_X1 i_34 (.A(n_30), .EN(n_0), .Z(c[34]));
   TBUF_X1 i_35 (.A(n_29), .EN(n_0), .Z(c[35]));
   TBUF_X1 i_36 (.A(n_28), .EN(n_0), .Z(c[36]));
   TBUF_X1 i_37 (.A(n_27), .EN(n_0), .Z(c[37]));
   TBUF_X1 i_38 (.A(n_26), .EN(n_0), .Z(c[38]));
   TBUF_X1 i_39 (.A(n_25), .EN(n_0), .Z(c[39]));
   TBUF_X1 i_40 (.A(n_24), .EN(n_0), .Z(c[40]));
   TBUF_X1 i_41 (.A(n_23), .EN(n_0), .Z(c[41]));
   TBUF_X1 i_42 (.A(n_22), .EN(n_0), .Z(c[42]));
   TBUF_X1 i_43 (.A(n_21), .EN(n_0), .Z(c[43]));
   TBUF_X1 i_44 (.A(n_20), .EN(n_0), .Z(c[44]));
   TBUF_X1 i_45 (.A(n_19), .EN(n_0), .Z(c[45]));
   TBUF_X1 i_46 (.A(n_18), .EN(n_0), .Z(c[46]));
   TBUF_X1 i_47 (.A(n_17), .EN(n_0), .Z(c[47]));
   TBUF_X1 i_48 (.A(n_16), .EN(n_0), .Z(c[48]));
   TBUF_X1 i_49 (.A(n_15), .EN(n_0), .Z(c[49]));
   TBUF_X1 i_50 (.A(n_14), .EN(n_0), .Z(c[50]));
   TBUF_X1 i_51 (.A(n_13), .EN(n_0), .Z(c[51]));
   TBUF_X1 i_52 (.A(n_12), .EN(n_0), .Z(c[52]));
   TBUF_X1 i_53 (.A(n_11), .EN(n_0), .Z(c[53]));
   TBUF_X1 i_54 (.A(n_10), .EN(n_0), .Z(c[54]));
   TBUF_X1 i_55 (.A(n_9), .EN(n_0), .Z(c[55]));
   TBUF_X1 i_56 (.A(n_8), .EN(n_0), .Z(c[56]));
   TBUF_X1 i_57 (.A(n_7), .EN(n_0), .Z(c[57]));
   TBUF_X1 i_58 (.A(n_6), .EN(n_0), .Z(c[58]));
   TBUF_X1 i_59 (.A(n_5), .EN(n_0), .Z(c[59]));
   TBUF_X1 i_60 (.A(n_4), .EN(n_0), .Z(c[60]));
   TBUF_X1 i_61 (.A(n_3), .EN(n_0), .Z(c[61]));
   TBUF_X1 i_62 (.A(n_2), .EN(n_0), .Z(c[62]));
   TBUF_X1 i_63 (.A(n_1), .EN(n_0), .Z(c[63]));
   INV_X1 i_64_0 (.A(n_64_3), .ZN(n_0));
   CLKGATETST_X1 clk_gate_c_reg (.CK(clk), .E(n_64_393), .SE(1'b0), .GCK(n_64_0));
   DFF_X1 \c_reg[63]  (.D(n_64_263), .CK(n_64_0), .Q(n_1), .QN());
   DFF_X1 \c_reg[62]  (.D(n_64_262), .CK(n_64_0), .Q(n_2), .QN());
   DFF_X1 \c_reg[61]  (.D(n_64_261), .CK(n_64_0), .Q(n_3), .QN());
   DFF_X1 \c_reg[60]  (.D(n_64_260), .CK(n_64_0), .Q(n_4), .QN());
   DFF_X1 \c_reg[59]  (.D(n_64_259), .CK(n_64_0), .Q(n_5), .QN());
   DFF_X1 \c_reg[58]  (.D(n_64_258), .CK(n_64_0), .Q(n_6), .QN());
   DFF_X1 \c_reg[57]  (.D(n_64_257), .CK(n_64_0), .Q(n_7), .QN());
   DFF_X1 \c_reg[56]  (.D(n_64_256), .CK(n_64_0), .Q(n_8), .QN());
   DFF_X1 \c_reg[55]  (.D(n_64_255), .CK(n_64_0), .Q(n_9), .QN());
   DFF_X1 \c_reg[54]  (.D(n_64_254), .CK(n_64_0), .Q(n_10), .QN());
   DFF_X1 \c_reg[53]  (.D(n_64_253), .CK(n_64_0), .Q(n_11), .QN());
   DFF_X1 \c_reg[52]  (.D(n_64_252), .CK(n_64_0), .Q(n_12), .QN());
   DFF_X1 \c_reg[51]  (.D(n_64_251), .CK(n_64_0), .Q(n_13), .QN());
   DFF_X1 \c_reg[50]  (.D(n_64_250), .CK(n_64_0), .Q(n_14), .QN());
   DFF_X1 \c_reg[49]  (.D(n_64_249), .CK(n_64_0), .Q(n_15), .QN());
   DFF_X1 \c_reg[48]  (.D(n_64_248), .CK(n_64_0), .Q(n_16), .QN());
   DFF_X1 \c_reg[47]  (.D(n_64_247), .CK(n_64_0), .Q(n_17), .QN());
   DFF_X1 \c_reg[46]  (.D(n_64_246), .CK(n_64_0), .Q(n_18), .QN());
   DFF_X1 \c_reg[45]  (.D(n_64_245), .CK(n_64_0), .Q(n_19), .QN());
   DFF_X1 \c_reg[44]  (.D(n_64_244), .CK(n_64_0), .Q(n_20), .QN());
   DFF_X1 \c_reg[43]  (.D(n_64_243), .CK(n_64_0), .Q(n_21), .QN());
   DFF_X1 \c_reg[42]  (.D(n_64_242), .CK(n_64_0), .Q(n_22), .QN());
   DFF_X1 \c_reg[41]  (.D(n_64_241), .CK(n_64_0), .Q(n_23), .QN());
   DFF_X1 \c_reg[40]  (.D(n_64_240), .CK(n_64_0), .Q(n_24), .QN());
   DFF_X1 \c_reg[39]  (.D(n_64_239), .CK(n_64_0), .Q(n_25), .QN());
   DFF_X1 \c_reg[38]  (.D(n_64_238), .CK(n_64_0), .Q(n_26), .QN());
   DFF_X1 \c_reg[37]  (.D(n_64_237), .CK(n_64_0), .Q(n_27), .QN());
   DFF_X1 \c_reg[36]  (.D(n_64_236), .CK(n_64_0), .Q(n_28), .QN());
   DFF_X1 \c_reg[35]  (.D(n_64_235), .CK(n_64_0), .Q(n_29), .QN());
   DFF_X1 \c_reg[34]  (.D(n_64_234), .CK(n_64_0), .Q(n_30), .QN());
   DFF_X1 \c_reg[33]  (.D(n_64_233), .CK(n_64_0), .Q(n_31), .QN());
   DFF_X1 \c_reg[32]  (.D(n_64_232), .CK(n_64_0), .Q(n_32), .QN());
   DFF_X1 \c_reg[31]  (.D(n_64_231), .CK(n_64_0), .Q(n_33), .QN());
   DFF_X1 \c_reg[30]  (.D(n_64_230), .CK(n_64_0), .Q(n_34), .QN());
   DFF_X1 \c_reg[29]  (.D(n_64_229), .CK(n_64_0), .Q(n_35), .QN());
   DFF_X1 \c_reg[28]  (.D(n_64_228), .CK(n_64_0), .Q(n_36), .QN());
   DFF_X1 \c_reg[27]  (.D(n_64_227), .CK(n_64_0), .Q(n_37), .QN());
   DFF_X1 \c_reg[26]  (.D(n_64_226), .CK(n_64_0), .Q(n_38), .QN());
   DFF_X1 \c_reg[25]  (.D(n_64_225), .CK(n_64_0), .Q(n_39), .QN());
   DFF_X1 \c_reg[24]  (.D(n_64_224), .CK(n_64_0), .Q(n_40), .QN());
   DFF_X1 \c_reg[23]  (.D(n_64_223), .CK(n_64_0), .Q(n_41), .QN());
   DFF_X1 \c_reg[22]  (.D(n_64_222), .CK(n_64_0), .Q(n_42), .QN());
   DFF_X1 \c_reg[21]  (.D(n_64_221), .CK(n_64_0), .Q(n_43), .QN());
   DFF_X1 \c_reg[20]  (.D(n_64_220), .CK(n_64_0), .Q(n_44), .QN());
   DFF_X1 \c_reg[19]  (.D(n_64_219), .CK(n_64_0), .Q(n_45), .QN());
   DFF_X1 \c_reg[18]  (.D(n_64_218), .CK(n_64_0), .Q(n_46), .QN());
   DFF_X1 \c_reg[17]  (.D(n_64_217), .CK(n_64_0), .Q(n_47), .QN());
   DFF_X1 \c_reg[16]  (.D(n_64_216), .CK(n_64_0), .Q(n_48), .QN());
   DFF_X1 \c_reg[15]  (.D(n_64_215), .CK(n_64_0), .Q(n_49), .QN());
   DFF_X1 \c_reg[14]  (.D(n_64_214), .CK(n_64_0), .Q(n_50), .QN());
   DFF_X1 \c_reg[13]  (.D(n_64_213), .CK(n_64_0), .Q(n_51), .QN());
   DFF_X1 \c_reg[12]  (.D(n_64_212), .CK(n_64_0), .Q(n_52), .QN());
   DFF_X1 \c_reg[11]  (.D(n_64_211), .CK(n_64_0), .Q(n_53), .QN());
   DFF_X1 \c_reg[10]  (.D(n_64_210), .CK(n_64_0), .Q(n_54), .QN());
   DFF_X1 \c_reg[9]  (.D(n_64_209), .CK(n_64_0), .Q(n_55), .QN());
   DFF_X1 \c_reg[8]  (.D(n_64_208), .CK(n_64_0), .Q(n_56), .QN());
   DFF_X1 \c_reg[7]  (.D(n_64_207), .CK(n_64_0), .Q(n_57), .QN());
   DFF_X1 \c_reg[6]  (.D(n_64_206), .CK(n_64_0), .Q(n_58), .QN());
   DFF_X1 \c_reg[5]  (.D(n_64_205), .CK(n_64_0), .Q(n_59), .QN());
   DFF_X1 \c_reg[4]  (.D(n_64_204), .CK(n_64_0), .Q(n_60), .QN());
   DFF_X1 \c_reg[3]  (.D(n_64_203), .CK(n_64_0), .Q(n_61), .QN());
   DFF_X1 \c_reg[2]  (.D(n_64_202), .CK(n_64_0), .Q(n_62), .QN());
   DFF_X1 \c_reg[1]  (.D(n_64_201), .CK(n_64_0), .Q(n_63), .QN());
   DFF_X1 \c_reg[0]  (.D(n_64_298), .CK(n_64_0), .Q(n_64), .QN());
   DFF_X1 i_64_64 (.D(n_64_394), .CK(clk), .Q(n_64_3), .QN());
   datapath i_64_194 (.p_0({n_64_34, n_64_33, n_64_32, n_64_31, n_64_30, n_64_29, 
      n_64_28, n_64_27, n_64_26, n_64_25, n_64_24, n_64_23, n_64_22, n_64_21, 
      n_64_20, n_64_19, n_64_18, n_64_17, n_64_16, n_64_15, n_64_14, n_64_13, 
      n_64_12, n_64_11, n_64_10, n_64_9, n_64_8, n_64_7, n_64_6, n_64_5, n_64_4, 
      uc_0}), .a(a));
   datapath__0_65 i_64_196 (.A({A[31], uc_1, A[29], A[28], A[27], A[26], A[25], 
      A[24], A[23], A[22], A[21], A[20], A[19], A[18], A[17], A[16], A[15], 
      A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], 
      A[3], A[2], A[1], A[0]}), .p_0({n_64_66, n_64_65, n_64_64, n_64_63, 
      n_64_62, n_64_61, n_64_60, n_64_59, n_64_58, n_64_57, n_64_56, n_64_55, 
      n_64_54, n_64_53, n_64_52, n_64_51, n_64_50, n_64_49, n_64_48, n_64_47, 
      n_64_46, n_64_45, n_64_44, n_64_43, n_64_42, n_64_41, n_64_40, n_64_39, 
      n_64_38, n_64_37, n_64_36, n_64_35}), .multiplicand({n_64_392, n_64_391, 
      n_64_390, n_64_389, n_64_388, n_64_387, n_64_386, n_64_385, n_64_384, 
      n_64_383, n_64_382, n_64_381, n_64_380, n_64_379, n_64_378, n_64_377, 
      n_64_376, n_64_375, n_64_374, n_64_373, n_64_372, n_64_371, n_64_370, 
      n_64_369, n_64_368, n_64_367, n_64_366, n_64_365, n_64_364, n_64_363, 
      n_64_362, n_64_361}));
   datapath__0_66 i_64_197 (.multiplicand({n_64_392, n_64_391, n_64_390, 
      n_64_389, n_64_388, n_64_387, n_64_386, n_64_385, n_64_384, n_64_383, 
      n_64_382, n_64_381, n_64_380, n_64_379, n_64_378, n_64_377, n_64_376, 
      n_64_375, n_64_374, n_64_373, n_64_372, n_64_371, n_64_370, n_64_369, 
      n_64_368, n_64_367, n_64_366, n_64_365, n_64_364, n_64_363, n_64_362, 
      n_64_361}), .A({A[31], uc_2, A[29], A[28], A[27], A[26], A[25], A[24], 
      A[23], A[22], A[21], A[20], A[19], A[18], A[17], A[16], A[15], A[14], 
      A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], 
      A[1], A[0]}), .p_0({n_64_98, n_64_97, n_64_96, n_64_95, n_64_94, n_64_93, 
      n_64_92, n_64_91, n_64_90, n_64_89, n_64_88, n_64_87, n_64_86, n_64_85, 
      n_64_84, n_64_83, n_64_82, n_64_81, n_64_80, n_64_79, n_64_78, n_64_77, 
      n_64_76, n_64_75, n_64_74, n_64_73, n_64_72, n_64_71, n_64_70, n_64_69, 
      n_64_68, n_64_67}));
   datapath__0_67 i_64_198 (.p_0({n_64_129, n_64_128, n_64_127, n_64_126, 
      n_64_125, n_64_124, n_64_123, n_64_122, n_64_121, n_64_120, n_64_119, 
      n_64_118, n_64_117, n_64_116, n_64_115, n_64_114, n_64_113, n_64_112, 
      n_64_111, n_64_110, n_64_109, n_64_108, n_64_107, n_64_106, n_64_105, 
      n_64_104, n_64_103, n_64_102, n_64_101, n_64_100, n_64_99, uc_3}), 
      .b(b));
   datapath__0_72 i_64_203 (.p_0({n_64_192, n_64_191, n_64_190, n_64_189, 
      n_64_188, n_64_187, n_64_186, n_64_185, n_64_184, n_64_183, n_64_182, 
      n_64_181, n_64_180, n_64_179, n_64_178, n_64_177, n_64_176, n_64_175, 
      n_64_174, n_64_173, n_64_172, n_64_171, n_64_170, n_64_169, n_64_168, 
      n_64_167, n_64_166, n_64_165, n_64_164, n_64_163, n_64_162, n_64_161, 
      n_64_160, n_64_159, n_64_158, n_64_157, n_64_156, n_64_155, n_64_154, 
      n_64_153, n_64_152, n_64_151, n_64_150, n_64_149, n_64_148, n_64_147, 
      n_64_146, n_64_145, n_64_144, n_64_143, n_64_142, n_64_141, n_64_140, 
      n_64_139, n_64_138, n_64_137, n_64_136, n_64_135, n_64_134, n_64_133, 
      n_64_132, n_64_131, n_64_130, uc_4}), .p_1({uc_5, n_64_360, n_64_359, 
      n_64_358, n_64_357, n_64_356, n_64_355, n_64_354, n_64_353, n_64_352, 
      n_64_351, n_64_350, n_64_349, n_64_348, n_64_347, n_64_346, n_64_345, 
      n_64_344, n_64_343, n_64_342, n_64_341, n_64_340, n_64_339, n_64_338, 
      n_64_337, n_64_336, n_64_335, n_64_334, n_64_333, n_64_332, n_64_331, 
      n_64_330, n_64_329, n_64_328, n_64_327, n_64_326, n_64_325, n_64_324, 
      n_64_323, n_64_322, n_64_321, n_64_320, n_64_319, n_64_318, n_64_317, 
      n_64_316, n_64_315, n_64_314, n_64_313, n_64_312, n_64_311, n_64_310, 
      n_64_309, n_64_308, n_64_307, n_64_306, n_64_305, n_64_304, n_64_303, 
      n_64_302, n_64_301, n_64_300, n_64_299, n_64_298}));
   DFF_X1 \A_reg[31]  (.D(n_64_295), .CK(n_64_1), .Q(A[31]), .QN());
   DFF_X1 \A_reg[29]  (.D(n_64_294), .CK(n_64_1), .Q(A[29]), .QN());
   DFF_X1 \A_reg[28]  (.D(n_64_293), .CK(n_64_1), .Q(A[28]), .QN());
   DFF_X1 \A_reg[27]  (.D(n_64_292), .CK(n_64_1), .Q(A[27]), .QN());
   DFF_X1 \A_reg[26]  (.D(n_64_291), .CK(n_64_1), .Q(A[26]), .QN());
   DFF_X1 \A_reg[25]  (.D(n_64_290), .CK(n_64_1), .Q(A[25]), .QN());
   DFF_X1 \A_reg[24]  (.D(n_64_289), .CK(n_64_1), .Q(A[24]), .QN());
   DFF_X1 \A_reg[23]  (.D(n_64_288), .CK(n_64_1), .Q(A[23]), .QN());
   DFF_X1 \A_reg[22]  (.D(n_64_287), .CK(n_64_1), .Q(A[22]), .QN());
   DFF_X1 \A_reg[21]  (.D(n_64_286), .CK(n_64_1), .Q(A[21]), .QN());
   DFF_X1 \A_reg[20]  (.D(n_64_285), .CK(n_64_1), .Q(A[20]), .QN());
   DFF_X1 \A_reg[19]  (.D(n_64_284), .CK(n_64_1), .Q(A[19]), .QN());
   DFF_X1 \A_reg[18]  (.D(n_64_283), .CK(n_64_1), .Q(A[18]), .QN());
   DFF_X1 \A_reg[17]  (.D(n_64_282), .CK(n_64_1), .Q(A[17]), .QN());
   DFF_X1 \A_reg[16]  (.D(n_64_281), .CK(n_64_1), .Q(A[16]), .QN());
   DFF_X1 \A_reg[15]  (.D(n_64_280), .CK(n_64_1), .Q(A[15]), .QN());
   DFF_X1 \A_reg[14]  (.D(n_64_279), .CK(n_64_1), .Q(A[14]), .QN());
   DFF_X1 \A_reg[13]  (.D(n_64_278), .CK(n_64_1), .Q(A[13]), .QN());
   DFF_X1 \A_reg[12]  (.D(n_64_277), .CK(n_64_1), .Q(A[12]), .QN());
   DFF_X1 \A_reg[11]  (.D(n_64_276), .CK(n_64_1), .Q(A[11]), .QN());
   DFF_X1 \A_reg[10]  (.D(n_64_275), .CK(n_64_1), .Q(A[10]), .QN());
   DFF_X1 \A_reg[9]  (.D(n_64_274), .CK(n_64_1), .Q(A[9]), .QN());
   DFF_X1 \A_reg[8]  (.D(n_64_273), .CK(n_64_1), .Q(A[8]), .QN());
   DFF_X1 \A_reg[7]  (.D(n_64_272), .CK(n_64_1), .Q(A[7]), .QN());
   DFF_X1 \A_reg[6]  (.D(n_64_271), .CK(n_64_1), .Q(A[6]), .QN());
   DFF_X1 \A_reg[5]  (.D(n_64_270), .CK(n_64_1), .Q(A[5]), .QN());
   DFF_X1 \A_reg[4]  (.D(n_64_269), .CK(n_64_1), .Q(A[4]), .QN());
   DFF_X1 \A_reg[3]  (.D(n_64_268), .CK(n_64_1), .Q(A[3]), .QN());
   DFF_X1 \A_reg[2]  (.D(n_64_267), .CK(n_64_1), .Q(A[2]), .QN());
   DFF_X1 \A_reg[1]  (.D(n_64_266), .CK(n_64_1), .Q(A[1]), .QN());
   DFF_X1 \A_reg[0]  (.D(n_64_265), .CK(n_64_1), .Q(A[0]), .QN());
   DFF_X1 \SC_reg[6]  (.D(n_64_199), .CK(n_64_1), .Q(SC[6]), .QN());
   DFF_X1 \SC_reg[5]  (.D(n_64_198), .CK(n_64_1), .Q(SC[5]), .QN());
   DFF_X1 \SC_reg[4]  (.D(n_64_197), .CK(n_64_1), .Q(SC[4]), .QN());
   DFF_X1 \SC_reg[3]  (.D(n_64_196), .CK(n_64_1), .Q(SC[3]), .QN());
   DFF_X1 \SC_reg[2]  (.D(n_64_195), .CK(n_64_1), .Q(SC[2]), .QN());
   DFF_X1 \SC_reg[1]  (.D(n_64_194), .CK(n_64_1), .Q(SC[1]), .QN());
   DFF_X1 \SC_reg[0]  (.D(n_64_193), .CK(n_64_1), .Q(SC[0]), .QN());
   DFF_X1 \multiplicand_reg[31]  (.D(n_64_392), .CK(n_64_2), .Q(multiplicand[31]), 
      .QN());
   DFF_X1 \multiplicand_reg[30]  (.D(n_64_391), .CK(n_64_2), .Q(multiplicand[30]), 
      .QN());
   DFF_X1 \multiplicand_reg[29]  (.D(n_64_390), .CK(n_64_2), .Q(multiplicand[29]), 
      .QN());
   DFF_X1 \multiplicand_reg[28]  (.D(n_64_389), .CK(n_64_2), .Q(multiplicand[28]), 
      .QN());
   DFF_X1 \multiplicand_reg[27]  (.D(n_64_388), .CK(n_64_2), .Q(multiplicand[27]), 
      .QN());
   DFF_X1 \multiplicand_reg[26]  (.D(n_64_387), .CK(n_64_2), .Q(multiplicand[26]), 
      .QN());
   DFF_X1 \multiplicand_reg[25]  (.D(n_64_386), .CK(n_64_2), .Q(multiplicand[25]), 
      .QN());
   DFF_X1 \multiplicand_reg[24]  (.D(n_64_385), .CK(n_64_2), .Q(multiplicand[24]), 
      .QN());
   DFF_X1 \multiplicand_reg[23]  (.D(n_64_384), .CK(n_64_2), .Q(multiplicand[23]), 
      .QN());
   DFF_X1 \multiplicand_reg[22]  (.D(n_64_383), .CK(n_64_2), .Q(multiplicand[22]), 
      .QN());
   DFF_X1 \multiplicand_reg[21]  (.D(n_64_382), .CK(n_64_2), .Q(multiplicand[21]), 
      .QN());
   DFF_X1 \multiplicand_reg[20]  (.D(n_64_381), .CK(n_64_2), .Q(multiplicand[20]), 
      .QN());
   DFF_X1 \multiplicand_reg[19]  (.D(n_64_380), .CK(n_64_2), .Q(multiplicand[19]), 
      .QN());
   DFF_X1 \multiplicand_reg[18]  (.D(n_64_379), .CK(n_64_2), .Q(multiplicand[18]), 
      .QN());
   DFF_X1 \multiplicand_reg[17]  (.D(n_64_378), .CK(n_64_2), .Q(multiplicand[17]), 
      .QN());
   DFF_X1 \multiplicand_reg[16]  (.D(n_64_377), .CK(n_64_2), .Q(multiplicand[16]), 
      .QN());
   DFF_X1 \multiplicand_reg[15]  (.D(n_64_376), .CK(n_64_2), .Q(multiplicand[15]), 
      .QN());
   DFF_X1 \multiplicand_reg[14]  (.D(n_64_375), .CK(n_64_2), .Q(multiplicand[14]), 
      .QN());
   DFF_X1 \multiplicand_reg[13]  (.D(n_64_374), .CK(n_64_2), .Q(multiplicand[13]), 
      .QN());
   DFF_X1 \multiplicand_reg[12]  (.D(n_64_373), .CK(n_64_2), .Q(multiplicand[12]), 
      .QN());
   DFF_X1 \multiplicand_reg[11]  (.D(n_64_372), .CK(n_64_2), .Q(multiplicand[11]), 
      .QN());
   DFF_X1 \multiplicand_reg[10]  (.D(n_64_371), .CK(n_64_2), .Q(multiplicand[10]), 
      .QN());
   DFF_X1 \multiplicand_reg[9]  (.D(n_64_370), .CK(n_64_2), .Q(multiplicand[9]), 
      .QN());
   DFF_X1 \multiplicand_reg[8]  (.D(n_64_369), .CK(n_64_2), .Q(multiplicand[8]), 
      .QN());
   DFF_X1 \multiplicand_reg[7]  (.D(n_64_368), .CK(n_64_2), .Q(multiplicand[7]), 
      .QN());
   DFF_X1 \multiplicand_reg[6]  (.D(n_64_367), .CK(n_64_2), .Q(multiplicand[6]), 
      .QN());
   DFF_X1 \multiplicand_reg[5]  (.D(n_64_366), .CK(n_64_2), .Q(multiplicand[5]), 
      .QN());
   DFF_X1 \multiplicand_reg[4]  (.D(n_64_365), .CK(n_64_2), .Q(multiplicand[4]), 
      .QN());
   DFF_X1 \multiplicand_reg[3]  (.D(n_64_364), .CK(n_64_2), .Q(multiplicand[3]), 
      .QN());
   DFF_X1 \multiplicand_reg[2]  (.D(n_64_363), .CK(n_64_2), .Q(multiplicand[2]), 
      .QN());
   DFF_X1 \multiplicand_reg[1]  (.D(n_64_362), .CK(n_64_2), .Q(multiplicand[1]), 
      .QN());
   DFF_X1 \multiplicand_reg[0]  (.D(n_64_361), .CK(n_64_2), .Q(multiplicand[0]), 
      .QN());
   DFF_X1 \Q_reg[32]  (.D(n_64_329), .CK(n_64_2), .Q(Q[32]), .QN());
   DFF_X1 \Q_reg[31]  (.D(n_64_328), .CK(n_64_2), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_64_327), .CK(n_64_2), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_64_326), .CK(n_64_2), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_64_325), .CK(n_64_2), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_64_324), .CK(n_64_2), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_64_323), .CK(n_64_2), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_64_322), .CK(n_64_2), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_64_321), .CK(n_64_2), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_64_320), .CK(n_64_2), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_64_319), .CK(n_64_2), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_64_318), .CK(n_64_2), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_64_317), .CK(n_64_2), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_64_316), .CK(n_64_2), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_64_315), .CK(n_64_2), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_64_314), .CK(n_64_2), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_64_313), .CK(n_64_2), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_64_312), .CK(n_64_2), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_64_311), .CK(n_64_2), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_64_310), .CK(n_64_2), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_64_309), .CK(n_64_2), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_64_308), .CK(n_64_2), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_64_307), .CK(n_64_2), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_64_306), .CK(n_64_2), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_64_305), .CK(n_64_2), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_64_304), .CK(n_64_2), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_64_303), .CK(n_64_2), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_64_302), .CK(n_64_2), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_64_301), .CK(n_64_2), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_64_300), .CK(n_64_2), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_64_299), .CK(n_64_2), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_64_298), .CK(n_64_2), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_64_297), .CK(n_64_2), .Q(Q[0]), .QN());
   DFF_X1 out_sign_reg (.D(n_64_200), .CK(n_64_2), .Q(out_sign), .QN());
   CLKGATETST_X1 clk_gate_SC_reg (.CK(clk), .E(n_64_296), .SE(1'b0), .GCK(n_64_1));
   CLKGATETST_X1 clk_gate_out_sign_reg (.CK(clk), .E(n_64_264), .SE(1'b0), 
      .GCK(n_64_2));
   HA_X1 i_64_1_0 (.A(SC[1]), .B(SC[0]), .CO(n_64_1_0), .S(n_64_1_5));
   HA_X1 i_64_1_1 (.A(SC[2]), .B(n_64_1_0), .CO(n_64_1_1), .S(n_64_1_6));
   HA_X1 i_64_1_2 (.A(SC[3]), .B(n_64_1_1), .CO(n_64_1_2), .S(n_64_1_7));
   HA_X1 i_64_1_3 (.A(SC[4]), .B(n_64_1_2), .CO(n_64_1_3), .S(n_64_1_8));
   HA_X1 i_64_1_4 (.A(SC[5]), .B(n_64_1_3), .CO(n_64_1_4), .S(n_64_1_9));
   NOR2_X1 i_64_1_5 (.A1(rst), .A2(SC[0]), .ZN(n_64_193));
   AND2_X1 i_64_1_6 (.A1(n_64_1_5), .A2(n_64_1_12), .ZN(n_64_194));
   AND2_X1 i_64_1_7 (.A1(n_64_1_6), .A2(n_64_1_12), .ZN(n_64_195));
   AND2_X1 i_64_1_8 (.A1(n_64_1_7), .A2(n_64_1_12), .ZN(n_64_196));
   AND2_X1 i_64_1_9 (.A1(n_64_1_8), .A2(n_64_1_12), .ZN(n_64_197));
   AND2_X1 i_64_1_10 (.A1(n_64_1_9), .A2(n_64_1_12), .ZN(n_64_198));
   INV_X1 i_64_1_11 (.A(n_64_1_10), .ZN(n_64_199));
   OAI211_X1 i_64_1_12 (.A(n_64_1_12), .B(n_64_1_11), .C1(SC[6]), .C2(n_64_1_4), 
      .ZN(n_64_1_10));
   NAND2_X1 i_64_1_13 (.A1(SC[6]), .A2(n_64_1_4), .ZN(n_64_1_11));
   OAI21_X1 i_64_1_14 (.A(n_64_296), .B1(rst), .B2(n_64_1_190), .ZN(n_64_1_12));
   AOI21_X1 i_64_1_15 (.A(n_64_1_15), .B1(en), .B2(n_64_1_13), .ZN(n_64_200));
   OAI21_X1 i_64_1_16 (.A(n_64_1_14), .B1(a[31]), .B2(n_64_1_109), .ZN(n_64_1_13));
   NAND2_X1 i_64_1_17 (.A1(b[31]), .A2(n_64_1_183), .ZN(n_64_1_14));
   AOI21_X1 i_64_1_18 (.A(out_sign), .B1(en), .B2(n_64_1_184), .ZN(n_64_1_15));
   OAI21_X1 i_64_1_19 (.A(n_64_1_16), .B1(n_64_1_80), .B2(n_64_1_78), .ZN(
      n_64_201));
   NAND2_X1 i_64_1_20 (.A1(n_64_130), .A2(n_64_1_78), .ZN(n_64_1_16));
   OAI21_X1 i_64_1_21 (.A(n_64_1_17), .B1(n_64_1_81), .B2(n_64_1_78), .ZN(
      n_64_202));
   NAND2_X1 i_64_1_22 (.A1(n_64_131), .A2(n_64_1_78), .ZN(n_64_1_17));
   OAI21_X1 i_64_1_23 (.A(n_64_1_18), .B1(n_64_1_82), .B2(n_64_1_78), .ZN(
      n_64_203));
   NAND2_X1 i_64_1_24 (.A1(n_64_132), .A2(n_64_1_78), .ZN(n_64_1_18));
   OAI21_X1 i_64_1_25 (.A(n_64_1_19), .B1(n_64_1_83), .B2(n_64_1_78), .ZN(
      n_64_204));
   NAND2_X1 i_64_1_26 (.A1(n_64_133), .A2(n_64_1_78), .ZN(n_64_1_19));
   OAI21_X1 i_64_1_27 (.A(n_64_1_20), .B1(n_64_1_84), .B2(n_64_1_78), .ZN(
      n_64_205));
   NAND2_X1 i_64_1_28 (.A1(n_64_134), .A2(n_64_1_78), .ZN(n_64_1_20));
   OAI21_X1 i_64_1_29 (.A(n_64_1_21), .B1(n_64_1_85), .B2(n_64_1_78), .ZN(
      n_64_206));
   NAND2_X1 i_64_1_30 (.A1(n_64_135), .A2(n_64_1_78), .ZN(n_64_1_21));
   OAI21_X1 i_64_1_31 (.A(n_64_1_22), .B1(n_64_1_86), .B2(n_64_1_78), .ZN(
      n_64_207));
   NAND2_X1 i_64_1_32 (.A1(n_64_136), .A2(n_64_1_78), .ZN(n_64_1_22));
   OAI21_X1 i_64_1_33 (.A(n_64_1_23), .B1(n_64_1_87), .B2(n_64_1_78), .ZN(
      n_64_208));
   NAND2_X1 i_64_1_34 (.A1(n_64_137), .A2(n_64_1_78), .ZN(n_64_1_23));
   OAI21_X1 i_64_1_35 (.A(n_64_1_24), .B1(n_64_1_88), .B2(n_64_1_78), .ZN(
      n_64_209));
   NAND2_X1 i_64_1_36 (.A1(n_64_138), .A2(n_64_1_78), .ZN(n_64_1_24));
   OAI21_X1 i_64_1_37 (.A(n_64_1_25), .B1(n_64_1_89), .B2(n_64_1_78), .ZN(
      n_64_210));
   NAND2_X1 i_64_1_38 (.A1(n_64_139), .A2(n_64_1_78), .ZN(n_64_1_25));
   OAI21_X1 i_64_1_39 (.A(n_64_1_26), .B1(n_64_1_90), .B2(n_64_1_78), .ZN(
      n_64_211));
   NAND2_X1 i_64_1_40 (.A1(n_64_140), .A2(n_64_1_78), .ZN(n_64_1_26));
   OAI21_X1 i_64_1_41 (.A(n_64_1_27), .B1(n_64_1_91), .B2(n_64_1_78), .ZN(
      n_64_212));
   NAND2_X1 i_64_1_42 (.A1(n_64_141), .A2(n_64_1_78), .ZN(n_64_1_27));
   OAI21_X1 i_64_1_43 (.A(n_64_1_28), .B1(n_64_1_92), .B2(n_64_1_78), .ZN(
      n_64_213));
   NAND2_X1 i_64_1_44 (.A1(n_64_142), .A2(n_64_1_78), .ZN(n_64_1_28));
   OAI21_X1 i_64_1_45 (.A(n_64_1_29), .B1(n_64_1_93), .B2(n_64_1_78), .ZN(
      n_64_214));
   NAND2_X1 i_64_1_46 (.A1(n_64_143), .A2(n_64_1_78), .ZN(n_64_1_29));
   OAI21_X1 i_64_1_47 (.A(n_64_1_30), .B1(n_64_1_94), .B2(n_64_1_78), .ZN(
      n_64_215));
   NAND2_X1 i_64_1_48 (.A1(n_64_144), .A2(n_64_1_78), .ZN(n_64_1_30));
   OAI21_X1 i_64_1_49 (.A(n_64_1_31), .B1(n_64_1_95), .B2(n_64_1_78), .ZN(
      n_64_216));
   NAND2_X1 i_64_1_50 (.A1(n_64_145), .A2(n_64_1_78), .ZN(n_64_1_31));
   OAI21_X1 i_64_1_51 (.A(n_64_1_32), .B1(n_64_1_96), .B2(n_64_1_78), .ZN(
      n_64_217));
   NAND2_X1 i_64_1_52 (.A1(n_64_146), .A2(n_64_1_78), .ZN(n_64_1_32));
   OAI21_X1 i_64_1_53 (.A(n_64_1_33), .B1(n_64_1_97), .B2(n_64_1_78), .ZN(
      n_64_218));
   NAND2_X1 i_64_1_54 (.A1(n_64_147), .A2(n_64_1_78), .ZN(n_64_1_33));
   OAI21_X1 i_64_1_55 (.A(n_64_1_34), .B1(n_64_1_98), .B2(n_64_1_78), .ZN(
      n_64_219));
   NAND2_X1 i_64_1_56 (.A1(n_64_148), .A2(n_64_1_78), .ZN(n_64_1_34));
   OAI21_X1 i_64_1_57 (.A(n_64_1_35), .B1(n_64_1_99), .B2(n_64_1_78), .ZN(
      n_64_220));
   NAND2_X1 i_64_1_58 (.A1(n_64_149), .A2(n_64_1_78), .ZN(n_64_1_35));
   OAI21_X1 i_64_1_59 (.A(n_64_1_36), .B1(n_64_1_100), .B2(n_64_1_78), .ZN(
      n_64_221));
   NAND2_X1 i_64_1_60 (.A1(n_64_150), .A2(n_64_1_78), .ZN(n_64_1_36));
   OAI21_X1 i_64_1_61 (.A(n_64_1_37), .B1(n_64_1_101), .B2(n_64_1_78), .ZN(
      n_64_222));
   NAND2_X1 i_64_1_62 (.A1(n_64_151), .A2(n_64_1_78), .ZN(n_64_1_37));
   OAI21_X1 i_64_1_63 (.A(n_64_1_38), .B1(n_64_1_102), .B2(n_64_1_78), .ZN(
      n_64_223));
   NAND2_X1 i_64_1_64 (.A1(n_64_152), .A2(n_64_1_78), .ZN(n_64_1_38));
   OAI21_X1 i_64_1_65 (.A(n_64_1_39), .B1(n_64_1_103), .B2(n_64_1_78), .ZN(
      n_64_224));
   NAND2_X1 i_64_1_66 (.A1(n_64_153), .A2(n_64_1_78), .ZN(n_64_1_39));
   OAI21_X1 i_64_1_67 (.A(n_64_1_40), .B1(n_64_1_104), .B2(n_64_1_78), .ZN(
      n_64_225));
   NAND2_X1 i_64_1_68 (.A1(n_64_154), .A2(n_64_1_78), .ZN(n_64_1_40));
   OAI21_X1 i_64_1_69 (.A(n_64_1_41), .B1(n_64_1_105), .B2(n_64_1_78), .ZN(
      n_64_226));
   NAND2_X1 i_64_1_70 (.A1(n_64_155), .A2(n_64_1_78), .ZN(n_64_1_41));
   OAI21_X1 i_64_1_71 (.A(n_64_1_42), .B1(n_64_1_106), .B2(n_64_1_78), .ZN(
      n_64_227));
   NAND2_X1 i_64_1_72 (.A1(n_64_156), .A2(n_64_1_78), .ZN(n_64_1_42));
   OAI21_X1 i_64_1_73 (.A(n_64_1_43), .B1(n_64_1_107), .B2(n_64_1_78), .ZN(
      n_64_228));
   NAND2_X1 i_64_1_74 (.A1(n_64_157), .A2(n_64_1_78), .ZN(n_64_1_43));
   OAI21_X1 i_64_1_75 (.A(n_64_1_44), .B1(n_64_1_108), .B2(n_64_1_78), .ZN(
      n_64_229));
   NAND2_X1 i_64_1_76 (.A1(n_64_158), .A2(n_64_1_78), .ZN(n_64_1_44));
   OAI21_X1 i_64_1_77 (.A(n_64_1_45), .B1(n_64_1_110), .B2(n_64_1_78), .ZN(
      n_64_230));
   NAND2_X1 i_64_1_78 (.A1(n_64_159), .A2(n_64_1_78), .ZN(n_64_1_45));
   OAI21_X1 i_64_1_79 (.A(n_64_1_46), .B1(n_64_1_113), .B2(n_64_1_78), .ZN(
      n_64_231));
   NAND2_X1 i_64_1_80 (.A1(n_64_160), .A2(n_64_1_78), .ZN(n_64_1_46));
   OAI21_X1 i_64_1_81 (.A(n_64_1_47), .B1(n_64_1_114), .B2(n_64_1_78), .ZN(
      n_64_232));
   NAND2_X1 i_64_1_82 (.A1(n_64_161), .A2(n_64_1_78), .ZN(n_64_1_47));
   OAI21_X1 i_64_1_83 (.A(n_64_1_48), .B1(n_64_1_115), .B2(n_64_1_78), .ZN(
      n_64_233));
   NAND2_X1 i_64_1_84 (.A1(n_64_162), .A2(n_64_1_78), .ZN(n_64_1_48));
   OAI21_X1 i_64_1_85 (.A(n_64_1_49), .B1(n_64_1_116), .B2(n_64_1_78), .ZN(
      n_64_234));
   NAND2_X1 i_64_1_86 (.A1(n_64_163), .A2(n_64_1_78), .ZN(n_64_1_49));
   OAI21_X1 i_64_1_87 (.A(n_64_1_50), .B1(n_64_1_117), .B2(n_64_1_78), .ZN(
      n_64_235));
   NAND2_X1 i_64_1_88 (.A1(n_64_164), .A2(n_64_1_78), .ZN(n_64_1_50));
   OAI21_X1 i_64_1_89 (.A(n_64_1_51), .B1(n_64_1_118), .B2(n_64_1_78), .ZN(
      n_64_236));
   NAND2_X1 i_64_1_90 (.A1(n_64_165), .A2(n_64_1_78), .ZN(n_64_1_51));
   OAI21_X1 i_64_1_91 (.A(n_64_1_52), .B1(n_64_1_119), .B2(n_64_1_78), .ZN(
      n_64_237));
   NAND2_X1 i_64_1_92 (.A1(n_64_166), .A2(n_64_1_78), .ZN(n_64_1_52));
   OAI21_X1 i_64_1_93 (.A(n_64_1_53), .B1(n_64_1_120), .B2(n_64_1_78), .ZN(
      n_64_238));
   NAND2_X1 i_64_1_94 (.A1(n_64_167), .A2(n_64_1_78), .ZN(n_64_1_53));
   OAI21_X1 i_64_1_95 (.A(n_64_1_54), .B1(n_64_1_121), .B2(n_64_1_78), .ZN(
      n_64_239));
   NAND2_X1 i_64_1_96 (.A1(n_64_168), .A2(n_64_1_78), .ZN(n_64_1_54));
   OAI21_X1 i_64_1_97 (.A(n_64_1_55), .B1(n_64_1_122), .B2(n_64_1_78), .ZN(
      n_64_240));
   NAND2_X1 i_64_1_98 (.A1(n_64_169), .A2(n_64_1_78), .ZN(n_64_1_55));
   OAI21_X1 i_64_1_99 (.A(n_64_1_56), .B1(n_64_1_123), .B2(n_64_1_78), .ZN(
      n_64_241));
   NAND2_X1 i_64_1_100 (.A1(n_64_170), .A2(n_64_1_78), .ZN(n_64_1_56));
   OAI21_X1 i_64_1_101 (.A(n_64_1_57), .B1(n_64_1_124), .B2(n_64_1_78), .ZN(
      n_64_242));
   NAND2_X1 i_64_1_102 (.A1(n_64_171), .A2(n_64_1_78), .ZN(n_64_1_57));
   OAI21_X1 i_64_1_103 (.A(n_64_1_58), .B1(n_64_1_125), .B2(n_64_1_78), .ZN(
      n_64_243));
   NAND2_X1 i_64_1_104 (.A1(n_64_172), .A2(n_64_1_78), .ZN(n_64_1_58));
   OAI21_X1 i_64_1_105 (.A(n_64_1_59), .B1(n_64_1_126), .B2(n_64_1_78), .ZN(
      n_64_244));
   NAND2_X1 i_64_1_106 (.A1(n_64_173), .A2(n_64_1_78), .ZN(n_64_1_59));
   OAI21_X1 i_64_1_107 (.A(n_64_1_60), .B1(n_64_1_127), .B2(n_64_1_78), .ZN(
      n_64_245));
   NAND2_X1 i_64_1_108 (.A1(n_64_174), .A2(n_64_1_78), .ZN(n_64_1_60));
   OAI21_X1 i_64_1_109 (.A(n_64_1_61), .B1(n_64_1_128), .B2(n_64_1_78), .ZN(
      n_64_246));
   NAND2_X1 i_64_1_110 (.A1(n_64_175), .A2(n_64_1_78), .ZN(n_64_1_61));
   OAI21_X1 i_64_1_111 (.A(n_64_1_62), .B1(n_64_1_129), .B2(n_64_1_78), .ZN(
      n_64_247));
   NAND2_X1 i_64_1_112 (.A1(n_64_176), .A2(n_64_1_78), .ZN(n_64_1_62));
   OAI21_X1 i_64_1_113 (.A(n_64_1_63), .B1(n_64_1_130), .B2(n_64_1_78), .ZN(
      n_64_248));
   NAND2_X1 i_64_1_114 (.A1(n_64_177), .A2(n_64_1_78), .ZN(n_64_1_63));
   OAI21_X1 i_64_1_115 (.A(n_64_1_64), .B1(n_64_1_131), .B2(n_64_1_78), .ZN(
      n_64_249));
   NAND2_X1 i_64_1_116 (.A1(n_64_178), .A2(n_64_1_78), .ZN(n_64_1_64));
   OAI21_X1 i_64_1_117 (.A(n_64_1_65), .B1(n_64_1_132), .B2(n_64_1_78), .ZN(
      n_64_250));
   NAND2_X1 i_64_1_118 (.A1(n_64_179), .A2(n_64_1_78), .ZN(n_64_1_65));
   OAI21_X1 i_64_1_119 (.A(n_64_1_66), .B1(n_64_1_133), .B2(n_64_1_78), .ZN(
      n_64_251));
   NAND2_X1 i_64_1_120 (.A1(n_64_180), .A2(n_64_1_78), .ZN(n_64_1_66));
   OAI21_X1 i_64_1_121 (.A(n_64_1_67), .B1(n_64_1_134), .B2(n_64_1_78), .ZN(
      n_64_252));
   NAND2_X1 i_64_1_122 (.A1(n_64_181), .A2(n_64_1_78), .ZN(n_64_1_67));
   OAI21_X1 i_64_1_123 (.A(n_64_1_68), .B1(n_64_1_135), .B2(n_64_1_78), .ZN(
      n_64_253));
   NAND2_X1 i_64_1_124 (.A1(n_64_182), .A2(n_64_1_78), .ZN(n_64_1_68));
   OAI21_X1 i_64_1_125 (.A(n_64_1_69), .B1(n_64_1_136), .B2(n_64_1_78), .ZN(
      n_64_254));
   NAND2_X1 i_64_1_126 (.A1(n_64_183), .A2(n_64_1_78), .ZN(n_64_1_69));
   OAI21_X1 i_64_1_127 (.A(n_64_1_70), .B1(n_64_1_137), .B2(n_64_1_78), .ZN(
      n_64_255));
   NAND2_X1 i_64_1_128 (.A1(n_64_184), .A2(n_64_1_78), .ZN(n_64_1_70));
   OAI21_X1 i_64_1_129 (.A(n_64_1_71), .B1(n_64_1_138), .B2(n_64_1_78), .ZN(
      n_64_256));
   NAND2_X1 i_64_1_130 (.A1(n_64_185), .A2(n_64_1_78), .ZN(n_64_1_71));
   OAI21_X1 i_64_1_131 (.A(n_64_1_72), .B1(n_64_1_139), .B2(n_64_1_78), .ZN(
      n_64_257));
   NAND2_X1 i_64_1_132 (.A1(n_64_186), .A2(n_64_1_78), .ZN(n_64_1_72));
   OAI21_X1 i_64_1_133 (.A(n_64_1_73), .B1(n_64_1_140), .B2(n_64_1_78), .ZN(
      n_64_258));
   NAND2_X1 i_64_1_134 (.A1(n_64_187), .A2(n_64_1_78), .ZN(n_64_1_73));
   OAI21_X1 i_64_1_135 (.A(n_64_1_74), .B1(n_64_1_141), .B2(n_64_1_78), .ZN(
      n_64_259));
   NAND2_X1 i_64_1_136 (.A1(n_64_188), .A2(n_64_1_78), .ZN(n_64_1_74));
   OAI21_X1 i_64_1_137 (.A(n_64_1_75), .B1(n_64_1_142), .B2(n_64_1_78), .ZN(
      n_64_260));
   NAND2_X1 i_64_1_138 (.A1(n_64_189), .A2(n_64_1_78), .ZN(n_64_1_75));
   NOR2_X1 i_64_1_145 (.A1(rst), .A2(n_64_1_114), .ZN(n_64_265));
   NOR2_X1 i_64_1_146 (.A1(rst), .A2(n_64_1_115), .ZN(n_64_266));
   NOR2_X1 i_64_1_147 (.A1(rst), .A2(n_64_1_116), .ZN(n_64_267));
   NOR2_X1 i_64_1_148 (.A1(rst), .A2(n_64_1_117), .ZN(n_64_268));
   NOR2_X1 i_64_1_149 (.A1(rst), .A2(n_64_1_118), .ZN(n_64_269));
   NOR2_X1 i_64_1_150 (.A1(rst), .A2(n_64_1_119), .ZN(n_64_270));
   NOR2_X1 i_64_1_151 (.A1(rst), .A2(n_64_1_120), .ZN(n_64_271));
   NOR2_X1 i_64_1_152 (.A1(rst), .A2(n_64_1_121), .ZN(n_64_272));
   NOR2_X1 i_64_1_153 (.A1(rst), .A2(n_64_1_122), .ZN(n_64_273));
   NOR2_X1 i_64_1_154 (.A1(rst), .A2(n_64_1_123), .ZN(n_64_274));
   NOR2_X1 i_64_1_155 (.A1(rst), .A2(n_64_1_124), .ZN(n_64_275));
   NOR2_X1 i_64_1_156 (.A1(rst), .A2(n_64_1_125), .ZN(n_64_276));
   NOR2_X1 i_64_1_157 (.A1(rst), .A2(n_64_1_126), .ZN(n_64_277));
   NOR2_X1 i_64_1_158 (.A1(rst), .A2(n_64_1_127), .ZN(n_64_278));
   NOR2_X1 i_64_1_159 (.A1(rst), .A2(n_64_1_128), .ZN(n_64_279));
   NOR2_X1 i_64_1_160 (.A1(rst), .A2(n_64_1_129), .ZN(n_64_280));
   NOR2_X1 i_64_1_161 (.A1(rst), .A2(n_64_1_130), .ZN(n_64_281));
   NOR2_X1 i_64_1_162 (.A1(rst), .A2(n_64_1_131), .ZN(n_64_282));
   NOR2_X1 i_64_1_163 (.A1(rst), .A2(n_64_1_132), .ZN(n_64_283));
   NOR2_X1 i_64_1_164 (.A1(rst), .A2(n_64_1_133), .ZN(n_64_284));
   NOR2_X1 i_64_1_165 (.A1(rst), .A2(n_64_1_134), .ZN(n_64_285));
   NOR2_X1 i_64_1_166 (.A1(rst), .A2(n_64_1_135), .ZN(n_64_286));
   NOR2_X1 i_64_1_167 (.A1(rst), .A2(n_64_1_136), .ZN(n_64_287));
   NOR2_X1 i_64_1_168 (.A1(rst), .A2(n_64_1_137), .ZN(n_64_288));
   NOR2_X1 i_64_1_169 (.A1(rst), .A2(n_64_1_138), .ZN(n_64_289));
   NOR2_X1 i_64_1_170 (.A1(rst), .A2(n_64_1_139), .ZN(n_64_290));
   NOR2_X1 i_64_1_171 (.A1(rst), .A2(n_64_1_140), .ZN(n_64_291));
   NOR2_X1 i_64_1_172 (.A1(rst), .A2(n_64_1_141), .ZN(n_64_292));
   NOR2_X1 i_64_1_173 (.A1(rst), .A2(n_64_1_142), .ZN(n_64_293));
   NOR2_X1 i_64_1_174 (.A1(rst), .A2(n_64_1_143), .ZN(n_64_294));
   NOR2_X1 i_64_1_175 (.A1(rst), .A2(n_64_1_144), .ZN(n_64_295));
   OR2_X1 i_64_1_176 (.A1(rst), .A2(en), .ZN(n_64_296));
   INV_X1 i_64_1_181 (.A(n_64_1_81), .ZN(n_64_300));
   OAI222_X1 i_64_1_182 (.A1(Q[4]), .A2(n_64_1_184), .B1(n_64_101), .B2(
      n_64_1_112), .C1(b[3]), .C2(n_64_1_109), .ZN(n_64_1_81));
   INV_X1 i_64_1_183 (.A(n_64_1_82), .ZN(n_64_301));
   OAI222_X1 i_64_1_184 (.A1(Q[5]), .A2(n_64_1_184), .B1(n_64_102), .B2(
      n_64_1_112), .C1(b[4]), .C2(n_64_1_109), .ZN(n_64_1_82));
   INV_X1 i_64_1_185 (.A(n_64_1_83), .ZN(n_64_302));
   OAI222_X1 i_64_1_186 (.A1(Q[6]), .A2(n_64_1_184), .B1(n_64_103), .B2(
      n_64_1_112), .C1(b[5]), .C2(n_64_1_109), .ZN(n_64_1_83));
   INV_X1 i_64_1_187 (.A(n_64_1_84), .ZN(n_64_303));
   OAI222_X1 i_64_1_188 (.A1(Q[7]), .A2(n_64_1_184), .B1(n_64_104), .B2(
      n_64_1_112), .C1(b[6]), .C2(n_64_1_109), .ZN(n_64_1_84));
   INV_X1 i_64_1_201 (.A(n_64_1_91), .ZN(n_64_310));
   OAI222_X1 i_64_1_202 (.A1(Q[14]), .A2(n_64_1_184), .B1(n_64_111), .B2(
      n_64_1_112), .C1(b[13]), .C2(n_64_1_109), .ZN(n_64_1_91));
   INV_X1 i_64_1_203 (.A(n_64_1_92), .ZN(n_64_311));
   OAI222_X1 i_64_1_204 (.A1(Q[15]), .A2(n_64_1_184), .B1(n_64_112), .B2(
      n_64_1_112), .C1(b[14]), .C2(n_64_1_109), .ZN(n_64_1_92));
   INV_X1 i_64_1_205 (.A(n_64_1_93), .ZN(n_64_312));
   OAI222_X1 i_64_1_206 (.A1(Q[16]), .A2(n_64_1_184), .B1(n_64_113), .B2(
      n_64_1_112), .C1(b[15]), .C2(n_64_1_109), .ZN(n_64_1_93));
   INV_X1 i_64_1_207 (.A(n_64_1_94), .ZN(n_64_313));
   OAI222_X1 i_64_1_208 (.A1(Q[17]), .A2(n_64_1_184), .B1(n_64_114), .B2(
      n_64_1_112), .C1(b[16]), .C2(n_64_1_109), .ZN(n_64_1_94));
   INV_X1 i_64_1_209 (.A(n_64_1_95), .ZN(n_64_314));
   OAI222_X1 i_64_1_210 (.A1(Q[18]), .A2(n_64_1_184), .B1(n_64_115), .B2(
      n_64_1_112), .C1(b[17]), .C2(n_64_1_109), .ZN(n_64_1_95));
   INV_X1 i_64_1_211 (.A(n_64_1_96), .ZN(n_64_315));
   OAI222_X1 i_64_1_212 (.A1(Q[19]), .A2(n_64_1_184), .B1(n_64_116), .B2(
      n_64_1_112), .C1(b[18]), .C2(n_64_1_109), .ZN(n_64_1_96));
   INV_X1 i_64_1_213 (.A(n_64_1_97), .ZN(n_64_316));
   OAI222_X1 i_64_1_214 (.A1(Q[20]), .A2(n_64_1_184), .B1(n_64_117), .B2(
      n_64_1_112), .C1(b[19]), .C2(n_64_1_109), .ZN(n_64_1_97));
   INV_X1 i_64_1_215 (.A(n_64_1_98), .ZN(n_64_317));
   OAI222_X1 i_64_1_216 (.A1(Q[21]), .A2(n_64_1_184), .B1(n_64_118), .B2(
      n_64_1_112), .C1(b[20]), .C2(n_64_1_109), .ZN(n_64_1_98));
   INV_X1 i_64_1_217 (.A(n_64_1_99), .ZN(n_64_318));
   OAI222_X1 i_64_1_218 (.A1(Q[22]), .A2(n_64_1_184), .B1(n_64_119), .B2(
      n_64_1_112), .C1(b[21]), .C2(n_64_1_109), .ZN(n_64_1_99));
   INV_X1 i_64_1_219 (.A(n_64_1_100), .ZN(n_64_319));
   OAI222_X1 i_64_1_220 (.A1(Q[23]), .A2(n_64_1_184), .B1(n_64_120), .B2(
      n_64_1_112), .C1(b[22]), .C2(n_64_1_109), .ZN(n_64_1_100));
   INV_X1 i_64_1_221 (.A(n_64_1_101), .ZN(n_64_320));
   OAI222_X1 i_64_1_222 (.A1(Q[24]), .A2(n_64_1_184), .B1(n_64_121), .B2(
      n_64_1_112), .C1(b[23]), .C2(n_64_1_109), .ZN(n_64_1_101));
   INV_X1 i_64_1_223 (.A(n_64_1_102), .ZN(n_64_321));
   OAI222_X1 i_64_1_224 (.A1(Q[25]), .A2(n_64_1_184), .B1(n_64_122), .B2(
      n_64_1_112), .C1(b[24]), .C2(n_64_1_109), .ZN(n_64_1_102));
   INV_X1 i_64_1_225 (.A(n_64_1_103), .ZN(n_64_322));
   OAI222_X1 i_64_1_226 (.A1(Q[26]), .A2(n_64_1_184), .B1(n_64_123), .B2(
      n_64_1_112), .C1(b[25]), .C2(n_64_1_109), .ZN(n_64_1_103));
   INV_X1 i_64_1_227 (.A(n_64_1_104), .ZN(n_64_323));
   OAI222_X1 i_64_1_228 (.A1(Q[27]), .A2(n_64_1_184), .B1(n_64_124), .B2(
      n_64_1_112), .C1(b[26]), .C2(n_64_1_109), .ZN(n_64_1_104));
   INV_X1 i_64_1_229 (.A(n_64_1_105), .ZN(n_64_324));
   OAI222_X1 i_64_1_230 (.A1(Q[28]), .A2(n_64_1_184), .B1(n_64_125), .B2(
      n_64_1_112), .C1(b[27]), .C2(n_64_1_109), .ZN(n_64_1_105));
   INV_X1 i_64_1_231 (.A(n_64_1_106), .ZN(n_64_325));
   OAI222_X1 i_64_1_232 (.A1(Q[29]), .A2(n_64_1_184), .B1(n_64_126), .B2(
      n_64_1_112), .C1(b[28]), .C2(n_64_1_109), .ZN(n_64_1_106));
   INV_X1 i_64_1_233 (.A(n_64_1_107), .ZN(n_64_326));
   OAI222_X1 i_64_1_234 (.A1(Q[30]), .A2(n_64_1_184), .B1(n_64_127), .B2(
      n_64_1_112), .C1(b[29]), .C2(n_64_1_109), .ZN(n_64_1_107));
   INV_X1 i_64_1_235 (.A(n_64_1_108), .ZN(n_64_327));
   OAI222_X1 i_64_1_236 (.A1(Q[31]), .A2(n_64_1_184), .B1(n_64_128), .B2(
      n_64_1_112), .C1(b[30]), .C2(n_64_1_109), .ZN(n_64_1_108));
   INV_X1 i_64_1_238 (.A(n_64_1_110), .ZN(n_64_328));
   AOI22_X1 i_64_1_239 (.A1(Q[32]), .A2(n_64_1_185), .B1(n_64_129), .B2(
      n_64_1_111), .ZN(n_64_1_110));
   INV_X1 i_64_1_240 (.A(n_64_1_112), .ZN(n_64_1_111));
   INV_X1 i_64_1_242 (.A(n_64_1_113), .ZN(n_64_329));
   AOI222_X1 i_64_1_243 (.A1(n_64_67), .A2(n_64_1_147), .B1(n_64_35), .B2(
      n_64_1_148), .C1(A[0]), .C2(n_64_1_146), .ZN(n_64_1_113));
   INV_X1 i_64_1_244 (.A(n_64_1_114), .ZN(n_64_330));
   AOI222_X1 i_64_1_245 (.A1(n_64_68), .A2(n_64_1_147), .B1(n_64_36), .B2(
      n_64_1_148), .C1(A[1]), .C2(n_64_1_146), .ZN(n_64_1_114));
   INV_X1 i_64_1_246 (.A(n_64_1_115), .ZN(n_64_331));
   AOI222_X1 i_64_1_247 (.A1(n_64_69), .A2(n_64_1_147), .B1(n_64_37), .B2(
      n_64_1_148), .C1(A[2]), .C2(n_64_1_146), .ZN(n_64_1_115));
   INV_X1 i_64_1_248 (.A(n_64_1_116), .ZN(n_64_332));
   AOI222_X1 i_64_1_249 (.A1(n_64_70), .A2(n_64_1_147), .B1(n_64_38), .B2(
      n_64_1_148), .C1(A[3]), .C2(n_64_1_146), .ZN(n_64_1_116));
   INV_X1 i_64_1_250 (.A(n_64_1_117), .ZN(n_64_333));
   AOI222_X1 i_64_1_251 (.A1(n_64_71), .A2(n_64_1_147), .B1(n_64_39), .B2(
      n_64_1_148), .C1(A[4]), .C2(n_64_1_146), .ZN(n_64_1_117));
   INV_X1 i_64_1_252 (.A(n_64_1_118), .ZN(n_64_334));
   AOI222_X1 i_64_1_253 (.A1(n_64_72), .A2(n_64_1_147), .B1(n_64_40), .B2(
      n_64_1_148), .C1(A[5]), .C2(n_64_1_146), .ZN(n_64_1_118));
   INV_X1 i_64_1_254 (.A(n_64_1_119), .ZN(n_64_335));
   AOI222_X1 i_64_1_255 (.A1(n_64_73), .A2(n_64_1_147), .B1(n_64_41), .B2(
      n_64_1_148), .C1(A[6]), .C2(n_64_1_146), .ZN(n_64_1_119));
   INV_X1 i_64_1_256 (.A(n_64_1_120), .ZN(n_64_336));
   AOI222_X1 i_64_1_257 (.A1(n_64_74), .A2(n_64_1_147), .B1(n_64_42), .B2(
      n_64_1_148), .C1(A[7]), .C2(n_64_1_146), .ZN(n_64_1_120));
   INV_X1 i_64_1_258 (.A(n_64_1_121), .ZN(n_64_337));
   AOI222_X1 i_64_1_259 (.A1(n_64_75), .A2(n_64_1_147), .B1(n_64_43), .B2(
      n_64_1_148), .C1(A[8]), .C2(n_64_1_146), .ZN(n_64_1_121));
   INV_X1 i_64_1_260 (.A(n_64_1_122), .ZN(n_64_338));
   AOI222_X1 i_64_1_261 (.A1(n_64_76), .A2(n_64_1_147), .B1(n_64_44), .B2(
      n_64_1_148), .C1(A[9]), .C2(n_64_1_146), .ZN(n_64_1_122));
   INV_X1 i_64_1_262 (.A(n_64_1_123), .ZN(n_64_339));
   AOI222_X1 i_64_1_263 (.A1(n_64_77), .A2(n_64_1_147), .B1(n_64_45), .B2(
      n_64_1_148), .C1(A[10]), .C2(n_64_1_146), .ZN(n_64_1_123));
   INV_X1 i_64_1_264 (.A(n_64_1_124), .ZN(n_64_340));
   AOI222_X1 i_64_1_265 (.A1(n_64_78), .A2(n_64_1_147), .B1(n_64_46), .B2(
      n_64_1_148), .C1(A[11]), .C2(n_64_1_146), .ZN(n_64_1_124));
   INV_X1 i_64_1_266 (.A(n_64_1_125), .ZN(n_64_341));
   AOI222_X1 i_64_1_267 (.A1(n_64_79), .A2(n_64_1_147), .B1(n_64_47), .B2(
      n_64_1_148), .C1(A[12]), .C2(n_64_1_146), .ZN(n_64_1_125));
   INV_X1 i_64_1_268 (.A(n_64_1_126), .ZN(n_64_342));
   AOI222_X1 i_64_1_269 (.A1(n_64_80), .A2(n_64_1_147), .B1(n_64_48), .B2(
      n_64_1_148), .C1(A[13]), .C2(n_64_1_146), .ZN(n_64_1_126));
   INV_X1 i_64_1_270 (.A(n_64_1_127), .ZN(n_64_343));
   AOI222_X1 i_64_1_271 (.A1(n_64_81), .A2(n_64_1_147), .B1(n_64_49), .B2(
      n_64_1_148), .C1(A[14]), .C2(n_64_1_146), .ZN(n_64_1_127));
   INV_X1 i_64_1_272 (.A(n_64_1_128), .ZN(n_64_344));
   AOI222_X1 i_64_1_273 (.A1(n_64_82), .A2(n_64_1_147), .B1(n_64_50), .B2(
      n_64_1_148), .C1(A[15]), .C2(n_64_1_146), .ZN(n_64_1_128));
   INV_X1 i_64_1_274 (.A(n_64_1_129), .ZN(n_64_345));
   AOI222_X1 i_64_1_275 (.A1(n_64_83), .A2(n_64_1_147), .B1(n_64_51), .B2(
      n_64_1_148), .C1(A[16]), .C2(n_64_1_146), .ZN(n_64_1_129));
   INV_X1 i_64_1_276 (.A(n_64_1_130), .ZN(n_64_346));
   AOI222_X1 i_64_1_277 (.A1(n_64_84), .A2(n_64_1_147), .B1(n_64_52), .B2(
      n_64_1_148), .C1(A[17]), .C2(n_64_1_146), .ZN(n_64_1_130));
   INV_X1 i_64_1_278 (.A(n_64_1_131), .ZN(n_64_347));
   AOI222_X1 i_64_1_279 (.A1(n_64_85), .A2(n_64_1_147), .B1(n_64_53), .B2(
      n_64_1_148), .C1(A[18]), .C2(n_64_1_146), .ZN(n_64_1_131));
   INV_X1 i_64_1_280 (.A(n_64_1_132), .ZN(n_64_348));
   AOI222_X1 i_64_1_281 (.A1(n_64_86), .A2(n_64_1_147), .B1(n_64_54), .B2(
      n_64_1_148), .C1(A[19]), .C2(n_64_1_146), .ZN(n_64_1_132));
   INV_X1 i_64_1_282 (.A(n_64_1_133), .ZN(n_64_349));
   AOI222_X1 i_64_1_283 (.A1(n_64_87), .A2(n_64_1_147), .B1(n_64_55), .B2(
      n_64_1_148), .C1(A[20]), .C2(n_64_1_146), .ZN(n_64_1_133));
   INV_X1 i_64_1_284 (.A(n_64_1_134), .ZN(n_64_350));
   AOI222_X1 i_64_1_285 (.A1(n_64_88), .A2(n_64_1_147), .B1(n_64_56), .B2(
      n_64_1_148), .C1(A[21]), .C2(n_64_1_146), .ZN(n_64_1_134));
   INV_X1 i_64_1_286 (.A(n_64_1_135), .ZN(n_64_351));
   AOI222_X1 i_64_1_287 (.A1(n_64_89), .A2(n_64_1_147), .B1(n_64_57), .B2(
      n_64_1_148), .C1(A[22]), .C2(n_64_1_146), .ZN(n_64_1_135));
   INV_X1 i_64_1_288 (.A(n_64_1_136), .ZN(n_64_352));
   AOI222_X1 i_64_1_289 (.A1(n_64_90), .A2(n_64_1_147), .B1(n_64_58), .B2(
      n_64_1_148), .C1(A[23]), .C2(n_64_1_146), .ZN(n_64_1_136));
   INV_X1 i_64_1_290 (.A(n_64_1_137), .ZN(n_64_353));
   AOI222_X1 i_64_1_291 (.A1(n_64_91), .A2(n_64_1_147), .B1(n_64_59), .B2(
      n_64_1_148), .C1(A[24]), .C2(n_64_1_146), .ZN(n_64_1_137));
   INV_X1 i_64_1_292 (.A(n_64_1_138), .ZN(n_64_354));
   AOI222_X1 i_64_1_293 (.A1(n_64_92), .A2(n_64_1_147), .B1(n_64_60), .B2(
      n_64_1_148), .C1(A[25]), .C2(n_64_1_146), .ZN(n_64_1_138));
   INV_X1 i_64_1_294 (.A(n_64_1_139), .ZN(n_64_355));
   AOI222_X1 i_64_1_295 (.A1(n_64_93), .A2(n_64_1_147), .B1(n_64_61), .B2(
      n_64_1_148), .C1(A[26]), .C2(n_64_1_146), .ZN(n_64_1_139));
   INV_X1 i_64_1_296 (.A(n_64_1_140), .ZN(n_64_356));
   AOI222_X1 i_64_1_297 (.A1(n_64_94), .A2(n_64_1_147), .B1(n_64_62), .B2(
      n_64_1_148), .C1(A[27]), .C2(n_64_1_146), .ZN(n_64_1_140));
   INV_X1 i_64_1_298 (.A(n_64_1_141), .ZN(n_64_357));
   AOI222_X1 i_64_1_299 (.A1(n_64_95), .A2(n_64_1_147), .B1(n_64_63), .B2(
      n_64_1_148), .C1(A[28]), .C2(n_64_1_146), .ZN(n_64_1_141));
   INV_X1 i_64_1_300 (.A(n_64_1_142), .ZN(n_64_358));
   AOI222_X1 i_64_1_301 (.A1(n_64_96), .A2(n_64_1_147), .B1(n_64_64), .B2(
      n_64_1_148), .C1(A[29]), .C2(n_64_1_146), .ZN(n_64_1_142));
   INV_X1 i_64_1_302 (.A(n_64_1_143), .ZN(n_64_359));
   INV_X1 i_64_1_304 (.A(n_64_1_144), .ZN(n_64_360));
   AND2_X1 i_64_1_306 (.A1(A[31]), .A2(n_64_1_146), .ZN(n_64_1_145));
   NOR2_X1 i_64_1_307 (.A1(n_64_1_148), .A2(n_64_1_147), .ZN(n_64_1_146));
   NOR3_X1 i_64_1_308 (.A1(n_64_1_193), .A2(n_64_1_184), .A3(Q[1]), .ZN(
      n_64_1_147));
   AOI21_X1 i_64_1_309 (.A(n_64_1_149), .B1(Q[0]), .B2(n_64_1_185), .ZN(
      n_64_1_148));
   INV_X1 i_64_1_310 (.A(n_64_1_149), .ZN(n_64_297));
   OAI22_X1 i_64_1_311 (.A1(Q[1]), .A2(n_64_1_184), .B1(b[0]), .B2(n_64_1_185), 
      .ZN(n_64_1_149));
   INV_X1 i_64_1_312 (.A(n_64_1_150), .ZN(n_64_361));
   AOI22_X1 i_64_1_313 (.A1(multiplicand[0]), .A2(n_64_1_185), .B1(a[0]), 
      .B2(n_64_1_184), .ZN(n_64_1_150));
   INV_X1 i_64_1_314 (.A(n_64_1_151), .ZN(n_64_362));
   AOI222_X1 i_64_1_315 (.A1(a[1]), .A2(n_64_1_181), .B1(multiplicand[1]), 
      .B2(n_64_1_185), .C1(n_64_4), .C2(n_64_1_183), .ZN(n_64_1_151));
   INV_X1 i_64_1_316 (.A(n_64_1_152), .ZN(n_64_363));
   AOI222_X1 i_64_1_317 (.A1(a[2]), .A2(n_64_1_181), .B1(multiplicand[2]), 
      .B2(n_64_1_185), .C1(n_64_5), .C2(n_64_1_183), .ZN(n_64_1_152));
   INV_X1 i_64_1_318 (.A(n_64_1_153), .ZN(n_64_364));
   AOI222_X1 i_64_1_319 (.A1(a[3]), .A2(n_64_1_181), .B1(multiplicand[3]), 
      .B2(n_64_1_185), .C1(n_64_6), .C2(n_64_1_183), .ZN(n_64_1_153));
   INV_X1 i_64_1_320 (.A(n_64_1_154), .ZN(n_64_365));
   AOI222_X1 i_64_1_321 (.A1(a[4]), .A2(n_64_1_181), .B1(multiplicand[4]), 
      .B2(n_64_1_185), .C1(n_64_7), .C2(n_64_1_183), .ZN(n_64_1_154));
   INV_X1 i_64_1_322 (.A(n_64_1_155), .ZN(n_64_366));
   AOI222_X1 i_64_1_323 (.A1(a[5]), .A2(n_64_1_181), .B1(multiplicand[5]), 
      .B2(n_64_1_185), .C1(n_64_8), .C2(n_64_1_183), .ZN(n_64_1_155));
   INV_X1 i_64_1_324 (.A(n_64_1_156), .ZN(n_64_367));
   AOI222_X1 i_64_1_325 (.A1(a[6]), .A2(n_64_1_181), .B1(multiplicand[6]), 
      .B2(n_64_1_185), .C1(n_64_9), .C2(n_64_1_183), .ZN(n_64_1_156));
   INV_X1 i_64_1_326 (.A(n_64_1_157), .ZN(n_64_368));
   AOI222_X1 i_64_1_327 (.A1(a[7]), .A2(n_64_1_181), .B1(multiplicand[7]), 
      .B2(n_64_1_185), .C1(n_64_10), .C2(n_64_1_183), .ZN(n_64_1_157));
   INV_X1 i_64_1_328 (.A(n_64_1_158), .ZN(n_64_369));
   AOI222_X1 i_64_1_329 (.A1(a[8]), .A2(n_64_1_181), .B1(multiplicand[8]), 
      .B2(n_64_1_185), .C1(n_64_11), .C2(n_64_1_183), .ZN(n_64_1_158));
   INV_X1 i_64_1_330 (.A(n_64_1_159), .ZN(n_64_370));
   AOI222_X1 i_64_1_331 (.A1(a[9]), .A2(n_64_1_181), .B1(multiplicand[9]), 
      .B2(n_64_1_185), .C1(n_64_12), .C2(n_64_1_183), .ZN(n_64_1_159));
   INV_X1 i_64_1_332 (.A(n_64_1_160), .ZN(n_64_371));
   AOI222_X1 i_64_1_333 (.A1(a[10]), .A2(n_64_1_181), .B1(multiplicand[10]), 
      .B2(n_64_1_185), .C1(n_64_13), .C2(n_64_1_183), .ZN(n_64_1_160));
   INV_X1 i_64_1_334 (.A(n_64_1_161), .ZN(n_64_372));
   AOI222_X1 i_64_1_335 (.A1(a[11]), .A2(n_64_1_181), .B1(multiplicand[11]), 
      .B2(n_64_1_185), .C1(n_64_14), .C2(n_64_1_183), .ZN(n_64_1_161));
   INV_X1 i_64_1_336 (.A(n_64_1_162), .ZN(n_64_373));
   AOI222_X1 i_64_1_337 (.A1(a[12]), .A2(n_64_1_181), .B1(multiplicand[12]), 
      .B2(n_64_1_185), .C1(n_64_15), .C2(n_64_1_183), .ZN(n_64_1_162));
   INV_X1 i_64_1_338 (.A(n_64_1_163), .ZN(n_64_374));
   AOI222_X1 i_64_1_339 (.A1(a[13]), .A2(n_64_1_181), .B1(multiplicand[13]), 
      .B2(n_64_1_185), .C1(n_64_16), .C2(n_64_1_183), .ZN(n_64_1_163));
   INV_X1 i_64_1_340 (.A(n_64_1_164), .ZN(n_64_375));
   AOI222_X1 i_64_1_341 (.A1(a[14]), .A2(n_64_1_181), .B1(multiplicand[14]), 
      .B2(n_64_1_185), .C1(n_64_17), .C2(n_64_1_183), .ZN(n_64_1_164));
   INV_X1 i_64_1_342 (.A(n_64_1_165), .ZN(n_64_376));
   AOI222_X1 i_64_1_343 (.A1(a[15]), .A2(n_64_1_181), .B1(multiplicand[15]), 
      .B2(n_64_1_185), .C1(n_64_18), .C2(n_64_1_183), .ZN(n_64_1_165));
   INV_X1 i_64_1_344 (.A(n_64_1_166), .ZN(n_64_377));
   AOI222_X1 i_64_1_345 (.A1(a[16]), .A2(n_64_1_181), .B1(multiplicand[16]), 
      .B2(n_64_1_185), .C1(n_64_19), .C2(n_64_1_183), .ZN(n_64_1_166));
   INV_X1 i_64_1_346 (.A(n_64_1_167), .ZN(n_64_378));
   AOI222_X1 i_64_1_347 (.A1(a[17]), .A2(n_64_1_181), .B1(multiplicand[17]), 
      .B2(n_64_1_185), .C1(n_64_20), .C2(n_64_1_183), .ZN(n_64_1_167));
   INV_X1 i_64_1_348 (.A(n_64_1_168), .ZN(n_64_379));
   AOI222_X1 i_64_1_349 (.A1(a[18]), .A2(n_64_1_181), .B1(multiplicand[18]), 
      .B2(n_64_1_185), .C1(n_64_21), .C2(n_64_1_183), .ZN(n_64_1_168));
   INV_X1 i_64_1_350 (.A(n_64_1_169), .ZN(n_64_380));
   AOI222_X1 i_64_1_351 (.A1(a[19]), .A2(n_64_1_181), .B1(multiplicand[19]), 
      .B2(n_64_1_185), .C1(n_64_22), .C2(n_64_1_183), .ZN(n_64_1_169));
   INV_X1 i_64_1_352 (.A(n_64_1_170), .ZN(n_64_381));
   AOI222_X1 i_64_1_353 (.A1(a[20]), .A2(n_64_1_181), .B1(multiplicand[20]), 
      .B2(n_64_1_185), .C1(n_64_23), .C2(n_64_1_183), .ZN(n_64_1_170));
   INV_X1 i_64_1_354 (.A(n_64_1_171), .ZN(n_64_382));
   AOI222_X1 i_64_1_355 (.A1(a[21]), .A2(n_64_1_181), .B1(multiplicand[21]), 
      .B2(n_64_1_185), .C1(n_64_24), .C2(n_64_1_183), .ZN(n_64_1_171));
   INV_X1 i_64_1_356 (.A(n_64_1_172), .ZN(n_64_383));
   AOI222_X1 i_64_1_357 (.A1(a[22]), .A2(n_64_1_181), .B1(multiplicand[22]), 
      .B2(n_64_1_185), .C1(n_64_25), .C2(n_64_1_183), .ZN(n_64_1_172));
   INV_X1 i_64_1_358 (.A(n_64_1_173), .ZN(n_64_384));
   AOI222_X1 i_64_1_359 (.A1(a[23]), .A2(n_64_1_181), .B1(multiplicand[23]), 
      .B2(n_64_1_185), .C1(n_64_26), .C2(n_64_1_183), .ZN(n_64_1_173));
   INV_X1 i_64_1_360 (.A(n_64_1_174), .ZN(n_64_385));
   AOI222_X1 i_64_1_361 (.A1(a[24]), .A2(n_64_1_181), .B1(multiplicand[24]), 
      .B2(n_64_1_185), .C1(n_64_27), .C2(n_64_1_183), .ZN(n_64_1_174));
   INV_X1 i_64_1_362 (.A(n_64_1_175), .ZN(n_64_386));
   AOI222_X1 i_64_1_363 (.A1(a[25]), .A2(n_64_1_181), .B1(multiplicand[25]), 
      .B2(n_64_1_185), .C1(n_64_28), .C2(n_64_1_183), .ZN(n_64_1_175));
   INV_X1 i_64_1_364 (.A(n_64_1_176), .ZN(n_64_387));
   AOI222_X1 i_64_1_365 (.A1(a[26]), .A2(n_64_1_181), .B1(multiplicand[26]), 
      .B2(n_64_1_185), .C1(n_64_29), .C2(n_64_1_183), .ZN(n_64_1_176));
   INV_X1 i_64_1_366 (.A(n_64_1_177), .ZN(n_64_388));
   AOI222_X1 i_64_1_367 (.A1(a[27]), .A2(n_64_1_181), .B1(multiplicand[27]), 
      .B2(n_64_1_185), .C1(n_64_30), .C2(n_64_1_183), .ZN(n_64_1_177));
   INV_X1 i_64_1_368 (.A(n_64_1_178), .ZN(n_64_389));
   AOI222_X1 i_64_1_369 (.A1(a[28]), .A2(n_64_1_181), .B1(multiplicand[28]), 
      .B2(n_64_1_185), .C1(n_64_31), .C2(n_64_1_183), .ZN(n_64_1_178));
   INV_X1 i_64_1_370 (.A(n_64_1_179), .ZN(n_64_390));
   AOI222_X1 i_64_1_371 (.A1(a[29]), .A2(n_64_1_181), .B1(multiplicand[29]), 
      .B2(n_64_1_185), .C1(n_64_32), .C2(n_64_1_183), .ZN(n_64_1_179));
   INV_X1 i_64_1_372 (.A(n_64_1_180), .ZN(n_64_391));
   AOI222_X1 i_64_1_373 (.A1(a[30]), .A2(n_64_1_181), .B1(multiplicand[30]), 
      .B2(n_64_1_185), .C1(n_64_33), .C2(n_64_1_183), .ZN(n_64_1_180));
   NOR2_X1 i_64_1_374 (.A1(a[31]), .A2(n_64_1_185), .ZN(n_64_1_181));
   INV_X1 i_64_1_375 (.A(n_64_1_182), .ZN(n_64_392));
   AOI22_X1 i_64_1_376 (.A1(multiplicand[31]), .A2(n_64_1_185), .B1(n_64_34), 
      .B2(n_64_1_183), .ZN(n_64_1_182));
   AND2_X1 i_64_1_377 (.A1(a[31]), .A2(n_64_1_184), .ZN(n_64_1_183));
   NOR4_X1 i_64_1_380 (.A1(SC[6]), .A2(SC[5]), .A3(SC[4]), .A4(SC[3]), .ZN(
      n_64_1_186));
   NOR3_X1 i_64_1_381 (.A1(SC[2]), .A2(SC[1]), .A3(SC[0]), .ZN(n_64_1_187));
   NAND2_X1 i_64_1_382 (.A1(n_64_264), .A2(n_64_1_189), .ZN(n_64_393));
   INV_X1 i_64_1_383 (.A(n_64_1_188), .ZN(n_64_394));
   OAI21_X1 i_64_1_384 (.A(n_64_264), .B1(n_64_3), .B2(n_64_1_190), .ZN(
      n_64_1_188));
   INV_X1 i_64_1_385 (.A(n_64_1_190), .ZN(n_64_1_189));
   NOR4_X1 i_64_1_386 (.A1(SC[6]), .A2(SC[5]), .A3(n_64_1_191), .A4(n_64_1_192), 
      .ZN(n_64_1_190));
   NAND2_X1 i_64_1_387 (.A1(SC[4]), .A2(SC[3]), .ZN(n_64_1_191));
   NAND3_X1 i_64_1_388 (.A1(SC[2]), .A2(SC[1]), .A3(SC[0]), .ZN(n_64_1_192));
   NOR2_X1 i_64_1_389 (.A1(rst), .A2(n_64_1_194), .ZN(n_64_264));
   INV_X1 i_64_1_390 (.A(Q[0]), .ZN(n_64_1_193));
   INV_X1 i_64_1_391 (.A(en), .ZN(n_64_1_194));
   INV_X1 i_64_1_139 (.A(n_64_1_79), .ZN(n_64_1_144));
   OAI21_X1 i_64_1_140 (.A(n_64_1_76), .B1(n_64_1_78), .B2(n_64_1_143), .ZN(
      n_64_261));
   AOI221_X1 i_64_1_141 (.A(n_64_1_145), .B1(n_64_65), .B2(n_64_1_148), .C1(
      n_64_97), .C2(n_64_1_147), .ZN(n_64_1_143));
   NAND2_X1 i_64_1_142 (.A1(n_64_190), .A2(n_64_1_78), .ZN(n_64_1_76));
   NAND2_X1 i_64_1_143 (.A1(n_64_1_200), .A2(n_64_1_77), .ZN(n_64_262));
   NAND2_X1 i_64_1_144 (.A1(n_64_1_79), .A2(n_64_1_202), .ZN(n_64_1_77));
   OAI221_X1 i_64_1_177 (.A(n_64_1_195), .B1(n_64_1_199), .B2(n_64_1_196), 
      .C1(n_64_1_198), .C2(n_64_1_197), .ZN(n_64_1_79));
   INV_X1 i_64_1_178 (.A(n_64_1_145), .ZN(n_64_1_195));
   INV_X1 i_64_1_179 (.A(n_64_1_148), .ZN(n_64_1_196));
   INV_X1 i_64_1_180 (.A(n_64_1_147), .ZN(n_64_1_197));
   INV_X1 i_64_1_189 (.A(n_64_98), .ZN(n_64_1_198));
   INV_X1 i_64_1_190 (.A(n_64_66), .ZN(n_64_1_199));
   NAND2_X1 i_64_1_191 (.A1(n_64_191), .A2(n_64_1_78), .ZN(n_64_1_200));
   INV_X1 i_64_1_192 (.A(n_64_1_201), .ZN(n_64_263));
   NAND2_X1 i_64_1_193 (.A1(n_64_192), .A2(n_64_1_78), .ZN(n_64_1_201));
   INV_X1 i_64_1_194 (.A(n_64_1_202), .ZN(n_64_1_78));
   NOR2_X1 i_64_1_195 (.A1(n_64_1_189), .A2(out_sign), .ZN(n_64_1_202));
   NOR2_X1 i_64_1_196 (.A1(n_64_1_204), .A2(n_64_1_203), .ZN(n_64_298));
   OAI22_X1 i_64_1_197 (.A1(n_64_1_109), .A2(b[1]), .B1(Q[2]), .B2(n_64_1_184), 
      .ZN(n_64_1_203));
   NOR2_X1 i_64_1_198 (.A1(n_64_99), .A2(n_64_1_112), .ZN(n_64_1_204));
   INV_X1 i_64_1_199 (.A(n_64_1_80), .ZN(n_64_299));
   OAI221_X1 i_64_1_200 (.A(n_64_1_205), .B1(Q[3]), .B2(n_64_1_184), .C1(
      n_64_100), .C2(n_64_1_112), .ZN(n_64_1_80));
   OR2_X1 i_64_1_237 (.A1(n_64_1_109), .A2(b[2]), .ZN(n_64_1_205));
   INV_X1 i_64_1_241 (.A(n_64_1_85), .ZN(n_64_304));
   OAI221_X1 i_64_1_303 (.A(n_64_1_206), .B1(Q[8]), .B2(n_64_1_184), .C1(
      n_64_105), .C2(n_64_1_112), .ZN(n_64_1_85));
   OR2_X1 i_64_1_305 (.A1(n_64_1_109), .A2(b[7]), .ZN(n_64_1_206));
   INV_X1 i_64_1_378 (.A(n_64_1_86), .ZN(n_64_305));
   OAI221_X1 i_64_1_379 (.A(n_64_1_207), .B1(Q[9]), .B2(n_64_1_184), .C1(
      n_64_106), .C2(n_64_1_112), .ZN(n_64_1_86));
   OR2_X1 i_64_1_392 (.A1(n_64_1_109), .A2(b[8]), .ZN(n_64_1_207));
   INV_X1 i_64_1_393 (.A(n_64_1_87), .ZN(n_64_306));
   OAI221_X1 i_64_1_394 (.A(n_64_1_208), .B1(Q[10]), .B2(n_64_1_184), .C1(
      n_64_107), .C2(n_64_1_112), .ZN(n_64_1_87));
   OR2_X1 i_64_1_395 (.A1(n_64_1_109), .A2(b[9]), .ZN(n_64_1_208));
   INV_X1 i_64_1_396 (.A(n_64_1_88), .ZN(n_64_307));
   OAI221_X1 i_64_1_397 (.A(n_64_1_209), .B1(Q[11]), .B2(n_64_1_184), .C1(
      n_64_108), .C2(n_64_1_112), .ZN(n_64_1_88));
   OR2_X1 i_64_1_398 (.A1(n_64_1_109), .A2(b[10]), .ZN(n_64_1_209));
   INV_X1 i_64_1_399 (.A(n_64_1_89), .ZN(n_64_308));
   OAI221_X1 i_64_1_400 (.A(n_64_1_210), .B1(Q[12]), .B2(n_64_1_184), .C1(
      n_64_109), .C2(n_64_1_112), .ZN(n_64_1_89));
   OR2_X1 i_64_1_401 (.A1(n_64_1_109), .A2(b[11]), .ZN(n_64_1_210));
   INV_X1 i_64_1_402 (.A(n_64_1_90), .ZN(n_64_309));
   OAI221_X1 i_64_1_403 (.A(n_64_1_211), .B1(Q[13]), .B2(n_64_1_184), .C1(
      n_64_110), .C2(n_64_1_112), .ZN(n_64_1_90));
   OR2_X1 i_64_1_404 (.A1(n_64_1_109), .A2(b[12]), .ZN(n_64_1_211));
   INV_X1 i_64_1_405 (.A(n_64_1_212), .ZN(n_64_1_109));
   NOR2_X1 i_64_1_406 (.A1(b[31]), .A2(n_64_1_185), .ZN(n_64_1_212));
   NAND2_X1 i_64_1_407 (.A1(n_64_1_184), .A2(b[31]), .ZN(n_64_1_112));
   INV_X1 i_64_1_408 (.A(n_64_1_185), .ZN(n_64_1_184));
   NAND2_X1 i_64_1_409 (.A1(n_64_1_186), .A2(n_64_1_187), .ZN(n_64_1_185));
endmodule
